DEPTH = 10240; % Memory depth and width are required % 
 % DEPTH is the number of addresses % 
WIDTH = 32; % WIDTH is the number of bits of data per word % 
% DEPTH and WIDTH should be entered as decimal numbers % 
ADDRESS_RADIX = HEX; % Address and value radixes are required % 
DATA_RADIX = HEX; % Enter BIN, DEC, HEX, OCT, or UNS; unless % 
 % otherwise specified, radixes = HEX % 
-- Specify values for addresses, which can be single address or range 
CONTENT 
BEGIN 
