
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80e5",
X"d0738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80e8",
X"f00c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580df",
X"fe2d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580de92",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80d9d404",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"775193b0",
X"3f83e080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3380e8f8",
X"0b80e8f8",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"52775192",
X"df3f83e0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583e0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"55b3923f",
X"83e08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"811451b2",
X"aa3f83e0",
X"80083070",
X"83e08008",
X"07802583",
X"e0800c53",
X"863d0d04",
X"fc3d0d76",
X"70525599",
X"cb3f83e0",
X"80085481",
X"5383e080",
X"0880c738",
X"7451998e",
X"3f83e080",
X"080b0b80",
X"e7b05383",
X"e0800852",
X"53ff8f3f",
X"83e08008",
X"a5380b0b",
X"80e7b452",
X"7251fefe",
X"3f83e080",
X"0894380b",
X"0b80e7b8",
X"527251fe",
X"ed3f83e0",
X"8008802e",
X"83388154",
X"73537283",
X"e0800c86",
X"3d0d04fd",
X"3d0d7570",
X"525498e4",
X"3f815383",
X"e0800898",
X"38735198",
X"ad3f83e0",
X"a0085283",
X"e0800851",
X"feb43f83",
X"e0800853",
X"7283e080",
X"0c853d0d",
X"04e03d0d",
X"a33d0870",
X"525e8ed3",
X"3f83e080",
X"0833943d",
X"56547394",
X"3880ea80",
X"52745184",
X"c7397d52",
X"785191d6",
X"3f84d139",
X"7d518ebb",
X"3f83e080",
X"08527451",
X"8deb3f83",
X"e0a80852",
X"933d7052",
X"5d94c63f",
X"83e08008",
X"59800b83",
X"e0800855",
X"5b83e080",
X"087b2e94",
X"38811b74",
X"525b97c7",
X"3f83e080",
X"085483e0",
X"8008ee38",
X"805aff7a",
X"437a427a",
X"415f7909",
X"709f2c7b",
X"065b547a",
X"7a248438",
X"ff1b5af6",
X"1a700970",
X"9f2c7206",
X"7bff125a",
X"5a525555",
X"80752595",
X"38765197",
X"863f83e0",
X"800876ff",
X"18585557",
X"738024ed",
X"38747f2e",
X"873880c2",
X"db3f745f",
X"78ff1b70",
X"585d5880",
X"7a259538",
X"775196db",
X"3f83e080",
X"0876ff18",
X"58555873",
X"8024ed38",
X"800b83e7",
X"bc0c800b",
X"83e7e00c",
X"0b0b80e7",
X"bc518bae",
X"3f81800b",
X"83e7e00c",
X"0b0b80e7",
X"c4518b9e",
X"3fa80b83",
X"e7bc0c76",
X"802e80e8",
X"3883e7bc",
X"08777932",
X"70307072",
X"07802570",
X"872b83e7",
X"e00c5156",
X"78535656",
X"968e3f83",
X"e0800880",
X"2e8a380b",
X"0b80e7cc",
X"518ae33f",
X"765195ce",
X"3f83e080",
X"08520b0b",
X"80e88051",
X"8ad03f76",
X"5195d43f",
X"83e08008",
X"83e7bc08",
X"55577574",
X"258638a8",
X"1656f739",
X"7583e7bc",
X"0c86f076",
X"24ff9438",
X"87980b83",
X"e7bc0c77",
X"802eb738",
X"7751958a",
X"3f83e080",
X"08785255",
X"95aa3f0b",
X"0b80e7d4",
X"5483e080",
X"088f3887",
X"39807634",
X"fd95390b",
X"0b80e7d0",
X"54745373",
X"520b0b80",
X"e7a05189",
X"e93f8054",
X"0b0b80e7",
X"a85189de",
X"3f811454",
X"73a82e09",
X"8106ed38",
X"868da051",
X"bed13f80",
X"52903d70",
X"525480cc",
X"e63f8352",
X"735180cc",
X"de3f6180",
X"2e80ff38",
X"7b5473ff",
X"2e963878",
X"802e8180",
X"38785194",
X"aa3f83e0",
X"8008ff15",
X"5559e739",
X"78802e80",
X"eb387851",
X"94a63f83",
X"e0800880",
X"2efc8338",
X"785193ee",
X"3f83e080",
X"08520b0b",
X"80e7ac51",
X"abcc3f83",
X"e08008a4",
X"387c51ad",
X"843f83e0",
X"80085574",
X"ff165654",
X"807425fb",
X"ee38741d",
X"70335556",
X"73af2efe",
X"c838e839",
X"785193ac",
X"3f83e080",
X"08527c51",
X"acbb3ffb",
X"ce397f88",
X"29601005",
X"7a056105",
X"5afbff39",
X"a23d0d04",
X"803d0d90",
X"80f83370",
X"81ff0670",
X"842a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"a80b9080",
X"f834b80b",
X"9080f834",
X"7083e080",
X"0c823d0d",
X"04803d0d",
X"9080f833",
X"7081ff06",
X"70852a81",
X"32708106",
X"51515151",
X"70802e8d",
X"38980b90",
X"80f834b8",
X"0b9080f8",
X"347083e0",
X"800c823d",
X"0d04930b",
X"9080fc34",
X"ff0b9080",
X"e83404ff",
X"3d0d028f",
X"05335280",
X"0b9080fc",
X"348a51bc",
X"a63fdf3f",
X"80f80b90",
X"80e03480",
X"0b9080c8",
X"34fa1252",
X"719080c0",
X"34800b90",
X"80d83471",
X"9080d034",
X"9080f852",
X"807234b8",
X"7234833d",
X"0d04803d",
X"0d028b05",
X"33517090",
X"80f434fe",
X"bf3f83e0",
X"8008802e",
X"f638823d",
X"0d04803d",
X"0d853980",
X"c5a23ffe",
X"d83f83e0",
X"8008802e",
X"f2389080",
X"f4337081",
X"ff0683e0",
X"800c5182",
X"3d0d0480",
X"3d0da30b",
X"9080fc34",
X"ff0b9080",
X"e8349080",
X"f851a871",
X"34b87134",
X"823d0d04",
X"803d0d90",
X"80fc3370",
X"81c00670",
X"30708025",
X"83e0800c",
X"51515182",
X"3d0d0480",
X"3d0d9080",
X"f8337081",
X"ff067083",
X"2a813270",
X"81065151",
X"51517080",
X"2ee838b0",
X"0b9080f8",
X"34b80b90",
X"80f83482",
X"3d0d0480",
X"3d0d9080",
X"ac088106",
X"83e0800c",
X"823d0d04",
X"fd3d0d75",
X"77545480",
X"73259438",
X"73708105",
X"55335280",
X"e7d85185",
X"a13fff13",
X"53e93985",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"80c8f53f",
X"83e08008",
X"7a27ed38",
X"74802e80",
X"e0387452",
X"755180c8",
X"df3f83e0",
X"80087553",
X"76525480",
X"c9853f83",
X"e080087a",
X"53755256",
X"80c8c53f",
X"83e08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"e08008c2",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9c",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fbfd3f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd13f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbad3f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83e0900c",
X"7183e094",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383e090",
X"085283e0",
X"940851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"99d25351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fd3d",
X"0d757052",
X"54a3c23f",
X"83e08008",
X"14537274",
X"2e9238ff",
X"13703353",
X"5371af2e",
X"098106ee",
X"38811353",
X"7283e080",
X"0c853d0d",
X"04fd3d0d",
X"75777053",
X"5454c73f",
X"83e08008",
X"732ea138",
X"83e08008",
X"733152ff",
X"125271ff",
X"2e8f3872",
X"70810554",
X"33747081",
X"055634eb",
X"39ff1454",
X"80743485",
X"3d0d0480",
X"3d0d7251",
X"ff903f82",
X"3d0d0471",
X"83e0800c",
X"04803d0d",
X"72518071",
X"34810bbc",
X"120c800b",
X"80c0120c",
X"823d0d04",
X"800b83e2",
X"d408248a",
X"38a4ac3f",
X"ff0b83e2",
X"d40c800b",
X"83e0800c",
X"04ff3d0d",
X"735283e0",
X"b008722e",
X"8d38d93f",
X"71519697",
X"3f7183e0",
X"b00c833d",
X"0d04f43d",
X"0d7e6062",
X"5c5a5581",
X"54bc1508",
X"81913874",
X"51cf3f79",
X"58807a25",
X"80f73883",
X"e3840870",
X"892a5783",
X"ff067884",
X"80723156",
X"56577378",
X"25833873",
X"557583e2",
X"d4082e84",
X"38ff893f",
X"83e2d408",
X"8025a638",
X"75892b51",
X"98da3f83",
X"e384088f",
X"3dfc1155",
X"5c548152",
X"f81b5196",
X"c43f7614",
X"83e3840c",
X"7583e2d4",
X"0c745376",
X"527851a2",
X"dd3f83e0",
X"800883e3",
X"84081683",
X"e3840c78",
X"7631761b",
X"5b595677",
X"8024ff8b",
X"38617a71",
X"0c547554",
X"75802e83",
X"38815473",
X"83e0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"9b3f7651",
X"feaf3f86",
X"3dfc0553",
X"78527751",
X"95e73f79",
X"75710c54",
X"83e08008",
X"5483e080",
X"08802e83",
X"38815473",
X"83e0800c",
X"863d0d04",
X"fe3d0d75",
X"83e2d408",
X"53538072",
X"24893871",
X"732e8438",
X"fdd63f74",
X"51fdea3f",
X"725197ac",
X"3f83e080",
X"085283e0",
X"8008802e",
X"83388152",
X"7183e080",
X"0c843d0d",
X"04803d0d",
X"7280c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d72bc11",
X"0883e080",
X"0c51823d",
X"0d0480c4",
X"0b83e080",
X"0c04fd3d",
X"0d757771",
X"54705355",
X"539f9a3f",
X"82c81308",
X"bc150c82",
X"c0130880",
X"c0150cfc",
X"eb3f7351",
X"93a93f73",
X"83e0b00c",
X"83e08008",
X"5383e080",
X"08802e83",
X"38815372",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"775553fc",
X"bf3f7280",
X"2ea538bc",
X"13085273",
X"519ea43f",
X"83e08008",
X"8f387752",
X"7251ff9a",
X"3f83e080",
X"08538a39",
X"82cc1308",
X"53d83981",
X"537283e0",
X"800c853d",
X"0d04fe3d",
X"0dff0b83",
X"e2d40c74",
X"83e0b40c",
X"7583e2d0",
X"0c9f913f",
X"83e08008",
X"81ff0652",
X"81537199",
X"3883e2ec",
X"518e933f",
X"83e08008",
X"5283e080",
X"08802e83",
X"38725271",
X"537283e0",
X"800c843d",
X"0d04fa3d",
X"0d787a82",
X"c4120882",
X"c4120870",
X"72245956",
X"56575773",
X"732e0981",
X"06913880",
X"c0165280",
X"c017519c",
X"953f83e0",
X"80085574",
X"83e0800c",
X"883d0d04",
X"f63d0d7c",
X"5b807b71",
X"5c54577a",
X"772e8c38",
X"811a82cc",
X"1408545a",
X"72f63880",
X"5980d939",
X"7a548157",
X"80707b7b",
X"315a5755",
X"ff185374",
X"732580c1",
X"3882cc14",
X"08527351",
X"ff8c3f80",
X"0b83e080",
X"0825a138",
X"82cc1408",
X"82cc1108",
X"82cc160c",
X"7482cc12",
X"0c537580",
X"2e863872",
X"82cc170c",
X"72548057",
X"7382cc15",
X"08811757",
X"5556ffb8",
X"39811959",
X"800bff1b",
X"54547873",
X"25833881",
X"54768132",
X"70750651",
X"5372ff90",
X"388c3d0d",
X"04f73d0d",
X"7b7d5a5a",
X"82d05283",
X"e2d00851",
X"bbfe3f83",
X"e0800857",
X"f9e23f79",
X"5283e2d8",
X"5195b43f",
X"83e08008",
X"54805383",
X"e0800873",
X"2e098106",
X"82833883",
X"e0b4080b",
X"0b80e7ac",
X"53705256",
X"9bd33f0b",
X"0b80e7ac",
X"5280c016",
X"519bc63f",
X"75bc170c",
X"7382c017",
X"0c810b82",
X"c4170c81",
X"0b82c817",
X"0c7382cc",
X"170cff17",
X"82d01755",
X"57819139",
X"83e0c033",
X"70822a70",
X"81065154",
X"55728180",
X"3874812a",
X"81065877",
X"80f63874",
X"842a8106",
X"82c4150c",
X"83e0c033",
X"810682c8",
X"150c7952",
X"73519aed",
X"3f73519b",
X"843f83e0",
X"80081453",
X"af737081",
X"05553472",
X"bc150c83",
X"e0c15272",
X"519ace3f",
X"83e0b808",
X"82c0150c",
X"83e0ce52",
X"80c01451",
X"9abb3f78",
X"802e8d38",
X"7351782d",
X"83e08008",
X"802e9938",
X"7782cc15",
X"0c75802e",
X"86387382",
X"cc170c73",
X"82d015ff",
X"19595556",
X"76802e9b",
X"3883e0b8",
X"5283e2d8",
X"5194aa3f",
X"83e08008",
X"8a3883e0",
X"c1335372",
X"fed23878",
X"802e8938",
X"83e0b408",
X"51fcb93f",
X"83e0b408",
X"537283e0",
X"800c8b3d",
X"0d04ff3d",
X"0d805273",
X"51fdb63f",
X"833d0d04",
X"f03d0d62",
X"705254f6",
X"913f83e0",
X"80087453",
X"873d7053",
X"5555f6b1",
X"3ff7913f",
X"7351d33f",
X"63537452",
X"83e08008",
X"51fab93f",
X"923d0d04",
X"7183e080",
X"0c0480c0",
X"1283e080",
X"0c04803d",
X"0d7282c0",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"cc110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"82c41108",
X"83e0800c",
X"51823d0d",
X"04f93d0d",
X"7983e098",
X"08575781",
X"77278196",
X"38768817",
X"0827818e",
X"38753355",
X"74822e89",
X"3874832e",
X"b33880fe",
X"39745476",
X"1083fe06",
X"5376882a",
X"8c170805",
X"52893dfc",
X"055199c0",
X"3f83e080",
X"0880df38",
X"029d0533",
X"893d3371",
X"882b0756",
X"5680d139",
X"84547682",
X"2b83fc06",
X"5376872a",
X"8c170805",
X"52893dfc",
X"05519990",
X"3f83e080",
X"08b03802",
X"9f053302",
X"84059e05",
X"3371982b",
X"71902b07",
X"028c059d",
X"05337088",
X"2b72078d",
X"3d337180",
X"fffffe80",
X"06075152",
X"53575856",
X"83398155",
X"7483e080",
X"0c893d0d",
X"04fb3d0d",
X"83e09808",
X"fe198812",
X"08fe0555",
X"56548056",
X"7473278d",
X"38821433",
X"75712994",
X"16080557",
X"537583e0",
X"800c873d",
X"0d04fc3d",
X"0d765280",
X"0b83e098",
X"08703351",
X"52537083",
X"2e098106",
X"91389512",
X"33941333",
X"71982b71",
X"902b0755",
X"55519b12",
X"339a1333",
X"71882b07",
X"740783e0",
X"800c5586",
X"3d0d04fc",
X"3d0d7683",
X"e0980855",
X"55807523",
X"88150853",
X"72812e88",
X"38881408",
X"73268538",
X"8152b239",
X"72903873",
X"33527183",
X"2e098106",
X"85389014",
X"0853728c",
X"160c7280",
X"2e8d3872",
X"51fed63f",
X"83e08008",
X"52853990",
X"14085271",
X"90160c80",
X"527183e0",
X"800c863d",
X"0d04fa3d",
X"0d7883e0",
X"98087122",
X"81057083",
X"ffff0657",
X"54575573",
X"802e8838",
X"90150853",
X"72863883",
X"5280e739",
X"738f0652",
X"7180da38",
X"81139016",
X"0c8c1508",
X"53729038",
X"830b8417",
X"22575273",
X"762780c6",
X"38bf3982",
X"1633ff05",
X"74842a06",
X"5271b238",
X"7251fcb1",
X"3f815271",
X"83e08008",
X"27a83883",
X"5283e080",
X"08881708",
X"279c3883",
X"e080088c",
X"160c83e0",
X"800851fd",
X"bc3f83e0",
X"80089016",
X"0c737523",
X"80527183",
X"e0800c88",
X"3d0d04f2",
X"3d0d6062",
X"64585e5b",
X"75335574",
X"a02e0981",
X"06883881",
X"16704456",
X"ef396270",
X"33565674",
X"af2e0981",
X"06843881",
X"1643800b",
X"881c0c62",
X"70335155",
X"749f2691",
X"387a51fd",
X"d23f83e0",
X"80085680",
X"7d348381",
X"39933d84",
X"1c087058",
X"595f8a55",
X"a0767081",
X"055834ff",
X"155574ff",
X"2e098106",
X"ef388070",
X"5a5c887f",
X"085f5a7b",
X"811d7081",
X"ff066013",
X"703370af",
X"327030a0",
X"73277180",
X"25075151",
X"525b535e",
X"57557480",
X"e73876ae",
X"2e098106",
X"83388155",
X"787a2775",
X"07557480",
X"2e9f3879",
X"88327030",
X"78ae3270",
X"30707307",
X"9f2a5351",
X"57515675",
X"bb388859",
X"8b5affab",
X"3976982b",
X"55748025",
X"873880e4",
X"e0173357",
X"ff9f1755",
X"74992689",
X"38e01770",
X"81ff0658",
X"5578811a",
X"7081ff06",
X"721b535b",
X"57557675",
X"34fef839",
X"7b1e7f0c",
X"805576a0",
X"26833881",
X"55748b19",
X"347a51fc",
X"823f83e0",
X"800880f5",
X"38a0547a",
X"2270852b",
X"83e00654",
X"55901b08",
X"527c5193",
X"cb3f83e0",
X"80085783",
X"e0800881",
X"81387c33",
X"5574802e",
X"80f4388b",
X"1d337083",
X"2a708106",
X"51565674",
X"b4388b7d",
X"841d0883",
X"e0800859",
X"5b5b58ff",
X"185877ff",
X"2e9a3879",
X"7081055b",
X"33797081",
X"055b3371",
X"71315256",
X"5675802e",
X"e2388639",
X"75802e96",
X"387a51fb",
X"e53fff86",
X"3983e080",
X"085683e0",
X"8008b638",
X"83397656",
X"841b088b",
X"11335155",
X"74a7388b",
X"1d337084",
X"2a708106",
X"51565674",
X"89388356",
X"94398156",
X"90397c51",
X"fa943f83",
X"e0800888",
X"1c0cfd81",
X"397583e0",
X"800c903d",
X"0d04f83d",
X"0d7a7c59",
X"57825483",
X"fe537752",
X"76519290",
X"3f835683",
X"e0800880",
X"ec388117",
X"33773371",
X"882b0756",
X"56825674",
X"82d4d52e",
X"09810680",
X"d4387554",
X"b6537752",
X"765191e4",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"ac388254",
X"80d25377",
X"52765191",
X"bb3f83e0",
X"80089838",
X"81173377",
X"3371882b",
X"0783e080",
X"08525656",
X"748182c6",
X"2e833881",
X"567583e0",
X"800c8a3d",
X"0d04eb3d",
X"0d675a80",
X"0b83e098",
X"0c90dd3f",
X"83e08008",
X"81065582",
X"567483ee",
X"38747553",
X"8f3d7053",
X"5759feca",
X"3f83e080",
X"0881ff06",
X"5776812e",
X"09810680",
X"d4389054",
X"83be5374",
X"52755190",
X"cf3f83e0",
X"800880c9",
X"388f3d33",
X"5574802e",
X"80c93802",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"70587b57",
X"5e525e57",
X"5957fdee",
X"3f83e080",
X"0881ff06",
X"5776832e",
X"09810686",
X"38815682",
X"f1397680",
X"2e863886",
X"5682e739",
X"a4548d53",
X"78527551",
X"8fe63f81",
X"5683e080",
X"0882d338",
X"02be0533",
X"028405bd",
X"05337188",
X"2b07595d",
X"77ab3802",
X"80ce0533",
X"02840580",
X"cd053371",
X"982b7190",
X"2b07973d",
X"3370882b",
X"72070294",
X"0580cb05",
X"33710754",
X"525e5759",
X"5602b705",
X"33787129",
X"028805b6",
X"0533028c",
X"05b50533",
X"71882b07",
X"701d707f",
X"8c050c5f",
X"5957595d",
X"8e3d3382",
X"1b3402b9",
X"0533903d",
X"3371882b",
X"075a5c78",
X"841b2302",
X"bb053302",
X"8405ba05",
X"3371882b",
X"07565c74",
X"ab380280",
X"ca053302",
X"840580c9",
X"05337198",
X"2b71902b",
X"07963d33",
X"70882b72",
X"07029405",
X"80c70533",
X"71075152",
X"53575e5c",
X"74763178",
X"3179842a",
X"903d3354",
X"71713153",
X"5656ace4",
X"3f83e080",
X"08820570",
X"881c0c83",
X"e08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83e0980c",
X"80567583",
X"e0800c97",
X"3d0d04e9",
X"3d0d83e0",
X"98085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e63f83e0",
X"80085483",
X"e0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f48a",
X"3f83e080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383e080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83e09808",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0ea3f",
X"83e08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"843f83e0",
X"80085583",
X"e0800880",
X"2eff8938",
X"83e08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"518a8d3f",
X"83e08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83e0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83e09808",
X"55568555",
X"73802e81",
X"e1388114",
X"33810653",
X"84557280",
X"2e81d338",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b7388214",
X"3370892b",
X"56537680",
X"2eb53874",
X"52ff1651",
X"a7e63f83",
X"e08008ff",
X"18765470",
X"535853a7",
X"d73f83e0",
X"80087326",
X"96387430",
X"70780670",
X"98170c77",
X"7131a417",
X"08525851",
X"538939a0",
X"140870a4",
X"160c5374",
X"7627b938",
X"7251eed9",
X"3f83e080",
X"0853810b",
X"83e08008",
X"278b3888",
X"140883e0",
X"80082688",
X"38800b81",
X"1534b039",
X"83e08008",
X"a4150c98",
X"14081598",
X"150c7575",
X"3156c439",
X"98140816",
X"7098160c",
X"735256ef",
X"c83f83e0",
X"80088c38",
X"83e08008",
X"81153481",
X"55943982",
X"1433ff05",
X"76892a06",
X"83e08008",
X"05a8150c",
X"80557483",
X"e0800c88",
X"3d0d04ef",
X"3d0d6356",
X"855583e0",
X"9808802e",
X"80d23893",
X"3df40584",
X"170c6453",
X"883d7053",
X"765257f1",
X"d23f83e0",
X"80085583",
X"e08008b4",
X"38883d33",
X"5473802e",
X"a13802a7",
X"05337084",
X"2a708106",
X"51555583",
X"5573802e",
X"97387651",
X"eef83f83",
X"e0800888",
X"170c7551",
X"efa93f83",
X"e0800855",
X"7483e080",
X"0c933d0d",
X"04e43d0d",
X"6ea13d08",
X"405e8556",
X"83e09808",
X"802e8485",
X"389e3df4",
X"05841f0c",
X"7e98387d",
X"51eef83f",
X"83e08008",
X"5683ee39",
X"814181f6",
X"39834181",
X"f139933d",
X"7f960541",
X"59807f82",
X"95055e56",
X"756081ff",
X"05348341",
X"901e0876",
X"2e81d338",
X"a0547d22",
X"70852b83",
X"e0065458",
X"901e0852",
X"78518698",
X"3f83e080",
X"084183e0",
X"8008ffb8",
X"3878335c",
X"7b802eff",
X"b4388b19",
X"3370bf06",
X"71810652",
X"43557480",
X"2e80de38",
X"7b81bf06",
X"55748f24",
X"80d3389a",
X"19335574",
X"80cb38f3",
X"1d70585d",
X"8156758b",
X"2e098106",
X"85388e56",
X"8b39759a",
X"2e098106",
X"83389c56",
X"75197070",
X"81055233",
X"7133811a",
X"821a5f5b",
X"525b5574",
X"86387977",
X"34853980",
X"df773477",
X"7b57577a",
X"a02e0981",
X"06c03881",
X"567b81e5",
X"32703070",
X"9f2a5151",
X"557bae2e",
X"93387480",
X"2e8e3861",
X"832a7081",
X"06515574",
X"802e9738",
X"7d51ede2",
X"3f83e080",
X"084183e0",
X"80088738",
X"901e08fe",
X"af388060",
X"3475802e",
X"88387c52",
X"7f5183a5",
X"3f60802e",
X"8638800b",
X"901f0c60",
X"5660832e",
X"85386081",
X"d038891f",
X"57901e08",
X"802e81a8",
X"38805675",
X"19703351",
X"5574a02e",
X"a0387485",
X"2e098106",
X"843881e5",
X"55747770",
X"81055934",
X"81167081",
X"ff065755",
X"877627d7",
X"38881933",
X"5574a02e",
X"a938ae77",
X"70810559",
X"34885675",
X"19703351",
X"5574a02e",
X"95387477",
X"70810559",
X"34811670",
X"81ff0657",
X"558a7627",
X"e2388b19",
X"337f8805",
X"349f1933",
X"9e1a3371",
X"982b7190",
X"2b079d1c",
X"3370882b",
X"72079c1e",
X"33710764",
X"0c52991d",
X"33981e33",
X"71882b07",
X"53515357",
X"5956747f",
X"84052397",
X"1933961a",
X"3371882b",
X"07565674",
X"7f860523",
X"8077347d",
X"51ebf33f",
X"83e08008",
X"83327030",
X"7072079f",
X"2c83e080",
X"08065256",
X"56961f33",
X"55748a38",
X"891f5296",
X"1f5181b1",
X"3f7583e0",
X"800c9e3d",
X"0d04fd3d",
X"0d757753",
X"54733351",
X"70893871",
X"33517080",
X"2ea13873",
X"33723352",
X"53727127",
X"8538ff51",
X"94397073",
X"27853881",
X"518b3981",
X"14811353",
X"54d33980",
X"517083e0",
X"800c853d",
X"0d04fd3d",
X"0d757754",
X"54723370",
X"81ff0652",
X"5270802e",
X"a3387181",
X"ff068114",
X"ffbf1253",
X"54527099",
X"268938a0",
X"127081ff",
X"06535171",
X"74708105",
X"5634d239",
X"80743485",
X"3d0d04ff",
X"bd3d0d80",
X"c63d0852",
X"a53d7052",
X"54ffb33f",
X"80c73d08",
X"52853d70",
X"5253ffa6",
X"3f725273",
X"51fedf3f",
X"80c53d0d",
X"04fe3d0d",
X"74765353",
X"71708105",
X"53335170",
X"73708105",
X"553470f0",
X"38843d0d",
X"04fe3d0d",
X"74528072",
X"33525370",
X"732e8d38",
X"81128114",
X"71335354",
X"5270f538",
X"7283e080",
X"0c843d0d",
X"04fc3d0d",
X"76557483",
X"e398082e",
X"af388053",
X"745187c1",
X"3f83e080",
X"0881ff06",
X"ff147081",
X"ff067230",
X"709f2a51",
X"52555354",
X"72802e84",
X"3871dd38",
X"73fe3874",
X"83e3980c",
X"863d0d04",
X"ff3d0dff",
X"0b83e398",
X"0c84a53f",
X"81518785",
X"3f83e080",
X"0881ff06",
X"5271ee38",
X"81d33f71",
X"83e0800c",
X"833d0d04",
X"fc3d0d76",
X"028405a2",
X"05220288",
X"05a60522",
X"7a545555",
X"55ff823f",
X"72802ea0",
X"3883e3ac",
X"14337570",
X"81055734",
X"81147083",
X"ffff06ff",
X"157083ff",
X"ff065652",
X"5552dd39",
X"800b83e0",
X"800c863d",
X"0d04fc3d",
X"0d76787a",
X"11565355",
X"80537174",
X"2e933872",
X"15517033",
X"83e3ac13",
X"34811281",
X"145452ea",
X"39800b83",
X"e0800c86",
X"3d0d04fd",
X"3d0d9054",
X"83e39808",
X"5186f43f",
X"83e08008",
X"81ff06ff",
X"15713071",
X"30707307",
X"9f2a729f",
X"2a065255",
X"52555372",
X"db38853d",
X"0d04803d",
X"0d83e3a4",
X"081083e3",
X"9c080790",
X"80a80c82",
X"3d0d0480",
X"0b83e3a4",
X"0ce43f04",
X"810b83e3",
X"a40cdb3f",
X"04ed3f04",
X"7183e3a0",
X"0c04803d",
X"0d8051f4",
X"3f810b83",
X"e3a40c81",
X"0b83e39c",
X"0cffbb3f",
X"823d0d04",
X"803d0d72",
X"30707407",
X"802583e3",
X"9c0c51ff",
X"a53f823d",
X"0d04803d",
X"0d028b05",
X"339080a4",
X"0c9080a8",
X"08708106",
X"515170f5",
X"389080a4",
X"087081ff",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d81ff51",
X"d13f83e0",
X"800881ff",
X"0683e080",
X"0c823d0d",
X"04803d0d",
X"73902b73",
X"079080b4",
X"0c823d0d",
X"0404fb3d",
X"0d780284",
X"059f0533",
X"70982b55",
X"57557280",
X"259b3875",
X"80ff0656",
X"805280f7",
X"51e03f83",
X"e0800881",
X"ff065473",
X"812680ff",
X"388051fe",
X"e73fffa2",
X"3f8151fe",
X"df3fff9a",
X"3f7551fe",
X"ed3f7498",
X"2a51fee6",
X"3f74902a",
X"7081ff06",
X"5253feda",
X"3f74882a",
X"7081ff06",
X"5253fece",
X"3f7481ff",
X"0651fec6",
X"3f815575",
X"80c02e09",
X"81068638",
X"8195558d",
X"397580c8",
X"2e098106",
X"84388187",
X"557451fe",
X"a53f8a55",
X"fec83f83",
X"e0800881",
X"ff067098",
X"2b545472",
X"80258c38",
X"ff157081",
X"ff065653",
X"74e23873",
X"83e0800c",
X"873d0d04",
X"fa3d0dfd",
X"c53f8051",
X"fdda3f8a",
X"54fe933f",
X"ff147081",
X"ff065553",
X"73f33873",
X"74535580",
X"c051fea6",
X"3f83e080",
X"0881ff06",
X"5473812e",
X"09810682",
X"9f3883aa",
X"5280c851",
X"fe8c3f83",
X"e0800881",
X"ff065372",
X"812e0981",
X"0681a838",
X"7454873d",
X"74115456",
X"fdc83f83",
X"e0800873",
X"34811470",
X"81ff0655",
X"53837427",
X"e538029a",
X"05335372",
X"812e0981",
X"0681d938",
X"029b0533",
X"5380ce90",
X"547281aa",
X"2e8d3881",
X"c73980e4",
X"518ac03f",
X"ff145473",
X"802e81b8",
X"38820a52",
X"81e951fd",
X"a53f83e0",
X"800881ff",
X"065372de",
X"38725280",
X"fa51fd92",
X"3f83e080",
X"0881ff06",
X"53728190",
X"38725473",
X"1653fcd6",
X"3f83e080",
X"08733481",
X"147081ff",
X"06555383",
X"7427e838",
X"873d3370",
X"862a7081",
X"06515454",
X"8c557280",
X"e3388455",
X"80de3974",
X"5281e951",
X"fccc3f83",
X"e0800881",
X"ff065382",
X"5581e956",
X"81732786",
X"38735580",
X"c15680ce",
X"90548a39",
X"80e45189",
X"b23fff14",
X"5473802e",
X"a9388052",
X"7551fc9a",
X"3f83e080",
X"0881ff06",
X"5372e138",
X"84805280",
X"d051fc86",
X"3f83e080",
X"0881ff06",
X"5372802e",
X"83388055",
X"7483e3a8",
X"348051fb",
X"873ffbc2",
X"3f883d0d",
X"04fb3d0d",
X"7754800b",
X"83e3a833",
X"70832a70",
X"81065155",
X"57557275",
X"2e098106",
X"85387389",
X"2b547352",
X"80d151fb",
X"bd3f83e0",
X"800881ff",
X"065372bd",
X"3882b8c0",
X"54fb833f",
X"83e08008",
X"81ff0653",
X"7281ff2e",
X"09810689",
X"38ff1454",
X"73e7389f",
X"397281fe",
X"2e098106",
X"963883e7",
X"ac5283e3",
X"ac51faed",
X"3ffad33f",
X"fad03f83",
X"39815580",
X"51fa893f",
X"fac43f74",
X"81ff0683",
X"e0800c87",
X"3d0d04fb",
X"3d0d7783",
X"e3ac5654",
X"8151f9ec",
X"3f83e3a8",
X"3370832a",
X"70810651",
X"54567285",
X"3873892b",
X"54735280",
X"d851fab6",
X"3f83e080",
X"0881ff06",
X"537280e4",
X"3881ff51",
X"f9d43f81",
X"fe51f9ce",
X"3f848053",
X"74708105",
X"563351f9",
X"c13fff13",
X"7083ffff",
X"06515372",
X"eb387251",
X"f9b03f72",
X"51f9ab3f",
X"f9d03f83",
X"e080089f",
X"0653a788",
X"5472852e",
X"8c389939",
X"80e45186",
X"ea3fff14",
X"54f9b33f",
X"83e08008",
X"81ff2e84",
X"3873e938",
X"8051f8e4",
X"3ff99f3f",
X"800b83e0",
X"800c873d",
X"0d047183",
X"e7b00c88",
X"80800b83",
X"e7ac0c84",
X"80800b83",
X"e7b40c04",
X"f03d0d83",
X"80805683",
X"e7b00816",
X"83e7ac08",
X"17565474",
X"33743483",
X"e7b40816",
X"54807434",
X"81165675",
X"8380a02e",
X"098106db",
X"3883d080",
X"5683e7b0",
X"081683e7",
X"ac081756",
X"54743374",
X"3483e7b4",
X"08165480",
X"74348116",
X"567583d0",
X"a02e0981",
X"06db3883",
X"a8805683",
X"e7b00816",
X"83e7ac08",
X"17565474",
X"33743483",
X"e7b40816",
X"54807434",
X"81165675",
X"83a8902e",
X"098106db",
X"38805683",
X"e7b00816",
X"83e7b408",
X"17555573",
X"33753481",
X"16567581",
X"80802e09",
X"8106e438",
X"86fe3f89",
X"3d58a253",
X"80e6e052",
X"77519afb",
X"3f80578c",
X"805683e7",
X"b4081677",
X"19555573",
X"33753481",
X"16811858",
X"5676a22e",
X"098106e6",
X"38860b87",
X"a8833480",
X"0b87a882",
X"34800b87",
X"809a34af",
X"0b878096",
X"34bf0b87",
X"80973480",
X"0b878098",
X"349f0b87",
X"80993480",
X"0b87809b",
X"34f80b87",
X"a8893476",
X"87a88034",
X"820b87d0",
X"8f34820b",
X"87a88134",
X"923d0d04",
X"fe3d0d80",
X"5383e7b4",
X"081383e7",
X"b0081452",
X"52703372",
X"34811353",
X"72818080",
X"2e098106",
X"e4388380",
X"805383e7",
X"b4081383",
X"e7b00814",
X"52527033",
X"72348113",
X"53728380",
X"a02e0981",
X"06e43883",
X"d0805383",
X"e7b40813",
X"83e7b008",
X"14525270",
X"33723481",
X"13537283",
X"d0a02e09",
X"8106e438",
X"83a88053",
X"83e7b408",
X"1383e7b0",
X"08145252",
X"70337234",
X"81135372",
X"83a8902e",
X"098106e4",
X"38843d0d",
X"04803d0d",
X"90809008",
X"810683e0",
X"800c823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087081",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fd0676",
X"1007720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870822c",
X"bf0683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe830676",
X"822b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087088",
X"2c870683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f1ff06",
X"76882b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"8b2cbf06",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f88f",
X"ff06768b",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870912c",
X"bf0683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fc87ffff",
X"0676912b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70992c81",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870ff",
X"bf0a0676",
X"992b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"80087088",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"892c8106",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708a2c81",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708b2c",
X"810683e0",
X"800c5182",
X"3d0d04fe",
X"3d0d7481",
X"e629872a",
X"9080a00c",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d818080",
X"53805288",
X"800a51ff",
X"b33fa080",
X"53805282",
X"800a51c7",
X"3f843d0d",
X"04803d0d",
X"8151fc92",
X"3f72802e",
X"90388051",
X"fe943fce",
X"3f80e9ec",
X"3351fe8a",
X"3f8151fc",
X"a33f8051",
X"fc9e3f80",
X"51fbef3f",
X"823d0d04",
X"fd3d0d75",
X"52805480",
X"ff722588",
X"38810bff",
X"80135354",
X"ffbf1251",
X"70992686",
X"38e01252",
X"9e39ff9f",
X"12519971",
X"279538d0",
X"12e01370",
X"54545189",
X"71278838",
X"8f732783",
X"38805273",
X"802e8538",
X"81801252",
X"7181ff06",
X"83e0800c",
X"853d0d04",
X"803d0d84",
X"d8c05180",
X"71708105",
X"53347084",
X"e0c02e09",
X"8106f038",
X"823d0d04",
X"fe3d0d02",
X"97053351",
X"ff863f83",
X"e0800881",
X"ff0683e7",
X"bc085452",
X"8073249b",
X"3883e7dc",
X"08137283",
X"e7e00807",
X"53537173",
X"3483e7bc",
X"08810583",
X"e7bc0c84",
X"3d0d04fa",
X"3d0d8280",
X"0a1b5580",
X"57883dfc",
X"05547953",
X"74527851",
X"cbe23f88",
X"3d0d04fe",
X"3d0d83e7",
X"d4085274",
X"51d2c53f",
X"83e08008",
X"8c387653",
X"755283e7",
X"d40851c7",
X"3f843d0d",
X"04fe3d0d",
X"83e7d408",
X"53755274",
X"51cd853f",
X"83e08008",
X"8d387753",
X"765283e7",
X"d40851ff",
X"a23f843d",
X"0d04fd3d",
X"0d83e7d4",
X"0851cbf9",
X"3f83e080",
X"0890802e",
X"098106ad",
X"38805483",
X"c1808053",
X"83e08008",
X"5283e7d4",
X"0851fef3",
X"3f87c180",
X"80143387",
X"c1908015",
X"34811454",
X"7390802e",
X"098106e9",
X"38853d0d",
X"0480e7e0",
X"0b83e080",
X"0c04f73d",
X"0d805a80",
X"59805880",
X"705757fd",
X"e73f800b",
X"83e7bc0c",
X"800b83e7",
X"e00c80e7",
X"e451c6de",
X"3f81800b",
X"83e7e00c",
X"80e7e851",
X"c6d03f80",
X"d00b83e7",
X"bc0c7530",
X"70770780",
X"2570872b",
X"83e7e00c",
X"5154f982",
X"3f83e080",
X"085280e7",
X"f051c6aa",
X"3f80f80b",
X"83e7bc0c",
X"75813270",
X"30707207",
X"80257087",
X"2b83e7e0",
X"0c515555",
X"ff833f83",
X"e0800852",
X"80e7fc51",
X"c6803f81",
X"a00b83e7",
X"bc0c7582",
X"32703070",
X"72078025",
X"70872b83",
X"e7e00c51",
X"5583e7d4",
X"085255c7",
X"9a3f83e0",
X"80085280",
X"e88451c5",
X"d13f81c8",
X"0b83e7bc",
X"0c758332",
X"70307072",
X"07802570",
X"872b83e7",
X"e00c5155",
X"80e88c52",
X"55c5af3f",
X"81f00b83",
X"e7bc0c75",
X"84327030",
X"70720780",
X"2570872b",
X"83e7e00c",
X"515580e8",
X"9c5255c5",
X"8d3f8298",
X"0b83e7bc",
X"0c758532",
X"70307072",
X"07802570",
X"872b83e7",
X"e00c5155",
X"80e8b452",
X"55c4eb3f",
X"82c00b83",
X"e7bc0c75",
X"86327030",
X"70720780",
X"2570872b",
X"83e7e00c",
X"515580e8",
X"cc5255c4",
X"c93f868d",
X"a051f9c7",
X"3f805288",
X"3d705254",
X"87dd3f83",
X"52735187",
X"d63f7816",
X"56758025",
X"85388056",
X"90398676",
X"25853886",
X"56873975",
X"862682db",
X"38758429",
X"80e78405",
X"54730804",
X"f6d43f83",
X"e0800878",
X"56547481",
X"2e098106",
X"893883e0",
X"80081054",
X"903974ff",
X"2e098106",
X"883883e0",
X"8008812c",
X"54907425",
X"85389054",
X"88397380",
X"24833881",
X"547351f6",
X"ae3f828f",
X"39f6c03f",
X"83e08008",
X"18547380",
X"25853880",
X"54883987",
X"74258338",
X"87547351",
X"f6ba3f81",
X"ee397787",
X"3879802e",
X"81e53883",
X"e0a40883",
X"e0a00c8b",
X"df0b83e0",
X"a80c83e7",
X"d40851ff",
X"b5e73ffb",
X"b53f81c7",
X"3979802e",
X"81c13883",
X"e09c0883",
X"e0a00c8b",
X"df0b83e0",
X"a80c83e7",
X"d00851ff",
X"b5c33f75",
X"832e0981",
X"06943881",
X"80805382",
X"80805283",
X"e7d00851",
X"fa993f81",
X"87397584",
X"2e098106",
X"af388280",
X"80538180",
X"805283e7",
X"d00851f9",
X"fe3f8054",
X"84828080",
X"14338481",
X"80801534",
X"81145473",
X"8180802e",
X"098106e8",
X"3880d139",
X"75852e09",
X"810680c8",
X"38805481",
X"80805380",
X"c0805283",
X"e7d00851",
X"f9c53f82",
X"80805380",
X"c0805283",
X"e7d00851",
X"f9b53f84",
X"81808014",
X"338481c0",
X"80153484",
X"82808014",
X"338482c0",
X"80153481",
X"14547380",
X"c0802e09",
X"8106dc38",
X"81548c39",
X"79873876",
X"802efac3",
X"38805473",
X"83e0800c",
X"8b3d0d04",
X"ff3d0df5",
X"d63f83e0",
X"8008802e",
X"86388051",
X"80dd39f5",
X"db3f83e0",
X"800880d1",
X"38f5fb3f",
X"83e08008",
X"802eaa38",
X"8151f38a",
X"3fefd13f",
X"800b83e7",
X"bc0cf9f2",
X"3f83e080",
X"0852ff0b",
X"83e7bc0c",
X"f1d63f71",
X"a4387151",
X"f2e83fa2",
X"39f5b23f",
X"83e08008",
X"802e9738",
X"8151f2d6",
X"3fef9d3f",
X"ff0b83e7",
X"bc0cf1b0",
X"3f8151f6",
X"ac3f833d",
X"0d04fc3d",
X"0d908080",
X"52868480",
X"8051c682",
X"3f83e080",
X"08b83880",
X"e9f051ca",
X"c53f83e0",
X"800883e7",
X"d4085480",
X"e8d85383",
X"e0800852",
X"55c5a13f",
X"83e08008",
X"8438f8aa",
X"3f818080",
X"54828080",
X"5380e8d4",
X"527451f7",
X"f43f8151",
X"f5d73ffe",
X"b73ffc39",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"0280e8e4",
X"0b83e0a4",
X"0c80e8e8",
X"0b83e09c",
X"0c80e8ec",
X"0b83e0ac",
X"0c83e08c",
X"08fc050c",
X"800b83e7",
X"c00b83e0",
X"8c08f805",
X"0c83e08c",
X"08f4050c",
X"c3f03f83",
X"e0800886",
X"05fc0683",
X"e08c08f0",
X"050c0283",
X"e08c08f0",
X"0508310d",
X"833d7083",
X"e08c08f8",
X"05087084",
X"0583e08c",
X"08f8050c",
X"0c51c0b9",
X"3f83e08c",
X"08f40508",
X"810583e0",
X"8c08f405",
X"0c83e08c",
X"08f40508",
X"872e0981",
X"06ffad38",
X"86948080",
X"51ed833f",
X"ff0b83e7",
X"bc0c800b",
X"83e7e00c",
X"84d8c00b",
X"83e7dc0c",
X"8151f0b6",
X"3f8151f0",
X"db3f8051",
X"f0d63f81",
X"51f0fc3f",
X"8151f1d1",
X"3f8251f1",
X"9f3f8051",
X"f1f53f80",
X"51f29f3f",
X"80d0c452",
X"8051ffbd",
X"f23ffdc6",
X"3f83e08c",
X"08fc0508",
X"0d800b83",
X"e0800c87",
X"3d0d83e0",
X"8c0c04fd",
X"3d0d7554",
X"80740c80",
X"0b84150c",
X"800b8815",
X"0c87d089",
X"3387d08f",
X"3370822a",
X"70810670",
X"30707207",
X"7009709f",
X"2c77069e",
X"06545151",
X"55515153",
X"53807298",
X"06525370",
X"882e0981",
X"06833881",
X"53709832",
X"70307080",
X"25757131",
X"84180c51",
X"51518072",
X"86065253",
X"70822e09",
X"81068338",
X"81537086",
X"32703070",
X"80257571",
X"31770c51",
X"51517194",
X"32703070",
X"80258817",
X"0c515185",
X"3d0d04fe",
X"3d0d7476",
X"54527151",
X"feed3f72",
X"812ea238",
X"8173268d",
X"3872822e",
X"ab387283",
X"2e9f38e6",
X"397108e2",
X"38841208",
X"dd388812",
X"08d838a0",
X"39881208",
X"812e0981",
X"06cc3894",
X"39881208",
X"812e8d38",
X"71088938",
X"84120880",
X"2effb738",
X"843d0d04",
X"83e08c08",
X"0283e08c",
X"0cfd3d0d",
X"805383e0",
X"8c088c05",
X"085283e0",
X"8c088805",
X"085183d4",
X"3f83e080",
X"087083e0",
X"800c5485",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"fd3d0d81",
X"5383e08c",
X"088c0508",
X"5283e08c",
X"08880508",
X"5183a13f",
X"83e08008",
X"7083e080",
X"0c54853d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cf9",
X"3d0d800b",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"05088025",
X"b93883e0",
X"8c088805",
X"083083e0",
X"8c088805",
X"0c800b83",
X"e08c08f4",
X"050c83e0",
X"8c08fc05",
X"088a3881",
X"0b83e08c",
X"08f4050c",
X"83e08c08",
X"f4050883",
X"e08c08fc",
X"050c83e0",
X"8c088c05",
X"088025b9",
X"3883e08c",
X"088c0508",
X"3083e08c",
X"088c050c",
X"800b83e0",
X"8c08f005",
X"0c83e08c",
X"08fc0508",
X"8a38810b",
X"83e08c08",
X"f0050c83",
X"e08c08f0",
X"050883e0",
X"8c08fc05",
X"0c805383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"05085181",
X"df3f83e0",
X"80087083",
X"e08c08f8",
X"050c5483",
X"e08c08fc",
X"0508802e",
X"903883e0",
X"8c08f805",
X"083083e0",
X"8c08f805",
X"0c83e08c",
X"08f80508",
X"7083e080",
X"0c54893d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cfb",
X"3d0d800b",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"05088025",
X"993883e0",
X"8c088805",
X"083083e0",
X"8c088805",
X"0c810b83",
X"e08c08fc",
X"050c83e0",
X"8c088c05",
X"08802590",
X"3883e08c",
X"088c0508",
X"3083e08c",
X"088c050c",
X"815383e0",
X"8c088c05",
X"085283e0",
X"8c088805",
X"0851bd3f",
X"83e08008",
X"7083e08c",
X"08f8050c",
X"5483e08c",
X"08fc0508",
X"802e9038",
X"83e08c08",
X"f8050830",
X"83e08c08",
X"f8050c83",
X"e08c08f8",
X"05087083",
X"e0800c54",
X"873d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cfd3d0d",
X"810b83e0",
X"8c08fc05",
X"0c800b83",
X"e08c08f8",
X"050c83e0",
X"8c088c05",
X"0883e08c",
X"08880508",
X"27b93883",
X"e08c08fc",
X"0508802e",
X"ae38800b",
X"83e08c08",
X"8c050824",
X"a23883e0",
X"8c088c05",
X"081083e0",
X"8c088c05",
X"0c83e08c",
X"08fc0508",
X"1083e08c",
X"08fc050c",
X"ffb83983",
X"e08c08fc",
X"0508802e",
X"80e13883",
X"e08c088c",
X"050883e0",
X"8c088805",
X"0826ad38",
X"83e08c08",
X"88050883",
X"e08c088c",
X"05083183",
X"e08c0888",
X"050c83e0",
X"8c08f805",
X"0883e08c",
X"08fc0508",
X"0783e08c",
X"08f8050c",
X"83e08c08",
X"fc050881",
X"2a83e08c",
X"08fc050c",
X"83e08c08",
X"8c050881",
X"2a83e08c",
X"088c050c",
X"ff953983",
X"e08c0890",
X"0508802e",
X"933883e0",
X"8c088805",
X"087083e0",
X"8c08f405",
X"0c519139",
X"83e08c08",
X"f8050870",
X"83e08c08",
X"f4050c51",
X"83e08c08",
X"f4050883",
X"e0800c85",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"ff3d0d80",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"88050881",
X"06ff1170",
X"097083e0",
X"8c088c05",
X"080683e0",
X"8c08fc05",
X"081183e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"812a83e0",
X"8c088805",
X"0c83e08c",
X"088c0508",
X"1083e08c",
X"088c050c",
X"51515151",
X"83e08c08",
X"88050880",
X"2e8438ff",
X"ab3983e0",
X"8c08fc05",
X"087083e0",
X"800c5183",
X"3d0d83e0",
X"8c0c04fc",
X"3d0d7670",
X"797b5555",
X"55558f72",
X"278c3872",
X"75078306",
X"5170802e",
X"a938ff12",
X"5271ff2e",
X"98387270",
X"81055433",
X"74708105",
X"5634ff12",
X"5271ff2e",
X"098106ea",
X"387483e0",
X"800c863d",
X"0d047451",
X"72708405",
X"54087170",
X"8405530c",
X"72708405",
X"54087170",
X"8405530c",
X"72708405",
X"54087170",
X"8405530c",
X"72708405",
X"54087170",
X"8405530c",
X"f0125271",
X"8f26c938",
X"83722795",
X"38727084",
X"05540871",
X"70840553",
X"0cfc1252",
X"718326ed",
X"387054ff",
X"81390000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00002aa8",
X"00002ae9",
X"00002b0a",
X"00002b31",
X"00002b31",
X"00002b31",
X"00002bf4",
X"25732025",
X"73000000",
X"20000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"31364b00",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"43617274",
X"72696467",
X"65203332",
X"6b000000",
X"43617274",
X"72696467",
X"65203136",
X"6b206f6e",
X"65206368",
X"69700000",
X"43617274",
X"72696467",
X"65203136",
X"6b207477",
X"6f206368",
X"69700000",
X"45786974",
X"00000000",
X"61636964",
X"35323030",
X"2e726f6d",
X"00000000",
X"524f4d00",
X"42494e00",
X"43415200",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"00000000",
X"2f617461",
X"72353230",
X"302f726f",
X"6d000000",
X"2f617461",
X"72353230",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
