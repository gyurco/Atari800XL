
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81eb",
X"8c738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81f3",
X"f80c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757580f7",
X"a62d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7580f6e5",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80e0e004",
X"fd3d0d75",
X"705254ae",
X"aa3f83c0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"c0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83c0",
X"8008732e",
X"a13883c0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183c0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83c2d008",
X"248a38b4",
X"fb3fff0b",
X"83c2d00c",
X"800b83c0",
X"800c04ff",
X"3d0d7352",
X"83c0ac08",
X"722e8d38",
X"d93f7151",
X"96a03f71",
X"83c0ac0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"55805681",
X"54bc1508",
X"762e0981",
X"06819138",
X"7451c83f",
X"7958757a",
X"2580f738",
X"83c38008",
X"70892a57",
X"83ff0678",
X"84807231",
X"56565773",
X"78258338",
X"73557583",
X"c2d0082e",
X"8438ff82",
X"3f83c2d0",
X"088025a6",
X"3875892b",
X"5198dc3f",
X"83c38008",
X"8f3dfc11",
X"555c5481",
X"52f81b51",
X"96c63f76",
X"1483c380",
X"0c7583c2",
X"d00c7453",
X"76527851",
X"b3a53f83",
X"c0800883",
X"c3800816",
X"83c3800c",
X"78763176",
X"1b5b5956",
X"778024ff",
X"8b38617a",
X"710c5475",
X"5475802e",
X"83388154",
X"7383c080",
X"0c8e3d0d",
X"04fc3d0d",
X"fe943f76",
X"51fea83f",
X"863dfc05",
X"53785277",
X"5195e93f",
X"7975710c",
X"5483c080",
X"085483c0",
X"8008802e",
X"83388154",
X"7383c080",
X"0c863d0d",
X"04fe3d0d",
X"7583c2d0",
X"08535380",
X"72248938",
X"71732e84",
X"38fdcf3f",
X"7451fde3",
X"3f725197",
X"ae3f83c0",
X"80085283",
X"c0800880",
X"2e833881",
X"527183c0",
X"800c843d",
X"0d04803d",
X"0d7280c0",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"3d0d72bc",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"c40b83c0",
X"800c04fd",
X"3d0d7577",
X"71547053",
X"5553a9fb",
X"3f82c813",
X"08bc150c",
X"82c01308",
X"80c0150c",
X"fce43f73",
X"5193ab3f",
X"7383c0ac",
X"0c83c080",
X"085383c0",
X"8008802e",
X"83388153",
X"7283c080",
X"0c853d0d",
X"04fd3d0d",
X"75775553",
X"fcb83f72",
X"802ea538",
X"bc130852",
X"7351a985",
X"3f83c080",
X"088f3877",
X"527251ff",
X"9a3f83c0",
X"8008538a",
X"3982cc13",
X"0853d839",
X"81537283",
X"c0800c85",
X"3d0d04fe",
X"3d0dff0b",
X"83c2d00c",
X"7483c0b0",
X"0c7583c2",
X"cc0cafd9",
X"3f83c080",
X"0881ff06",
X"52815371",
X"993883c2",
X"e8518e94",
X"3f83c080",
X"085283c0",
X"8008802e",
X"83387252",
X"71537283",
X"c0800c84",
X"3d0d04fa",
X"3d0d787a",
X"82c41208",
X"82c41208",
X"70722459",
X"56565757",
X"73732e09",
X"81069138",
X"80c01652",
X"80c01751",
X"a6f63f83",
X"c0800855",
X"7483c080",
X"0c883d0d",
X"04f63d0d",
X"7c5b807b",
X"715c5457",
X"7a772e8c",
X"38811a82",
X"cc140854",
X"5a72f638",
X"805980d9",
X"397a5481",
X"5780707b",
X"7b315a57",
X"55ff1853",
X"74732580",
X"c13882cc",
X"14085273",
X"51ff8c3f",
X"800b83c0",
X"800825a1",
X"3882cc14",
X"0882cc11",
X"0882cc16",
X"0c7482cc",
X"120c5375",
X"802e8638",
X"7282cc17",
X"0c725480",
X"577382cc",
X"15088117",
X"575556ff",
X"b8398119",
X"59800bff",
X"1b545478",
X"73258338",
X"81547681",
X"32707506",
X"515372ff",
X"90388c3d",
X"0d04f73d",
X"0d7b7d5a",
X"5a82d052",
X"83c2cc08",
X"5180e5e1",
X"3f83c080",
X"0857f9da",
X"3f795283",
X"c2d45195",
X"b73f83c0",
X"80085480",
X"5383c080",
X"08732e09",
X"81068283",
X"3883c0b0",
X"080b0b81",
X"f0a85370",
X"5256a6b3",
X"3f0b0b81",
X"f0a85280",
X"c01651a6",
X"a63f75bc",
X"170c7382",
X"c0170c81",
X"0b82c417",
X"0c810b82",
X"c8170c73",
X"82cc170c",
X"ff1782d0",
X"17555781",
X"913983c0",
X"bc337082",
X"2a708106",
X"51545572",
X"81803874",
X"812a8106",
X"587780f6",
X"3874842a",
X"810682c4",
X"150c83c0",
X"bc338106",
X"82c8150c",
X"79527351",
X"a5cd3f73",
X"51a5e43f",
X"83c08008",
X"1453af73",
X"70810555",
X"3472bc15",
X"0c83c0bd",
X"527251a5",
X"ae3f83c0",
X"b40882c0",
X"150c83c0",
X"ca5280c0",
X"1451a59b",
X"3f78802e",
X"8d387351",
X"782d83c0",
X"8008802e",
X"99387782",
X"cc150c75",
X"802e8638",
X"7382cc17",
X"0c7382d0",
X"15ff1959",
X"55567680",
X"2e9b3883",
X"c0b45283",
X"c2d45194",
X"ad3f83c0",
X"80088a38",
X"83c0bd33",
X"5372fed2",
X"3878802e",
X"893883c0",
X"b00851fc",
X"b83f83c0",
X"b0085372",
X"83c0800c",
X"8b3d0d04",
X"ff3d0d80",
X"527351fd",
X"b53f833d",
X"0d04f03d",
X"0d627052",
X"54f6893f",
X"83c08008",
X"7453873d",
X"70535555",
X"f6a93ff7",
X"893f7351",
X"d33f6353",
X"745283c0",
X"800851fa",
X"b83f923d",
X"0d047183",
X"c0800c04",
X"80c01283",
X"c0800c04",
X"803d0d72",
X"82c01108",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"7282cc11",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d7282c4",
X"110883c0",
X"800c5182",
X"3d0d04f9",
X"3d0d7983",
X"c0900857",
X"57817727",
X"81963876",
X"88170827",
X"818e3875",
X"33557482",
X"2e893874",
X"832eb338",
X"80fe3974",
X"54761083",
X"fe065376",
X"882a8c17",
X"08055289",
X"3dfc0551",
X"aa873f83",
X"c0800880",
X"df38029d",
X"0533893d",
X"3371882b",
X"07565680",
X"d1398454",
X"76822b83",
X"fc065376",
X"872a8c17",
X"08055289",
X"3dfc0551",
X"a9d73f83",
X"c08008b0",
X"38029f05",
X"33028405",
X"9e053371",
X"982b7190",
X"2b07028c",
X"059d0533",
X"70882b72",
X"078d3d33",
X"7180ffff",
X"fe800607",
X"51525357",
X"58568339",
X"81557483",
X"c0800c89",
X"3d0d04fb",
X"3d0d83c0",
X"9008fe19",
X"881208fe",
X"05555654",
X"80567473",
X"278d3882",
X"14337571",
X"29941608",
X"05575375",
X"83c0800c",
X"873d0d04",
X"fc3d0d76",
X"52800b83",
X"c0900870",
X"33515253",
X"70832e09",
X"81069138",
X"95123394",
X"13337198",
X"2b71902b",
X"07555551",
X"9b12339a",
X"13337188",
X"2b077407",
X"83c0800c",
X"55863d0d",
X"04fc3d0d",
X"7683c090",
X"08555580",
X"75238815",
X"08537281",
X"2e883888",
X"14087326",
X"85388152",
X"b2397290",
X"38733352",
X"71832e09",
X"81068538",
X"90140853",
X"728c160c",
X"72802e8d",
X"387251fe",
X"d63f83c0",
X"80085285",
X"39901408",
X"52719016",
X"0c805271",
X"83c0800c",
X"863d0d04",
X"fa3d0d78",
X"83c09008",
X"71228105",
X"7083ffff",
X"06575457",
X"5573802e",
X"88389015",
X"08537286",
X"38835280",
X"e739738f",
X"06527180",
X"da388113",
X"90160c8c",
X"15085372",
X"9038830b",
X"84172257",
X"52737627",
X"80c638bf",
X"39821633",
X"ff057484",
X"2a065271",
X"b2387251",
X"fcb13f81",
X"527183c0",
X"800827a8",
X"38835283",
X"c0800888",
X"1708279c",
X"3883c080",
X"088c160c",
X"83c08008",
X"51fdbc3f",
X"83c08008",
X"90160c73",
X"75238052",
X"7183c080",
X"0c883d0d",
X"04f23d0d",
X"60626458",
X"5e5b7533",
X"5574a02e",
X"09810688",
X"38811670",
X"4456ef39",
X"62703356",
X"5674af2e",
X"09810684",
X"38811643",
X"800b881c",
X"0c627033",
X"5155749f",
X"2691387a",
X"51fdd23f",
X"83c08008",
X"56807d34",
X"83813993",
X"3d841c08",
X"7058595f",
X"8a55a076",
X"70810558",
X"34ff1555",
X"74ff2e09",
X"8106ef38",
X"80705a5c",
X"887f085f",
X"5a7b811d",
X"7081ff06",
X"60137033",
X"70af3270",
X"30a07327",
X"71802507",
X"5151525b",
X"535e5755",
X"7480e738",
X"76ae2e09",
X"81068338",
X"8155787a",
X"27750755",
X"74802e9f",
X"38798832",
X"703078ae",
X"32703070",
X"73079f2a",
X"53515751",
X"5675bb38",
X"88598b5a",
X"ffab3976",
X"982b5574",
X"80258738",
X"81ea9c17",
X"3357ff9f",
X"17557499",
X"268938e0",
X"177081ff",
X"06585578",
X"811a7081",
X"ff06721b",
X"535b5755",
X"767534fe",
X"f8397b1e",
X"7f0c8055",
X"76a02683",
X"38815574",
X"8b19347a",
X"51fc823f",
X"83c08008",
X"80f538a0",
X"547a2270",
X"852b83e0",
X"06545590",
X"1b08527c",
X"51a4923f",
X"83c08008",
X"5783c080",
X"08818138",
X"7c335574",
X"802e80f4",
X"388b1d33",
X"70832a70",
X"81065156",
X"5674b438",
X"8b7d841d",
X"0883c080",
X"08595b5b",
X"58ff1858",
X"77ff2e9a",
X"38797081",
X"055b3379",
X"7081055b",
X"33717131",
X"52565675",
X"802ee238",
X"86397580",
X"2e96387a",
X"51fbe53f",
X"ff863983",
X"c0800856",
X"83c08008",
X"b6388339",
X"7656841b",
X"088b1133",
X"515574a7",
X"388b1d33",
X"70842a70",
X"81065156",
X"56748938",
X"83569439",
X"81569039",
X"7c51fa94",
X"3f83c080",
X"08881c0c",
X"fd813975",
X"83c0800c",
X"903d0d04",
X"f83d0d7a",
X"7c595782",
X"5483fe53",
X"77527651",
X"a2d73f83",
X"5683c080",
X"0880ec38",
X"81173377",
X"3371882b",
X"07565682",
X"567482d4",
X"d52e0981",
X"0680d438",
X"7554b653",
X"77527651",
X"a2ab3f83",
X"c0800898",
X"38811733",
X"77337188",
X"2b0783c0",
X"80085256",
X"56748182",
X"c62eac38",
X"825480d2",
X"53775276",
X"51a2823f",
X"83c08008",
X"98388117",
X"33773371",
X"882b0783",
X"c0800852",
X"56567481",
X"82c62e83",
X"38815675",
X"83c0800c",
X"8a3d0d04",
X"eb3d0d67",
X"5a800b83",
X"c0900ca1",
X"a43f83c0",
X"80088106",
X"55825674",
X"83ef3874",
X"75538f3d",
X"70535759",
X"feca3f83",
X"c0800881",
X"ff065776",
X"812e0981",
X"0680d438",
X"905483be",
X"53745275",
X"51a1963f",
X"83c08008",
X"80c9388f",
X"3d335574",
X"802e80c9",
X"3802bf05",
X"33028405",
X"be053371",
X"982b7190",
X"2b07028c",
X"05bd0533",
X"70882b72",
X"07953d33",
X"71077058",
X"7b575e52",
X"5e575957",
X"fdee3f83",
X"c0800881",
X"ff065776",
X"832e0981",
X"06863881",
X"5682f239",
X"76802e86",
X"38865682",
X"e839a454",
X"8d537852",
X"7551a0ad",
X"3f815683",
X"c0800882",
X"d43802be",
X"05330284",
X"05bd0533",
X"71882b07",
X"595d77ab",
X"380280ce",
X"05330284",
X"0580cd05",
X"3371982b",
X"71902b07",
X"973d3370",
X"882b7207",
X"02940580",
X"cb053371",
X"0754525e",
X"57595602",
X"b7053378",
X"71290288",
X"05b60533",
X"028c05b5",
X"05337188",
X"2b07701d",
X"707f8c05",
X"0c5f5957",
X"595d8e3d",
X"33821b34",
X"02b90533",
X"903d3371",
X"882b075a",
X"5c78841b",
X"2302bb05",
X"33028405",
X"ba053371",
X"882b0756",
X"5c74ab38",
X"0280ca05",
X"33028405",
X"80c90533",
X"71982b71",
X"902b0796",
X"3d337088",
X"2b720702",
X"940580c7",
X"05337107",
X"51525357",
X"5e5c7476",
X"31783179",
X"842a903d",
X"33547171",
X"31535656",
X"80d6c63f",
X"83c08008",
X"82057088",
X"1c0c83c0",
X"8008e08a",
X"05565674",
X"83dffe26",
X"83388257",
X"83fff676",
X"27853883",
X"57893986",
X"5676802e",
X"80db3876",
X"7a347683",
X"2e098106",
X"b0380280",
X"d6053302",
X"840580d5",
X"05337198",
X"2b71902b",
X"07993d33",
X"70882b72",
X"07029405",
X"80d30533",
X"71077f90",
X"050c525e",
X"57585686",
X"39771b90",
X"1b0c841a",
X"228c1b08",
X"1971842a",
X"05941c0c",
X"5d800b81",
X"1b347983",
X"c0900c80",
X"567583c0",
X"800c973d",
X"0d04e93d",
X"0d83c090",
X"08568554",
X"75802e81",
X"8238800b",
X"81173499",
X"3de01146",
X"6a548a3d",
X"705458ec",
X"0551f6e5",
X"3f83c080",
X"085483c0",
X"800880df",
X"38893d33",
X"5473802e",
X"913802ab",
X"05337084",
X"2a810651",
X"5574802e",
X"86388354",
X"80c13976",
X"51f4893f",
X"83c08008",
X"a0170c02",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"9c1c0c52",
X"78981b0c",
X"53565957",
X"810b8117",
X"34745473",
X"83c0800c",
X"993d0d04",
X"f53d0d7d",
X"7f617283",
X"c090085a",
X"5d5d595c",
X"807b0c85",
X"5775802e",
X"81e03881",
X"16338106",
X"55845774",
X"802e81d2",
X"38913974",
X"81173486",
X"39800b81",
X"17348157",
X"81c0399c",
X"16089817",
X"08315574",
X"78278338",
X"74587780",
X"2e81a938",
X"98160870",
X"83ff0656",
X"577480cf",
X"38821633",
X"ff057789",
X"2a067081",
X"ff065a55",
X"78a03876",
X"8738a016",
X"08558d39",
X"a4160851",
X"f0e93f83",
X"c0800855",
X"817527ff",
X"a83874a4",
X"170ca416",
X"0851f283",
X"3f83c080",
X"085583c0",
X"8008802e",
X"ff893883",
X"c0800819",
X"a8170c98",
X"160883ff",
X"06848071",
X"31515577",
X"75278338",
X"77557483",
X"ffff0654",
X"98160883",
X"ff0653a8",
X"16085279",
X"577b8338",
X"7b577651",
X"9ad33f83",
X"c08008fe",
X"d0389816",
X"08159817",
X"0c741a78",
X"76317c08",
X"177d0c59",
X"5afed339",
X"80577683",
X"c0800c8d",
X"3d0d04fa",
X"3d0d7883",
X"c0900855",
X"56855573",
X"802e81e3",
X"38811433",
X"81065384",
X"5572802e",
X"81d5389c",
X"14085372",
X"76278338",
X"72569814",
X"0857800b",
X"98150c75",
X"802e81b9",
X"38821433",
X"70892b56",
X"5376802e",
X"b7387452",
X"ff165180",
X"d1c73f83",
X"c08008ff",
X"18765470",
X"53585380",
X"d1b73f83",
X"c0800873",
X"26963874",
X"30707806",
X"7098170c",
X"777131a4",
X"17085258",
X"51538939",
X"a0140870",
X"a4160c53",
X"747627b9",
X"387251ee",
X"d63f83c0",
X"80085381",
X"0b83c080",
X"08278b38",
X"88140883",
X"c0800826",
X"8838800b",
X"811534b0",
X"3983c080",
X"08a4150c",
X"98140815",
X"98150c75",
X"753156c4",
X"39981408",
X"16709816",
X"0c735256",
X"efc53f83",
X"c080088c",
X"3883c080",
X"08811534",
X"81559439",
X"821433ff",
X"0576892a",
X"0683c080",
X"0805a815",
X"0c805574",
X"83c0800c",
X"883d0d04",
X"ef3d0d63",
X"56855583",
X"c0900880",
X"2e80d238",
X"933df405",
X"84170c64",
X"53883d70",
X"53765257",
X"f1cf3f83",
X"c0800855",
X"83c08008",
X"b438883d",
X"33547380",
X"2ea13802",
X"a7053370",
X"842a7081",
X"06515555",
X"83557380",
X"2e973876",
X"51eef53f",
X"83c08008",
X"88170c75",
X"51efa63f",
X"83c08008",
X"557483c0",
X"800c933d",
X"0d04e43d",
X"0d6ea13d",
X"08405e85",
X"5683c090",
X"08802e84",
X"85389e3d",
X"f405841f",
X"0c7e9838",
X"7d51eef5",
X"3f83c080",
X"085683ee",
X"39814181",
X"f6398341",
X"81f13993",
X"3d7f9605",
X"4159807f",
X"8295055e",
X"56756081",
X"ff053483",
X"41901e08",
X"762e81d3",
X"38a0547d",
X"2270852b",
X"83e00654",
X"58901e08",
X"52785196",
X"dc3f83c0",
X"80084183",
X"c08008ff",
X"b8387833",
X"5c7b802e",
X"ffb4388b",
X"193370bf",
X"06718106",
X"52435574",
X"802e80de",
X"387b81bf",
X"0655748f",
X"2480d338",
X"9a193355",
X"7480cb38",
X"f31d7058",
X"5d815675",
X"8b2e0981",
X"0685388e",
X"568b3975",
X"9a2e0981",
X"0683389c",
X"56751970",
X"70810552",
X"33713381",
X"1a821a5f",
X"5b525b55",
X"74863879",
X"77348539",
X"80df7734",
X"777b5757",
X"7aa02e09",
X"8106c038",
X"81567b81",
X"e5327030",
X"709f2a51",
X"51557bae",
X"2e933874",
X"802e8e38",
X"61832a70",
X"81065155",
X"74802e97",
X"387d51ed",
X"df3f83c0",
X"80084183",
X"c0800887",
X"38901e08",
X"feaf3880",
X"60347580",
X"2e88387c",
X"527f518e",
X"823f6080",
X"2e863880",
X"0b901f0c",
X"60566083",
X"2e853860",
X"81d03889",
X"1f57901e",
X"08802e81",
X"a8388056",
X"75197033",
X"515574a0",
X"2ea03874",
X"852e0981",
X"06843881",
X"e5557477",
X"70810559",
X"34811670",
X"81ff0657",
X"55877627",
X"d7388819",
X"335574a0",
X"2ea938ae",
X"77708105",
X"59348856",
X"75197033",
X"515574a0",
X"2e953874",
X"77708105",
X"59348116",
X"7081ff06",
X"57558a76",
X"27e2388b",
X"19337f88",
X"05349f19",
X"339e1a33",
X"71982b71",
X"902b079d",
X"1c337088",
X"2b72079c",
X"1e337107",
X"640c5299",
X"1d33981e",
X"3371882b",
X"07535153",
X"57595674",
X"7f840523",
X"97193396",
X"1a337188",
X"2b075656",
X"747f8605",
X"23807734",
X"7d51ebf0",
X"3f83c080",
X"08833270",
X"30707207",
X"9f2c83c0",
X"80080652",
X"5656961f",
X"3355748a",
X"38891f52",
X"961f518c",
X"8e3f7583",
X"c0800c9e",
X"3d0d04f4",
X"3d0d7e8f",
X"3dec1156",
X"56589053",
X"f0155277",
X"51e0d23f",
X"83c08008",
X"80d63878",
X"902e0981",
X"0680cd38",
X"02ab0533",
X"81f4800b",
X"81f48033",
X"5758568c",
X"3974762e",
X"8a388417",
X"70335657",
X"74f33876",
X"33705755",
X"74802eac",
X"38821722",
X"708a2b90",
X"3dec0556",
X"70555656",
X"96800a52",
X"7751e081",
X"3f83c080",
X"08863878",
X"752e8538",
X"80568539",
X"81173356",
X"7583c080",
X"0c8e3d0d",
X"04fc3d0d",
X"76705255",
X"8b953f83",
X"c0800815",
X"ff055473",
X"752e8e38",
X"73335372",
X"ae2e8638",
X"ff1454ef",
X"39775281",
X"14518aad",
X"3f83c080",
X"08307083",
X"c0800807",
X"802583c0",
X"800c5386",
X"3d0d04fc",
X"3d0d7670",
X"5255e6ee",
X"3f83c080",
X"08548153",
X"83c08008",
X"80c13874",
X"51e6b13f",
X"83c08008",
X"81f0b853",
X"83c08008",
X"5253ff91",
X"3f83c080",
X"08a13881",
X"f0bc5272",
X"51ff823f",
X"83c08008",
X"923881f0",
X"c0527251",
X"fef33f83",
X"c0800880",
X"2e833881",
X"54735372",
X"83c0800c",
X"863d0d04",
X"fd3d0d75",
X"705254e6",
X"8d3f8153",
X"83c08008",
X"98387351",
X"e5d63f83",
X"c3980852",
X"83c08008",
X"51feba3f",
X"83c08008",
X"537283c0",
X"800c853d",
X"0d04df3d",
X"0da43d08",
X"70525edb",
X"f43f83c0",
X"80083395",
X"3d565473",
X"963881f7",
X"c8527451",
X"898d3f9a",
X"397d5278",
X"51defc3f",
X"84d0397d",
X"51dbda3f",
X"83c08008",
X"527451db",
X"8a3f8043",
X"80428041",
X"804083c3",
X"a0085294",
X"3d70525d",
X"e1e43f83",
X"c0800859",
X"800b83c0",
X"8008555b",
X"83c08008",
X"7b2e9438",
X"811b7452",
X"5be4e63f",
X"83c08008",
X"5483c080",
X"08ee3880",
X"5aff5f79",
X"09709f2c",
X"7b065b54",
X"7a7a2484",
X"38ff1b5a",
X"f61a7009",
X"709f2c72",
X"067bff12",
X"5a5a5255",
X"55807525",
X"95387651",
X"e4ab3f83",
X"c0800876",
X"ff185855",
X"57738024",
X"ed38747f",
X"2e8638a1",
X"b53f745f",
X"78ff1b70",
X"585d5880",
X"7a259538",
X"7751e481",
X"3f83c080",
X"0876ff18",
X"58555873",
X"8024ed38",
X"800b83c7",
X"d00c800b",
X"83c8980c",
X"81f0c451",
X"8d8c3f81",
X"800b83c8",
X"980c81f0",
X"cc518cfe",
X"3fa80b83",
X"c7d00c76",
X"802e80e4",
X"3883c7d0",
X"08777932",
X"70307072",
X"07802570",
X"872b83c8",
X"980c5156",
X"78535656",
X"e3b83f83",
X"c0800880",
X"2e883881",
X"f0d4518c",
X"c53f7651",
X"e2fa3f83",
X"c0800852",
X"81f2b451",
X"8cb43f76",
X"51e3823f",
X"83c08008",
X"83c7d008",
X"55577574",
X"258638a8",
X"1656f739",
X"7583c7d0",
X"0c86f076",
X"24ff9838",
X"87980b83",
X"c7d00c77",
X"802eb138",
X"7751e2b8",
X"3f83c080",
X"08785255",
X"e2d83f81",
X"f0dc5483",
X"c080088d",
X"38873980",
X"763481d0",
X"3981f0d8",
X"54745373",
X"5281f0ac",
X"518bd33f",
X"805481f0",
X"b4518bca",
X"3f811454",
X"73a82e09",
X"8106ef38",
X"868da051",
X"9da83f80",
X"52903d70",
X"525780c7",
X"bc3f8352",
X"765180c7",
X"b43f6281",
X"8f386180",
X"2e80fb38",
X"7b5473ff",
X"2e963878",
X"802e818a",
X"387851e1",
X"dc3f83c0",
X"8008ff15",
X"5559e739",
X"78802e80",
X"f5387851",
X"e1d83f83",
X"c0800880",
X"2efc8e38",
X"7851e1a0",
X"3f83c080",
X"085281f0",
X"a85183e0",
X"3f83c080",
X"08a3387c",
X"5185983f",
X"83c08008",
X"5574ff16",
X"56548074",
X"25ae3874",
X"1d703355",
X"5673af2e",
X"fecd38e9",
X"397851e0",
X"e13f83c0",
X"8008527c",
X"5184d03f",
X"8f397f88",
X"29601005",
X"7a056105",
X"5afc9039",
X"62802efb",
X"d1388052",
X"765180c6",
X"943fa33d",
X"0d04803d",
X"0d9088b8",
X"337081ff",
X"0670842a",
X"81327081",
X"06515151",
X"5170802e",
X"8d38a80b",
X"9088b834",
X"b80b9088",
X"b8347083",
X"c0800c82",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067085",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d3898",
X"0b9088b8",
X"34b80b90",
X"88b83470",
X"83c0800c",
X"823d0d04",
X"930b9088",
X"bc34ff0b",
X"9088a834",
X"04ff3d0d",
X"028f0533",
X"52800b90",
X"88bc348a",
X"519aef3f",
X"df3f80f8",
X"0b9088a0",
X"34800b90",
X"888834fa",
X"12527190",
X"88803480",
X"0b908898",
X"34719088",
X"90349088",
X"b8528072",
X"34b87234",
X"833d0d04",
X"803d0d02",
X"8b053351",
X"709088b4",
X"34febf3f",
X"83c08008",
X"802ef638",
X"823d0d04",
X"803d0d84",
X"39a8de3f",
X"fed93f83",
X"c0800880",
X"2ef33890",
X"88b43370",
X"81ff0683",
X"c0800c51",
X"823d0d04",
X"803d0da3",
X"0b9088bc",
X"34ff0b90",
X"88a83490",
X"88b851a8",
X"7134b871",
X"34823d0d",
X"04803d0d",
X"9088bc33",
X"70982b70",
X"802583c0",
X"800c5151",
X"823d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"832a8132",
X"70810651",
X"51515170",
X"802ee838",
X"b00b9088",
X"b834b80b",
X"9088b834",
X"823d0d04",
X"803d0d90",
X"80ac0881",
X"0683c080",
X"0c823d0d",
X"04fd3d0d",
X"75775454",
X"80732594",
X"38737081",
X"05553352",
X"81f0e051",
X"87843fff",
X"1353e939",
X"853d0d04",
X"fd3d0d75",
X"77535473",
X"33517089",
X"38713351",
X"70802ea1",
X"38733372",
X"33525372",
X"71278538",
X"ff519439",
X"70732785",
X"3881518b",
X"39811481",
X"135354d3",
X"39805170",
X"83c0800c",
X"853d0d04",
X"fd3d0d75",
X"77545472",
X"337081ff",
X"06525270",
X"802ea338",
X"7181ff06",
X"8114ffbf",
X"12535452",
X"70992689",
X"38a01270",
X"81ff0653",
X"51717470",
X"81055634",
X"d2398074",
X"34853d0d",
X"04ffbd3d",
X"0d80c63d",
X"0852a53d",
X"705254ff",
X"b33f80c7",
X"3d085285",
X"3d705253",
X"ffa63f72",
X"527351fe",
X"df3f80c5",
X"3d0d04fe",
X"3d0d7476",
X"53537170",
X"81055333",
X"51707370",
X"81055534",
X"70f03884",
X"3d0d04fe",
X"3d0d7452",
X"80723352",
X"5370732e",
X"8d388112",
X"81147133",
X"53545270",
X"f5387283",
X"c0800c84",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"be9f3f83",
X"c080087a",
X"27ee3874",
X"802e80dd",
X"38745275",
X"51be8a3f",
X"83c08008",
X"75537652",
X"54be8e3f",
X"83c08008",
X"7a537552",
X"56bdf23f",
X"83c08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"c08008c5",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9f",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fc813f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd53f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbb13f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83c0940c",
X"7183c098",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383c094",
X"085283c0",
X"980851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"bdbe5351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fc3d",
X"0d765574",
X"83c3ac08",
X"2eaf3880",
X"53745187",
X"c13f83c0",
X"800881ff",
X"06ff1470",
X"81ff0672",
X"30709f2a",
X"51525553",
X"5472802e",
X"843871dd",
X"3873fe38",
X"7483c3ac",
X"0c863d0d",
X"04ff3d0d",
X"ff0b83c3",
X"ac0c84a5",
X"3f815187",
X"853f83c0",
X"800881ff",
X"065271ee",
X"3881d33f",
X"7183c080",
X"0c833d0d",
X"04fc3d0d",
X"76028405",
X"a2052202",
X"8805a605",
X"227a5455",
X"5555ff82",
X"3f72802e",
X"a03883c3",
X"c0143375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552dd",
X"39800b83",
X"c0800c86",
X"3d0d04fc",
X"3d0d7678",
X"7a115653",
X"55805371",
X"742e9338",
X"72155170",
X"3383c3c0",
X"13348112",
X"81145452",
X"ea39800b",
X"83c0800c",
X"863d0d04",
X"fd3d0d90",
X"5483c3ac",
X"085186f4",
X"3f83c080",
X"0881ff06",
X"ff157130",
X"71307073",
X"079f2a72",
X"9f2a0652",
X"55525553",
X"72db3885",
X"3d0d0480",
X"3d0d83c3",
X"b8081083",
X"c3b00807",
X"9080a80c",
X"823d0d04",
X"800b83c3",
X"b80ce43f",
X"04810b83",
X"c3b80cdb",
X"3f04ed3f",
X"047183c3",
X"b40c0480",
X"3d0d8051",
X"f43f810b",
X"83c3b80c",
X"810b83c3",
X"b00cffbb",
X"3f823d0d",
X"04803d0d",
X"72307074",
X"07802583",
X"c3b00c51",
X"ffa53f82",
X"3d0d0480",
X"3d0d028b",
X"05339080",
X"a40c9080",
X"a8087081",
X"06515170",
X"f5389080",
X"a4087081",
X"ff0683c0",
X"800c5182",
X"3d0d0480",
X"3d0d81ff",
X"51d13f83",
X"c0800881",
X"ff0683c0",
X"800c823d",
X"0d04803d",
X"0d73902b",
X"73079080",
X"b40c823d",
X"0d0404fb",
X"3d0d7802",
X"84059f05",
X"3370982b",
X"55575572",
X"80259b38",
X"7580ff06",
X"56805280",
X"f751e03f",
X"83c08008",
X"81ff0654",
X"73812680",
X"ff388051",
X"fee73fff",
X"a23f8151",
X"fedf3fff",
X"9a3f7551",
X"feed3f74",
X"982a51fe",
X"e63f7490",
X"2a7081ff",
X"065253fe",
X"da3f7488",
X"2a7081ff",
X"065253fe",
X"ce3f7481",
X"ff0651fe",
X"c63f8155",
X"7580c02e",
X"09810686",
X"38819555",
X"8d397580",
X"c82e0981",
X"06843881",
X"87557451",
X"fea53f8a",
X"55fec83f",
X"83c08008",
X"81ff0670",
X"982b5454",
X"7280258c",
X"38ff1570",
X"81ff0656",
X"5374e238",
X"7383c080",
X"0c873d0d",
X"04fa3d0d",
X"fdc53f80",
X"51fdda3f",
X"8a54fe93",
X"3fff1470",
X"81ff0655",
X"5373f338",
X"73745355",
X"80c051fe",
X"a63f83c0",
X"800881ff",
X"06547381",
X"2e098106",
X"829f3883",
X"aa5280c8",
X"51fe8c3f",
X"83c08008",
X"81ff0653",
X"72812e09",
X"810681a8",
X"38745487",
X"3d741154",
X"56fdc83f",
X"83c08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e53802",
X"9a053353",
X"72812e09",
X"810681d9",
X"38029b05",
X"335380ce",
X"90547281",
X"aa2e8d38",
X"81c73980",
X"e4518b9a",
X"3fff1454",
X"73802e81",
X"b838820a",
X"5281e951",
X"fda53f83",
X"c0800881",
X"ff065372",
X"de387252",
X"80fa51fd",
X"923f83c0",
X"800881ff",
X"06537281",
X"90387254",
X"731653fc",
X"d63f83c0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e8",
X"38873d33",
X"70862a70",
X"81065154",
X"548c5572",
X"80e33884",
X"5580de39",
X"745281e9",
X"51fccc3f",
X"83c08008",
X"81ff0653",
X"825581e9",
X"56817327",
X"86387355",
X"80c15680",
X"ce90548a",
X"3980e451",
X"8a8c3fff",
X"14547380",
X"2ea93880",
X"527551fc",
X"9a3f83c0",
X"800881ff",
X"065372e1",
X"38848052",
X"80d051fc",
X"863f83c0",
X"800881ff",
X"06537280",
X"2e833880",
X"557483c3",
X"bc348051",
X"fb873ffb",
X"c23f883d",
X"0d04fb3d",
X"0d775480",
X"0b83c3bc",
X"3370832a",
X"70810651",
X"55575572",
X"752e0981",
X"06853873",
X"892b5473",
X"5280d151",
X"fbbd3f83",
X"c0800881",
X"ff065372",
X"bd3882b8",
X"c054fb83",
X"3f83c080",
X"0881ff06",
X"537281ff",
X"2e098106",
X"8938ff14",
X"5473e738",
X"9f397281",
X"fe2e0981",
X"06963883",
X"c7c05283",
X"c3c051fa",
X"ed3ffad3",
X"3ffad03f",
X"83398155",
X"8051fa89",
X"3ffac43f",
X"7481ff06",
X"83c0800c",
X"873d0d04",
X"fb3d0d77",
X"83c3c056",
X"548151f9",
X"ec3f83c3",
X"bc337083",
X"2a708106",
X"51545672",
X"85387389",
X"2b547352",
X"80d851fa",
X"b63f83c0",
X"800881ff",
X"06537280",
X"e43881ff",
X"51f9d43f",
X"81fe51f9",
X"ce3f8480",
X"53747081",
X"05563351",
X"f9c13fff",
X"137083ff",
X"ff065153",
X"72eb3872",
X"51f9b03f",
X"7251f9ab",
X"3ff9d03f",
X"83c08008",
X"9f0653a7",
X"88547285",
X"2e8c3899",
X"3980e451",
X"87c43fff",
X"1454f9b3",
X"3f83c080",
X"0881ff2e",
X"843873e9",
X"388051f8",
X"e43ff99f",
X"3f800b83",
X"c0800c87",
X"3d0d0471",
X"83c7c40c",
X"8880800b",
X"83c7c00c",
X"8480800b",
X"83c7c80c",
X"04fd3d0d",
X"77701755",
X"7705ff1a",
X"535371ff",
X"2e943873",
X"70810555",
X"33517073",
X"70810555",
X"34ff1252",
X"e939853d",
X"0d04fb3d",
X"0d87a681",
X"0b83c7c4",
X"08565675",
X"3383a680",
X"1634a054",
X"83a08053",
X"83c7c408",
X"5283c7c0",
X"0851ffb1",
X"3fa05483",
X"a4805383",
X"c7c40852",
X"83c7c008",
X"51ff9e3f",
X"905483a8",
X"805383c7",
X"c4085283",
X"c7c00851",
X"ff8b3fa0",
X"53805283",
X"c7c80883",
X"a0800551",
X"86953fa0",
X"53805283",
X"c7c80883",
X"a4800551",
X"86853f90",
X"53805283",
X"c7c80883",
X"a8800551",
X"85f53fff",
X"763483a0",
X"80548053",
X"83c7c408",
X"5283c7c8",
X"0851fec5",
X"3f80d080",
X"5483b080",
X"5383c7c4",
X"085283c7",
X"c80851fe",
X"b03f87ba",
X"3fa25480",
X"5383c7c8",
X"088c8005",
X"5281f4f4",
X"51fe9a3f",
X"860b87a8",
X"8334800b",
X"87a88234",
X"800b87a0",
X"9a34af0b",
X"87a09634",
X"bf0b87a0",
X"9734800b",
X"87a09834",
X"9f0b87a0",
X"9934800b",
X"87a09b34",
X"e00b87a8",
X"8934a20b",
X"87a88034",
X"830b87a4",
X"8f34820b",
X"87a88134",
X"873d0d04",
X"fc3d0d83",
X"a0805480",
X"5383c7c8",
X"085283c7",
X"c40851fd",
X"b83f80d0",
X"805483b0",
X"805383c7",
X"c8085283",
X"c7c40851",
X"fda33fa0",
X"5483a080",
X"5383c7c8",
X"085283c7",
X"c40851fd",
X"903fa054",
X"83a48053",
X"83c7c808",
X"5283c7c4",
X"0851fcfd",
X"3f905483",
X"a8805383",
X"c7c80852",
X"83c7c408",
X"51fcea3f",
X"83c7c408",
X"5583a680",
X"153387a6",
X"8134863d",
X"0d04fa3d",
X"0d787052",
X"55c1e33f",
X"83ffff0b",
X"83c08008",
X"25a93874",
X"51c1e43f",
X"83c08008",
X"9e3883c0",
X"80085788",
X"3dfc0554",
X"84808053",
X"83c7c408",
X"527451ff",
X"bf963fff",
X"bedc3f88",
X"3d0d04fa",
X"3d0d7870",
X"5255c1a2",
X"3f83ffff",
X"0b83c080",
X"08259638",
X"8057883d",
X"fc055484",
X"80805383",
X"c7c40852",
X"7451c095",
X"3f883d0d",
X"04803d0d",
X"90809008",
X"810683c0",
X"800c823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087081",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fd0676",
X"1007720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870822c",
X"bf0683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe830676",
X"822b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087088",
X"2c870683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f1ff06",
X"76882b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"912cbf06",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fc87",
X"ffff0676",
X"912b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087099",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70ffbf0a",
X"0676992b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90808008",
X"70882c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"0870892c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708a",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8b2c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708c2cbf",
X"0683c080",
X"0c51823d",
X"0d04fe3d",
X"0d7481e6",
X"29872a90",
X"80a00c84",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70810554",
X"34ff1151",
X"f039843d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"8405540c",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"84808053",
X"80528880",
X"0a51ffb3",
X"3f818080",
X"53805282",
X"800a51c6",
X"3f843d0d",
X"04803d0d",
X"8151fcaa",
X"3f72802e",
X"90388051",
X"fdfe3fcd",
X"3f83c7cc",
X"3351fdf4",
X"3f8151fc",
X"bb3f8051",
X"fcb63f80",
X"51fc873f",
X"823d0d04",
X"fd3d0d75",
X"52805480",
X"ff722588",
X"38810bff",
X"80135354",
X"ffbf1251",
X"70992686",
X"38e01252",
X"b039ff9f",
X"12519971",
X"27a738d0",
X"12e01354",
X"51708926",
X"85387252",
X"9839728f",
X"26853872",
X"528f3971",
X"ba2e0981",
X"0685389a",
X"52833980",
X"5273802e",
X"85388180",
X"12527181",
X"ff0683c0",
X"800c853d",
X"0d04803d",
X"0d84d8c0",
X"51807170",
X"81055334",
X"7084e0c0",
X"2e098106",
X"f038823d",
X"0d04fe3d",
X"0d029705",
X"3351fef4",
X"3f83c080",
X"0881ff06",
X"83c7d008",
X"54528073",
X"249b3883",
X"c8940813",
X"7283c898",
X"08075353",
X"71733483",
X"c7d00881",
X"0583c7d0",
X"0c843d0d",
X"04fa3d0d",
X"82800a1b",
X"55805788",
X"3dfc0554",
X"79537452",
X"7851ffba",
X"ac3f883d",
X"0d04fe3d",
X"0d83c7e8",
X"08527451",
X"c1903f83",
X"c080088c",
X"38765375",
X"5283c7e8",
X"0851c63f",
X"843d0d04",
X"fe3d0d83",
X"c7e80853",
X"75527451",
X"ffbbce3f",
X"83c08008",
X"8d387753",
X"765283c7",
X"e80851ff",
X"a03f843d",
X"0d04f73d",
X"0daabd3f",
X"83c08008",
X"81ff06ff",
X"05577683",
X"38815780",
X"feff3f83",
X"c0800883",
X"c0800856",
X"5a871533",
X"5473802e",
X"80df3874",
X"0881ecc8",
X"2e098106",
X"80d33880",
X"0b911633",
X"55597379",
X"2e80c638",
X"74569a16",
X"33547383",
X"2e098106",
X"a438a416",
X"70335558",
X"80527351",
X"a8a73f80",
X"53805273",
X"51a8c73f",
X"81145476",
X"74258338",
X"80547378",
X"34811980",
X"d8179117",
X"33565759",
X"78742e09",
X"8106ffbe",
X"3881c415",
X"98c01b55",
X"5574742e",
X"098106ff",
X"88388b3d",
X"0d04f63d",
X"0d80fdf1",
X"3f83c080",
X"087d83c0",
X"80085859",
X"5b7783c7",
X"d00c8716",
X"33557480",
X"2e81a738",
X"75085473",
X"81f0802e",
X"09810693",
X"38901633",
X"53871633",
X"5281f0e8",
X"51e8f33f",
X"81883973",
X"81ecc82e",
X"09810680",
X"fd387452",
X"81f0fc51",
X"e8dc3f80",
X"70911833",
X"565b5973",
X"792e80e6",
X"38a41657",
X"f6173355",
X"79802e91",
X"38ff1554",
X"73822689",
X"38a81870",
X"83c7d00c",
X"5874812e",
X"09810687",
X"3881f184",
X"518d3974",
X"822e0981",
X"068a3881",
X"f18c51e8",
X"953f9539",
X"74832e09",
X"81068f38",
X"76338105",
X"5281f198",
X"51e7ff3f",
X"815a8119",
X"80d81891",
X"18335658",
X"5978742e",
X"098106ff",
X"9f38a818",
X"81c41798",
X"c01d5657",
X"5875742e",
X"098106fe",
X"b8388c3d",
X"0d04fe3d",
X"0d83c7e8",
X"0851ffb7",
X"c13f83c0",
X"80088180",
X"802e0981",
X"06883883",
X"c1808053",
X"9c3983c7",
X"e80851ff",
X"b7a43f83",
X"c0800880",
X"d0802e09",
X"81069338",
X"83c1b080",
X"5383c080",
X"085283c7",
X"e80851fb",
X"d43f843d",
X"0d04803d",
X"0df6fc3f",
X"83c08008",
X"842981f5",
X"98057008",
X"83c0800c",
X"51823d0d",
X"04ed3d0d",
X"80448043",
X"80428041",
X"80705a5b",
X"facc3f80",
X"0b83c7d0",
X"0c800b83",
X"c8980c81",
X"f1ec51e6",
X"c53f8180",
X"0b83c898",
X"0c81f1f0",
X"51e6b73f",
X"80d00b83",
X"c7d00c78",
X"30707a07",
X"80257087",
X"2b83c898",
X"0c5155f5",
X"ed3f83c0",
X"80085281",
X"f1f851e6",
X"913f80f8",
X"0b83c7d0",
X"0c788132",
X"70307072",
X"07802570",
X"872b83c8",
X"980c5156",
X"569eb03f",
X"83c08008",
X"5281f288",
X"51e5e73f",
X"81a00b83",
X"c7d00c78",
X"82327030",
X"70720780",
X"2570872b",
X"83c8980c",
X"515656fe",
X"c53f83c0",
X"80085281",
X"f29851e5",
X"bd3f81c8",
X"0b83c7d0",
X"0c788332",
X"70307072",
X"07802570",
X"872b83c8",
X"980c5156",
X"83c7e808",
X"5256ffb2",
X"983f83c0",
X"80085281",
X"f2a051e5",
X"8d3f8298",
X"0b83c7d0",
X"0c810b83",
X"c7d45b58",
X"83c7d008",
X"83197a32",
X"70307072",
X"07802570",
X"872b83c8",
X"980c5157",
X"8e3d7055",
X"ff1b5457",
X"57579bf2",
X"3f797084",
X"055b0851",
X"ffb1ce3f",
X"745483c0",
X"80085377",
X"5281f2a8",
X"51e4bf3f",
X"a81783c7",
X"d00c8118",
X"5877852e",
X"098106ff",
X"af3883b8",
X"0b83c7d0",
X"0c788832",
X"70307072",
X"07802570",
X"872b83c8",
X"980c5156",
X"56f4b93f",
X"81f2b855",
X"83c08008",
X"802e8f38",
X"83c7e408",
X"51ffb0f9",
X"3f83c080",
X"08557452",
X"81f2c051",
X"e3ec3f83",
X"e00b83c7",
X"d00c7889",
X"32703070",
X"72078025",
X"70872b83",
X"c8980c51",
X"5681f2cc",
X"5256e3ca",
X"3f84b00b",
X"83c7d00c",
X"788a3270",
X"30707207",
X"80257087",
X"2b83c898",
X"0c515681",
X"f2e45256",
X"e3a83f80",
X"0b83c898",
X"0c858051",
X"f9ec3f86",
X"8da051f5",
X"853f8052",
X"913d7052",
X"559f9a3f",
X"83527451",
X"9f933f63",
X"557483a6",
X"38611959",
X"78802585",
X"38745990",
X"398a7925",
X"85388a59",
X"8739788a",
X"26838538",
X"78822b55",
X"81ec9c15",
X"0804f2a6",
X"3f83c080",
X"08615755",
X"75812e09",
X"81068938",
X"83c08008",
X"10559039",
X"75ff2e09",
X"81068838",
X"83c08008",
X"812c5590",
X"75258538",
X"90558839",
X"74802483",
X"38815574",
X"51f2803f",
X"82ba399a",
X"c93f83c0",
X"80086105",
X"55748025",
X"85388055",
X"88398775",
X"25833887",
X"5574518e",
X"983f8298",
X"39f1f03f",
X"83c08008",
X"61055574",
X"80258538",
X"80558839",
X"86752583",
X"38865574",
X"51f1e93f",
X"81f63960",
X"87386280",
X"2e81ed38",
X"83c39c08",
X"83c3980c",
X"adec0b83",
X"c3a00c83",
X"c7e80851",
X"d2b43ff9",
X"e13f81d0",
X"39605680",
X"76259838",
X"ad8b0b83",
X"c3a00c83",
X"c7c41570",
X"085255d2",
X"953f7408",
X"52923975",
X"80259238",
X"83c7c415",
X"0851ffae",
X"923f8052",
X"fc1951b8",
X"3962802e",
X"81963883",
X"c7c41570",
X"0883c7d4",
X"08720c83",
X"c7d40cfc",
X"1a705351",
X"558ce53f",
X"83c08008",
X"5680518c",
X"db3f83c0",
X"80085274",
X"5188f43f",
X"75528051",
X"88ed3f80",
X"df396055",
X"807525b6",
X"3883c3a8",
X"0883c398",
X"0cadec0b",
X"83c3a00c",
X"83c7e408",
X"51d19f3f",
X"83c7e408",
X"51cec03f",
X"83c08008",
X"81ff0670",
X"5255f0c9",
X"3f74802e",
X"a7388155",
X"ab397480",
X"259e3883",
X"c7e40851",
X"ffad843f",
X"8051f0ad",
X"3f8e3962",
X"802e8938",
X"f5943f84",
X"39628738",
X"7a802ef8",
X"ff388055",
X"7483c080",
X"0c953d0d",
X"04fe3d0d",
X"83c88451",
X"8183d73f",
X"83c7f451",
X"8183cf3f",
X"f0bf3f83",
X"c0800880",
X"2e863880",
X"51818a39",
X"f0c43f83",
X"c0800880",
X"fe38f0e4",
X"3f83c080",
X"08802eb9",
X"388151ee",
X"a13f8051",
X"effa3fea",
X"993f800b",
X"83c7d00c",
X"f8973f83",
X"c0800853",
X"ff0b83c7",
X"d00cec8c",
X"3f7280cb",
X"3883c7cc",
X"3351efd4",
X"3f7251ed",
X"f13f80c0",
X"39f08c3f",
X"83c08008",
X"802eb538",
X"8151edde",
X"3f8051ef",
X"b73fe9d6",
X"3fad8b0b",
X"83c3a00c",
X"83c7d408",
X"51cfb73f",
X"ff0b83c7",
X"d00cebc8",
X"3f83c7d4",
X"08528051",
X"86d13f81",
X"51f0fe3f",
X"843d0d04",
X"fb3d0d80",
X"5283c884",
X"5180f2de",
X"3f815283",
X"c7f45180",
X"f2d43f80",
X"0b83c7cc",
X"34908080",
X"52868480",
X"8051ffaf",
X"963f83c0",
X"800881a0",
X"3883c7f0",
X"08518189",
X"8a3f8a99",
X"3f81f7b8",
X"51ffb3cc",
X"3f83c080",
X"08559c80",
X"0a5480c0",
X"805381f2",
X"ec5283c0",
X"800851f2",
X"c73f83c7",
X"e8085381",
X"f2fc5274",
X"51ffae95",
X"3f83c080",
X"088438f5",
X"d53f83c7",
X"ec085381",
X"f3885274",
X"51ffadfd",
X"3f83c080",
X"08b63887",
X"3dfc0554",
X"84808053",
X"86a88080",
X"5283c7ec",
X"0851ffac",
X"883f83c0",
X"80089338",
X"75848080",
X"2e098106",
X"8938810b",
X"83c7cc34",
X"8739800b",
X"83c7cc34",
X"83c7cc33",
X"51edc13f",
X"8151efad",
X"3f93de3f",
X"8151efa5",
X"3f8151fc",
X"f43ffa39",
X"83c08c08",
X"0283c08c",
X"0cfb3d0d",
X"0281f394",
X"0b83c39c",
X"0c81f398",
X"0b83c394",
X"0c81f39c",
X"0b83c3a8",
X"0c81f3a0",
X"0b83c3a4",
X"0c83c08c",
X"08fc050c",
X"800b83c7",
X"d40b83c0",
X"8c08f805",
X"0c83c08c",
X"08f4050c",
X"ffac903f",
X"83c08008",
X"8605fc06",
X"83c08c08",
X"f0050c02",
X"83c08c08",
X"f0050831",
X"0d833d70",
X"83c08c08",
X"f8050870",
X"840583c0",
X"8c08f805",
X"0c0c51ff",
X"a8d13f83",
X"c08c08f4",
X"05088105",
X"83c08c08",
X"f4050c83",
X"c08c08f4",
X"0508882e",
X"098106ff",
X"ab388694",
X"808051e5",
X"ea3fff0b",
X"83c7d00c",
X"800b83c8",
X"980c84d8",
X"c00b83c8",
X"940c8151",
X"ea903f81",
X"51eab53f",
X"8051eab0",
X"3f8151ea",
X"d63f8251",
X"eafe3f80",
X"51eba63f",
X"8051ebd0",
X"3f80d1ae",
X"528051da",
X"ce3ffcbc",
X"3f83c08c",
X"08fc0508",
X"0d800b83",
X"c0800c87",
X"3d0d83c0",
X"8c0c0480",
X"3d0d81ff",
X"51800b83",
X"c8a81234",
X"ff115170",
X"f438823d",
X"0d04ff3d",
X"0d737033",
X"53518111",
X"33713471",
X"81123483",
X"3d0d04ff",
X"3d0d83ca",
X"c408a82e",
X"0981068b",
X"3883cadc",
X"0883cac4",
X"0c8739a8",
X"0b83cac4",
X"0c83cac4",
X"08860570",
X"81ff0652",
X"52d0d63f",
X"833d0d04",
X"fb3d0d77",
X"79565680",
X"70715555",
X"52717525",
X"ac387216",
X"70337014",
X"7081ff06",
X"55515151",
X"71742789",
X"38811270",
X"81ff0653",
X"51718114",
X"7083ffff",
X"06555254",
X"747324d6",
X"387183c0",
X"800c873d",
X"0d04fb3d",
X"0d775689",
X"39f9c63f",
X"8351eafe",
X"3fd1dd3f",
X"83c08008",
X"802eee38",
X"83cac408",
X"86057081",
X"ff065253",
X"cfe33f81",
X"0b9088d4",
X"34f99e3f",
X"8351ead6",
X"3f9088d4",
X"337081ff",
X"06555373",
X"802eea38",
X"73862a70",
X"81065153",
X"72ffbe38",
X"73982b53",
X"80732480",
X"de38d0cd",
X"3f83c080",
X"085583c0",
X"800880cf",
X"38741675",
X"822b5454",
X"9088c013",
X"33743481",
X"15557485",
X"2e098106",
X"e8387533",
X"83c8a834",
X"81163383",
X"c8a93482",
X"163383c8",
X"aa348316",
X"3383c8ab",
X"34845283",
X"c8a851fe",
X"933f83c0",
X"800881ff",
X"06841733",
X"55537274",
X"2e8738fd",
X"ce3ffed1",
X"3980e451",
X"e9c83f87",
X"3d0d04f4",
X"3d0d7e60",
X"5955805d",
X"8075822b",
X"7183cac8",
X"120c83ca",
X"e0175b5b",
X"57767934",
X"77772e83",
X"b7387652",
X"7751ffa6",
X"ec3f8e3d",
X"fc055490",
X"5383cab0",
X"527751ff",
X"a6a73f7c",
X"5675902e",
X"09810683",
X"933883ca",
X"b051fcde",
X"3f83cab2",
X"51fcd73f",
X"83cab451",
X"fcd03f76",
X"83cac00c",
X"7751ffa3",
X"ec3f81f0",
X"bc5283c0",
X"800851c6",
X"8c3f83c0",
X"8008812e",
X"09810680",
X"d4387683",
X"cad80c82",
X"0b83cab0",
X"34ff960b",
X"83cab134",
X"7751ffa6",
X"b93f83c0",
X"80085583",
X"c0800877",
X"25883883",
X"c080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583cab2",
X"347483ca",
X"b3347683",
X"cab434ff",
X"800b83ca",
X"b5348190",
X"3983cab0",
X"3383cab1",
X"3371882b",
X"07565b74",
X"83ffff2e",
X"09810680",
X"e838fe80",
X"0b83cad8",
X"0c810b83",
X"cac00cff",
X"0b83cab0",
X"34ff0b83",
X"cab13477",
X"51ffa5c6",
X"3f83c080",
X"0883cae4",
X"0c83c080",
X"085583c0",
X"80088025",
X"883883c0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83cab234",
X"7483cab3",
X"347683ca",
X"b434ff80",
X"0b83cab5",
X"34810b83",
X"cabf34a5",
X"39748596",
X"2e098106",
X"80fe3875",
X"83cad80c",
X"7751ffa4",
X"fa3f83ca",
X"bf3383c0",
X"80080755",
X"7483cabf",
X"3483cabf",
X"33810655",
X"74802e83",
X"38845783",
X"cab43383",
X"cab53371",
X"882b0756",
X"5c748180",
X"2e098106",
X"a13883ca",
X"b23383ca",
X"b3337188",
X"2b07565b",
X"ad807527",
X"87387682",
X"07579c39",
X"76810757",
X"96397482",
X"802e0981",
X"06873876",
X"83075787",
X"397481ff",
X"268a3877",
X"83cac81b",
X"0c767934",
X"8e3d0d04",
X"803d0d72",
X"842983ca",
X"c8057008",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"727083c8",
X"a00c7084",
X"2981f6ec",
X"05700883",
X"cadc0c51",
X"51823d0d",
X"04fe3d0d",
X"8151de3f",
X"800b83ca",
X"ac0c800b",
X"83caa80c",
X"ff0b83c8",
X"a40ca80b",
X"83cac40c",
X"ae51ca91",
X"3f800b83",
X"cac85452",
X"80737084",
X"05550c81",
X"12527184",
X"2e098106",
X"ef38843d",
X"0d04fe3d",
X"0d740284",
X"05960522",
X"53537180",
X"2e963872",
X"70810554",
X"3351ca9c",
X"3fff1270",
X"83ffff06",
X"5152e739",
X"843d0d04",
X"fe3d0d02",
X"92052253",
X"82ac51e4",
X"bd3f80c3",
X"51c9f93f",
X"819651e4",
X"b13f7252",
X"83c8a851",
X"ffb43f72",
X"5283c8a8",
X"51f8cd3f",
X"83c08008",
X"81ff0651",
X"c9d63f84",
X"3d0d04ff",
X"b23d0d80",
X"d03df805",
X"51f8f73f",
X"83caac08",
X"810583ca",
X"ac0c80ce",
X"3d33cf11",
X"7081ff06",
X"51565674",
X"832688fa",
X"38758f06",
X"ff055675",
X"83c8a408",
X"2e9b3875",
X"83269638",
X"7583c8a4",
X"0c758429",
X"83cac805",
X"70085355",
X"7551f9fb",
X"3f807624",
X"88d63875",
X"842983ca",
X"c8055574",
X"08802e88",
X"c73883c8",
X"a4088429",
X"83cac805",
X"70080288",
X"0582b505",
X"33525a55",
X"7480d22e",
X"84b03874",
X"80d22490",
X"3874bf2e",
X"9c387480",
X"d02e81d5",
X"38888539",
X"7480d32e",
X"80d33874",
X"80d72e81",
X"c43887f4",
X"390282b7",
X"05330284",
X"0582b605",
X"33718280",
X"29055656",
X"c8d23f80",
X"c151c88c",
X"3ff6983f",
X"83cadf33",
X"83c8a834",
X"815283c8",
X"a851c9a9",
X"3f8151fd",
X"e73f748b",
X"3883cadc",
X"0883cac4",
X"0c8739a8",
X"0b83cac4",
X"0cc89d3f",
X"80c151c7",
X"d73ff5e3",
X"3f900b83",
X"cabf3381",
X"06565674",
X"802e8338",
X"985683ca",
X"b43383ca",
X"b5337188",
X"2b075659",
X"7481802e",
X"0981069c",
X"3883cab2",
X"3383cab3",
X"3371882b",
X"075657ad",
X"8075278c",
X"38758180",
X"07568539",
X"75a00756",
X"7583c8a8",
X"34ff0b83",
X"c8a934e0",
X"0b83c8aa",
X"34800b83",
X"c8ab3484",
X"5283c8a8",
X"51c89e3f",
X"845186ae",
X"390282b7",
X"05330284",
X"0582b605",
X"33718280",
X"2905565a",
X"c7923f78",
X"51ff9fa7",
X"3f83c080",
X"08802e8a",
X"3880ce51",
X"c6be3f86",
X"843980c1",
X"51c6b53f",
X"c7a63fc5",
X"df3f83ca",
X"d8085883",
X"75259b38",
X"83cab433",
X"83cab533",
X"71882b07",
X"fc177129",
X"7a058380",
X"055a5157",
X"8d397481",
X"802918ff",
X"80055881",
X"80578056",
X"76762e92",
X"38c6913f",
X"83c08008",
X"83c8a817",
X"34811656",
X"eb39c680",
X"3f83c080",
X"0881ff06",
X"775383c8",
X"a85256f4",
X"bf3f83c0",
X"800881ff",
X"06557575",
X"2e098106",
X"81953894",
X"51dffb3f",
X"c5fa3f80",
X"c151c5b4",
X"3fc6a53f",
X"77527851",
X"ff9dba3f",
X"805d80d0",
X"3dfdf405",
X"54765383",
X"c8a85278",
X"51ff9bc0",
X"3f0282b5",
X"05335581",
X"5a7480d7",
X"2e098106",
X"80c53877",
X"527851ff",
X"9d8b3f80",
X"d03dfdf0",
X"05547653",
X"8e3d7053",
X"795258ff",
X"9cc33f80",
X"5676762e",
X"a2387518",
X"83c8a817",
X"33713370",
X"72327030",
X"70802570",
X"30600681",
X"1d5d4051",
X"5151525a",
X"55db3982",
X"ac51def6",
X"3f79802e",
X"863880c3",
X"51843980",
X"ce51c4a8",
X"3fc5993f",
X"c3d23f83",
X"eb390282",
X"b7053302",
X"840582b6",
X"05337182",
X"80290558",
X"5a80705c",
X"5680e451",
X"dec03fc4",
X"bf3f7676",
X"2e098106",
X"8a3880ce",
X"51c3f13f",
X"83ba3980",
X"c151c3e8",
X"3f83cac0",
X"08802e82",
X"d83883ca",
X"e40880fc",
X"055580fd",
X"52745185",
X"c43f83c0",
X"80085a76",
X"8224b238",
X"ff177087",
X"2b83ffff",
X"800681f5",
X"b80583c8",
X"a8595755",
X"81805575",
X"70810557",
X"33777081",
X"055934ff",
X"157081ff",
X"06515574",
X"ea388287",
X"397682e8",
X"2e81a538",
X"7682e92e",
X"09810681",
X"ac387576",
X"5a587787",
X"32703070",
X"72078025",
X"7a8a3270",
X"30707207",
X"80257307",
X"53545a51",
X"57557580",
X"2e973878",
X"78269238",
X"a00b83c8",
X"a81a3481",
X"197081ff",
X"065a55eb",
X"39811870",
X"81ff0659",
X"558a7827",
X"ffbc388f",
X"5883c8a3",
X"183383c8",
X"a81934ff",
X"187081ff",
X"06595577",
X"8426ea38",
X"9058800b",
X"83c8a819",
X"34811870",
X"81ff0670",
X"982b5259",
X"55748025",
X"e93880c6",
X"5579858f",
X"24843880",
X"c2557483",
X"c8a83480",
X"f10b83c8",
X"ab34810b",
X"83c8ac34",
X"7983c8a9",
X"3479882c",
X"557483c8",
X"aa3480cb",
X"3982f077",
X"2580c438",
X"7680fd29",
X"fd97d305",
X"527851ff",
X"99d33f80",
X"d03dfdec",
X"055480fd",
X"5383c8a8",
X"527851ff",
X"998b3f7a",
X"81185858",
X"7780fc24",
X"83387557",
X"76882c55",
X"7483c9a5",
X"347683c9",
X"a6347783",
X"c9a73481",
X"805680cc",
X"3983cad8",
X"08588377",
X"259b3883",
X"cab43383",
X"cab53371",
X"882b07fc",
X"1971297a",
X"05838005",
X"5a575a8d",
X"39768180",
X"2918ff80",
X"05588180",
X"56775278",
X"51ff98e1",
X"3f80d03d",
X"fdec0554",
X"755383c8",
X"a8527851",
X"ff989a3f",
X"7551f6ac",
X"3fc1a93f",
X"ffbfe13f",
X"8b3983ca",
X"a8088105",
X"83caa80c",
X"80d03d0d",
X"04f6cc3f",
X"fc39fc3d",
X"0d767871",
X"842983ca",
X"c8057008",
X"51535353",
X"709e3880",
X"ce723480",
X"cf0b8113",
X"3480ce0b",
X"82133480",
X"c50b8313",
X"34708413",
X"3480e739",
X"83cae013",
X"335480d2",
X"72347382",
X"2a708106",
X"515180cf",
X"53708438",
X"80d75372",
X"811334a0",
X"0b821334",
X"73830651",
X"70812e9e",
X"38708124",
X"88387080",
X"2e8f389f",
X"3970822e",
X"92387083",
X"2e923893",
X"3980d855",
X"8e3980d3",
X"55893980",
X"cd558439",
X"80c45574",
X"83133480",
X"c40b8413",
X"34800b85",
X"1334863d",
X"0d0483c8",
X"a00883c0",
X"800c0480",
X"3d0d83c8",
X"a0088429",
X"81f78c05",
X"700883c0",
X"800c5182",
X"3d0d04fc",
X"3d0d7678",
X"53548153",
X"80558739",
X"71107310",
X"54527372",
X"26517280",
X"2ea73870",
X"802e8638",
X"718025e8",
X"3872802e",
X"98387174",
X"26893873",
X"72317574",
X"07565472",
X"812a7281",
X"2a5353e5",
X"39735178",
X"83387451",
X"7083c080",
X"0c863d0d",
X"04fe3d0d",
X"80537552",
X"7451ffa3",
X"3f843d0d",
X"04fe3d0d",
X"81537552",
X"7451ff93",
X"3f843d0d",
X"04fb3d0d",
X"77795555",
X"80567476",
X"25863874",
X"30558156",
X"73802588",
X"38733076",
X"81325754",
X"80537352",
X"7451fee7",
X"3f83c080",
X"08547580",
X"2e873883",
X"c0800830",
X"547383c0",
X"800c873d",
X"0d04fa3d",
X"0d787a57",
X"55805774",
X"77258638",
X"74305581",
X"57759f2c",
X"54815375",
X"74327431",
X"527451fe",
X"aa3f83c0",
X"80085476",
X"802e8738",
X"83c08008",
X"30547383",
X"c0800c88",
X"3d0d04fc",
X"3d0d7655",
X"80750c80",
X"0b84160c",
X"800b8816",
X"0c800b8c",
X"160c83c8",
X"845180e9",
X"b13f83c7",
X"f45180e9",
X"a93f87a6",
X"80337081",
X"ff067071",
X"842a0651",
X"5152d6dd",
X"3f71812a",
X"81327281",
X"32718106",
X"71810631",
X"84180c54",
X"5471832a",
X"81327282",
X"2a813270",
X"81067271",
X"31780c51",
X"535387a0",
X"903387a0",
X"91337081",
X"ff067073",
X"06813281",
X"0688190c",
X"51535383",
X"c0800880",
X"2e80c238",
X"83c08008",
X"812a7081",
X"0683c080",
X"08810631",
X"84170c52",
X"83c08008",
X"832a83c0",
X"8008822a",
X"71810671",
X"81063177",
X"0c535383",
X"c0800884",
X"2a810688",
X"160c83c0",
X"8008852a",
X"81068c16",
X"0c863d0d",
X"04fe3d0d",
X"74765452",
X"7151feab",
X"3f72812e",
X"a2388173",
X"268d3872",
X"822ea838",
X"72832e9c",
X"38e63971",
X"08e23884",
X"1208dd38",
X"881208d8",
X"38a53988",
X"1208812e",
X"9e389139",
X"88120881",
X"2e953871",
X"08913884",
X"12088c38",
X"8c120881",
X"2e098106",
X"ffb23884",
X"3d0d04fb",
X"3d0d7802",
X"84059f05",
X"33555680",
X"0b81eeb4",
X"56538173",
X"2b740652",
X"71802e83",
X"38815274",
X"70820556",
X"22707390",
X"2b079080",
X"9c0c5181",
X"13537288",
X"2e098106",
X"d9388053",
X"83caec13",
X"33517081",
X"ff2eb238",
X"701081ec",
X"d4057022",
X"55518073",
X"17703370",
X"1081ecd4",
X"05702251",
X"51515252",
X"73712e91",
X"38811252",
X"71862e09",
X"8106f138",
X"7390809c",
X"0c811353",
X"72862e09",
X"8106ffb8",
X"38805372",
X"16703351",
X"517081ff",
X"2e943870",
X"1081ecd4",
X"05702270",
X"84808007",
X"90809c0c",
X"51518113",
X"5372862e",
X"098106d7",
X"38805372",
X"16517033",
X"83caec14",
X"34811353",
X"72862e09",
X"8106ec38",
X"873d0d04",
X"04fe3d0d",
X"75028405",
X"93053381",
X"06525270",
X"88387190",
X"80940c8e",
X"3970812e",
X"09810686",
X"38719080",
X"980c843d",
X"0d04fb3d",
X"0d78982b",
X"70982c7b",
X"982b7098",
X"2c029005",
X"9f053381",
X"0683cb88",
X"11703370",
X"982b7098",
X"2c51585c",
X"5a565155",
X"51547074",
X"2e098106",
X"943883ca",
X"e8123370",
X"982b7098",
X"2c515256",
X"70732eb1",
X"38737534",
X"7283cae8",
X"133483ca",
X"e93383cb",
X"89337198",
X"2b71902b",
X"0783cae8",
X"3370882b",
X"720783cb",
X"88337107",
X"9080b80c",
X"52595354",
X"52873d0d",
X"04fe3d0d",
X"74811133",
X"71337188",
X"2b0783c0",
X"800c5351",
X"843d0d04",
X"83caf433",
X"83c0800c",
X"04f53d0d",
X"02bb0533",
X"028405bf",
X"05330288",
X"0580c305",
X"33028c05",
X"80c60522",
X"665c5a5e",
X"5c567a55",
X"7b548953",
X"a1527d51",
X"80df843f",
X"83c08008",
X"81ff0683",
X"c0800c8d",
X"3d0d0483",
X"c08c0802",
X"83c08c0c",
X"f53d0d83",
X"c08c0888",
X"050883c0",
X"8c088f05",
X"3383c08c",
X"08920522",
X"028c0573",
X"900583c0",
X"8c08e805",
X"0c83c08c",
X"08f8050c",
X"83c08c08",
X"f0050c83",
X"c08c08ec",
X"050c83c0",
X"8c08f405",
X"0c800b83",
X"c08c08f0",
X"050883c0",
X"8c08e005",
X"0c83c08c",
X"08fc050c",
X"83c08c08",
X"f0050889",
X"278a3889",
X"0b83c08c",
X"08e0050c",
X"83c08c08",
X"e0050886",
X"0587fffc",
X"0683c08c",
X"08e0050c",
X"0283c08c",
X"08e00508",
X"310d853d",
X"705583c0",
X"8c08ec05",
X"085483c0",
X"8c08f005",
X"085383c0",
X"8c08f405",
X"085283c0",
X"8c08e405",
X"0c80e8dd",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"e4050883",
X"c08c08ec",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"802e8c38",
X"83c08c08",
X"f805080d",
X"89c83983",
X"c08c08f0",
X"0508802e",
X"89a63883",
X"c08c08ec",
X"05088105",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e0050884",
X"2ea93884",
X"0b83c08c",
X"08e00508",
X"2588c738",
X"83c08c08",
X"e0050885",
X"2e859b38",
X"83c08c08",
X"e00508a1",
X"2e87ad38",
X"88ac3980",
X"0b83c08c",
X"08ec0508",
X"85053383",
X"c08c08e0",
X"050c83c0",
X"8c08fc05",
X"0c83c08c",
X"08e00508",
X"832e0981",
X"06888338",
X"83c08c08",
X"e8050881",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"812687e6",
X"38810b83",
X"c08c08e0",
X"050880d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"fc050c83",
X"c08c08ec",
X"05088205",
X"3383c08c",
X"08e00508",
X"87053483",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c80",
X"0b83c08c",
X"08e00508",
X"8b053483",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"f4050c80",
X"0b83c08c",
X"08e00508",
X"8c053483",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c80",
X"0b83c08c",
X"08e00508",
X"8d053483",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"f4050c80",
X"0b83c08c",
X"08e00508",
X"8e052383",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c80",
X"0b83c08c",
X"08e00508",
X"8a053483",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"05709405",
X"08fcffff",
X"06719405",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"ec050886",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"83c08c08",
X"e0050883",
X"c08c08fc",
X"05082e09",
X"8106b638",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"83c08c08",
X"fc050883",
X"c08c08e0",
X"05088b05",
X"3483c08c",
X"08ec0508",
X"87053383",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08812e8f",
X"3883c08c",
X"08e00508",
X"822eb738",
X"848c3983",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"f4050c82",
X"0b83c08c",
X"08e00508",
X"8a053483",
X"d93983c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c83c0",
X"8c08fc05",
X"0883c08c",
X"08e00508",
X"8a053483",
X"a13983c0",
X"8c08fc05",
X"08802e83",
X"953883c0",
X"8c08ec05",
X"08830533",
X"830683c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"832e0981",
X"0682f338",
X"83c08c08",
X"ec050882",
X"05337098",
X"2b83c08c",
X"08e0050c",
X"83c08c08",
X"e4050c83",
X"c08c08e0",
X"05088025",
X"82cc3883",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"f4050c83",
X"c08c08ec",
X"05088605",
X"3383c08c",
X"08e00508",
X"80d60534",
X"83c08c08",
X"e0050884",
X"0583c08c",
X"08ec0508",
X"8205338f",
X"0683c08c",
X"08e4050c",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050883c0",
X"8c08e005",
X"083483c0",
X"8c08ec05",
X"08840533",
X"83c08c08",
X"e0050881",
X"0534800b",
X"83c08c08",
X"e0050882",
X"053483c0",
X"8c08e005",
X"0808ff83",
X"ff068280",
X"0783c08c",
X"08e00508",
X"0c83c08c",
X"08e80508",
X"81053381",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e0050883",
X"c08c08e8",
X"05088105",
X"34818339",
X"83c08c08",
X"fc050880",
X"2e80f738",
X"83c08c08",
X"ec050886",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"a22e0981",
X"0680d738",
X"83c08c08",
X"ec050888",
X"053383c0",
X"8c08ec05",
X"08870533",
X"71828029",
X"0583c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c5283",
X"c08c08e4",
X"050c83c0",
X"8c08f405",
X"0c83c08c",
X"08e40508",
X"83c08c08",
X"e0050888",
X"052383c0",
X"8c08ec05",
X"083383c0",
X"8c08f005",
X"08713170",
X"83ffff06",
X"83c08c08",
X"f0050c83",
X"c08c08e0",
X"050c83c0",
X"8c08ec05",
X"080583c0",
X"8c08ec05",
X"0cf6d039",
X"83c08c08",
X"f805080d",
X"83c08c08",
X"f0050883",
X"c08c08e0",
X"050c83c0",
X"8c08f805",
X"080d83c0",
X"8c08e005",
X"0883c080",
X"0c8d3d0d",
X"83c08c0c",
X"0483c08c",
X"080283c0",
X"8c0ce73d",
X"0d83c08c",
X"08880508",
X"02840583",
X"c08c08e8",
X"050c83c0",
X"8c08d405",
X"0c800b83",
X"cb903483",
X"c08c08d4",
X"05089005",
X"83c08c08",
X"c4050c80",
X"0b83c08c",
X"08c40508",
X"34800b83",
X"c08c08c4",
X"05088105",
X"34800b83",
X"c08c08c8",
X"050c83c0",
X"8c08c805",
X"0880d829",
X"83c08c08",
X"c4050805",
X"83c08c08",
X"ffb8050c",
X"800b83c0",
X"8c08ffb8",
X"050880d8",
X"050c83c0",
X"8c08ffb8",
X"05088405",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"c8050883",
X"c08c08ff",
X"b8050834",
X"880b83c0",
X"8c08ffb8",
X"05088105",
X"34800b83",
X"c08c08ff",
X"b8050882",
X"053483c0",
X"8c08ffb8",
X"050808ff",
X"a1ff06a0",
X"800783c0",
X"8c08ffb8",
X"05080c83",
X"c08c08c8",
X"05088105",
X"7081ff06",
X"83c08c08",
X"c8050c83",
X"c08c08ff",
X"b8050c81",
X"0b83c08c",
X"08c80508",
X"27fedb38",
X"83c08c08",
X"ec057054",
X"83c08c08",
X"cc050c92",
X"5283c08c",
X"08d40508",
X"5180dc84",
X"3f83c080",
X"0881ff06",
X"7083c08c",
X"08ffb805",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffbc05",
X"0891c638",
X"83c08c08",
X"f40551f1",
X"8c3f83c0",
X"800883ff",
X"ff0683c0",
X"8c08f605",
X"5283c08c",
X"08e0050c",
X"f0f33f83",
X"c0800883",
X"ffff0683",
X"c08c08fd",
X"053383c0",
X"8c08ffbc",
X"050883c0",
X"8c08c805",
X"0c83c08c",
X"08c0050c",
X"83c08c08",
X"dc050c83",
X"c08c08c8",
X"050883c0",
X"8c08c005",
X"082780fe",
X"3883c08c",
X"08cc0508",
X"5483c08c",
X"08c80508",
X"53895283",
X"c08c08d4",
X"05085180",
X"db8b3f83",
X"c0800881",
X"ff0683c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffbc",
X"050883eb",
X"3883c08c",
X"08ee0551",
X"eff33f83",
X"c0800883",
X"ffff0653",
X"83c08c08",
X"c8050852",
X"83c08c08",
X"d4050851",
X"f0b53f83",
X"c08c08c8",
X"05088105",
X"7081ff06",
X"83c08c08",
X"c8050c83",
X"c08c08ff",
X"b8050cfe",
X"f23983c0",
X"8c08c405",
X"08810533",
X"83c08c08",
X"c0050c83",
X"c08c08c0",
X"0508839e",
X"3883c08c",
X"08c00508",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"e0050888",
X"de2e0981",
X"068b3881",
X"0b83c08c",
X"08ffb805",
X"0c83c08c",
X"08dc0508",
X"858e2e09",
X"810682c5",
X"38817083",
X"c08c08ff",
X"b8050806",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"c8050c83",
X"c08c08ff",
X"b8050880",
X"2e829e38",
X"83c08c08",
X"c8050883",
X"c08c08c4",
X"05088105",
X"3483c08c",
X"08c00508",
X"83c08c08",
X"c4050887",
X"053483c0",
X"8c08c005",
X"0883c08c",
X"08c40508",
X"8b053483",
X"c08c08c0",
X"050883c0",
X"8c08c405",
X"088c0534",
X"830b83c0",
X"8c08c405",
X"088d0534",
X"83c08c08",
X"c0050883",
X"c08c08c4",
X"05088e05",
X"23830b83",
X"c08c08c4",
X"05088a05",
X"3483c08c",
X"08c40508",
X"94050883",
X"80800783",
X"c08c08c4",
X"05089405",
X"0c83caf4",
X"337083c0",
X"8c08c805",
X"080583c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb8",
X"050883ca",
X"f43483c0",
X"8c08ffbc",
X"050883c0",
X"8c08c405",
X"08940534",
X"83c08c08",
X"c8050883",
X"c08c08c4",
X"050880d6",
X"053483c0",
X"8c08c805",
X"0883c08c",
X"08c40508",
X"8405348e",
X"0b83c08c",
X"08c40508",
X"85053483",
X"c08c08c0",
X"050883c0",
X"8c08c405",
X"08860534",
X"83c08c08",
X"c4050884",
X"0508ff83",
X"ff068280",
X"0783c08c",
X"08c40508",
X"84050ca2",
X"3981db0b",
X"83c08c08",
X"ffb8050c",
X"8cc33983",
X"c08c08ff",
X"bc050883",
X"c08c08ff",
X"b8050c8c",
X"b03983c0",
X"8c08f105",
X"335283c0",
X"8c08d405",
X"085180d7",
X"903f800b",
X"83c08c08",
X"c4050881",
X"053383c0",
X"8c08ffb8",
X"050c83c0",
X"8c08c805",
X"0c83c08c",
X"08c80508",
X"83c08c08",
X"ffb80508",
X"278acb38",
X"83c08c08",
X"c8050880",
X"d8297083",
X"c08c08c4",
X"05080570",
X"88057083",
X"053383c0",
X"8c08ffb8",
X"050c83c0",
X"8c08cc05",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08d8050c",
X"83c08c08",
X"ffb80508",
X"88893883",
X"c08c08ff",
X"bc05088d",
X"053383c0",
X"8c08d005",
X"0c83c08c",
X"08d00508",
X"87ed3883",
X"c08c08cc",
X"05082202",
X"84057186",
X"0587fffc",
X"0683c08c",
X"08ffb805",
X"0c83c08c",
X"08e4050c",
X"83c08c08",
X"c0050c02",
X"83c08c08",
X"ffb80508",
X"310d893d",
X"705983c0",
X"8c08c005",
X"085883c0",
X"8c08ffbc",
X"05088705",
X"335783c0",
X"8c08ffb8",
X"050ca255",
X"83c08c08",
X"d0050854",
X"86538181",
X"5283c08c",
X"08d40508",
X"5180c9c3",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"d0050c83",
X"c08c08d0",
X"050881c0",
X"3883c08c",
X"08ffbc05",
X"08960553",
X"83c08c08",
X"c0050852",
X"83c08c08",
X"ffb80508",
X"51acf73f",
X"83c08008",
X"81ff0683",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b8050880",
X"2e818538",
X"83c08c08",
X"ffbc0508",
X"940583c0",
X"8c08ffbc",
X"05089605",
X"3370862a",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"c0050c83",
X"c08c08ff",
X"b8050883",
X"2e098106",
X"80c63883",
X"c08c08ff",
X"b8050883",
X"c08c08cc",
X"05088205",
X"3483caf4",
X"33708105",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb80508",
X"83caf434",
X"83c08c08",
X"ffbc0508",
X"83c08c08",
X"c0050834",
X"83c08c08",
X"e405080d",
X"83c08c08",
X"d0050881",
X"ff0683c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffbc",
X"0508fbe3",
X"3883c08c",
X"08d80508",
X"83c08c08",
X"c4050805",
X"88057082",
X"05335183",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b8050883",
X"2e098106",
X"80e33883",
X"c08c08ff",
X"bc050883",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b8050881",
X"057081ff",
X"065183c0",
X"8c08ffb8",
X"050c810b",
X"83c08c08",
X"ffb80508",
X"27dd3880",
X"0b83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"08810570",
X"81ff0651",
X"83c08c08",
X"ffb8050c",
X"970b83c0",
X"8c08ffb8",
X"050827dd",
X"3883c08c",
X"08e00508",
X"80f93270",
X"30708025",
X"515183c0",
X"8c08ffb8",
X"050c83c0",
X"8c08dc05",
X"08912e09",
X"810680f9",
X"3883c08c",
X"08ffb805",
X"08802e80",
X"ec3883c0",
X"8c08c805",
X"0880e238",
X"850b83c0",
X"8c08c405",
X"08a60534",
X"a00b83c0",
X"8c08c405",
X"08a70534",
X"850b83c0",
X"8c08c405",
X"08a80534",
X"80c00b83",
X"c08c08c4",
X"0508a905",
X"34860b83",
X"c08c08c4",
X"0508aa05",
X"34900b83",
X"c08c08c4",
X"0508ab05",
X"34860b83",
X"c08c08c4",
X"0508ac05",
X"34a00b83",
X"c08c08c4",
X"0508ad05",
X"3483c08c",
X"08e00508",
X"89d83270",
X"30708025",
X"515183c0",
X"8c08ffb8",
X"050c83c0",
X"8c08dc05",
X"0883edec",
X"2e098106",
X"80f63881",
X"7083c08c",
X"08ffb805",
X"080683c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb8",
X"0508802e",
X"80ce3883",
X"c08c08c8",
X"050880c4",
X"38840b83",
X"c08c08c4",
X"0508aa05",
X"3480c00b",
X"83c08c08",
X"c40508ab",
X"0534840b",
X"83c08c08",
X"c40508ac",
X"0534900b",
X"83c08c08",
X"c40508ad",
X"053483c0",
X"8c08ffbc",
X"050883c0",
X"8c08c405",
X"088c0534",
X"83c08c08",
X"e0050880",
X"f9327030",
X"70802551",
X"5183c08c",
X"08ffb805",
X"0c83c08c",
X"08dc0508",
X"862e0981",
X"0680c338",
X"817083c0",
X"8c08ffb8",
X"05080683",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"b8050880",
X"2e9c3883",
X"c08c08c8",
X"05089338",
X"83c08c08",
X"ffbc0508",
X"83c08c08",
X"c405088d",
X"053483c0",
X"8c08e005",
X"08b4b432",
X"70307080",
X"25515183",
X"c08c08ff",
X"b8050c83",
X"c08c08dc",
X"05089089",
X"2e098106",
X"a23883c0",
X"8c08ffb8",
X"0508802e",
X"963883c0",
X"8c08c805",
X"088d3882",
X"0b83c08c",
X"08c40508",
X"8d053483",
X"c08c08c8",
X"050880d8",
X"2983c08c",
X"08c40508",
X"05708405",
X"70830533",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"cc050c83",
X"c08c08c0",
X"050c8058",
X"805783c0",
X"8c08ffb8",
X"05085680",
X"5580548a",
X"53a15283",
X"c08c08d4",
X"05085180",
X"c1f53f83",
X"c0800881",
X"ff067030",
X"709f2a51",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffbc0508",
X"a02e8c38",
X"83c08c08",
X"ffb80508",
X"f5dd3883",
X"c08c08c0",
X"05088b05",
X"3383c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"08802eb4",
X"3883c08c",
X"08cc0508",
X"83053383",
X"c08c08ff",
X"b8050c80",
X"58805783",
X"c08c08ff",
X"b8050856",
X"80558054",
X"8b53a152",
X"83c08c08",
X"d4050851",
X"80c0f03f",
X"83c08c08",
X"c8050881",
X"057081ff",
X"0683c08c",
X"08c40508",
X"81053352",
X"83c08c08",
X"c8050c83",
X"c08c08ff",
X"b8050cf5",
X"a439800b",
X"83c08c08",
X"c8050c83",
X"c08c08c8",
X"050880d8",
X"2983c08c",
X"08d40508",
X"05709a05",
X"3383c08c",
X"08ffb805",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffb805",
X"08822e09",
X"8106a938",
X"83cb9056",
X"81558054",
X"83c08c08",
X"ffb80508",
X"5383c08c",
X"08ffbc05",
X"08970533",
X"5283c08c",
X"08d40508",
X"51e0ae3f",
X"83c08c08",
X"c8050881",
X"057081ff",
X"0683c08c",
X"08c8050c",
X"83c08c08",
X"ffb8050c",
X"810b83c0",
X"8c08c805",
X"0827fefb",
X"38810b83",
X"c08c08c4",
X"05083480",
X"0b83c08c",
X"08ffb805",
X"0c83c08c",
X"08e80508",
X"0d83c08c",
X"08ffb805",
X"0883c080",
X"0c9b3d0d",
X"83c08c0c",
X"04f43d0d",
X"901f5980",
X"0b811a33",
X"555b7a74",
X"2781ad38",
X"7a80d829",
X"198a1133",
X"55557383",
X"2e098106",
X"81883894",
X"15335780",
X"527651dd",
X"e03f8053",
X"80527651",
X"de803fb3",
X"e43f83c0",
X"80085c80",
X"587781c4",
X"291c8711",
X"33555573",
X"802e80c0",
X"38740881",
X"ecc82e09",
X"8106b538",
X"80755b56",
X"7580d829",
X"1a9a1133",
X"55557383",
X"2e098106",
X"9238a415",
X"70335555",
X"76742787",
X"38ff1454",
X"73753481",
X"167081ff",
X"06575481",
X"7627d138",
X"81187081",
X"ff065954",
X"8f7827ff",
X"a43883ca",
X"f433ff05",
X"547383ca",
X"f434811b",
X"7081ff06",
X"811b335f",
X"5c547c7b",
X"26fed538",
X"800b83c0",
X"800c8e3d",
X"0d0483c0",
X"8c080283",
X"c08c0ce6",
X"3d0d83c0",
X"8c088805",
X"08028405",
X"71900570",
X"337083c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08cc05",
X"0c83c08c",
X"08dc050c",
X"83c08c08",
X"e0050c83",
X"c08c08ff",
X"a4050880",
X"2e9f8c38",
X"800b83c0",
X"8c08cc05",
X"08810533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"d4050c83",
X"c08c08d4",
X"050883c0",
X"8c08ffa4",
X"0508259e",
X"d43883c0",
X"8c08d405",
X"0880d829",
X"83c08c08",
X"cc050805",
X"84057086",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"9de038b1",
X"8a3f83c0",
X"8c08ffbc",
X"050880d4",
X"050883c0",
X"8008269d",
X"c9380283",
X"c08c08ff",
X"bc050881",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08d805",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08fc0523",
X"83c08c08",
X"ffa40508",
X"860583fc",
X"0683c08c",
X"08ffa405",
X"0c0283c0",
X"8c08ffa4",
X"0508310d",
X"853d7055",
X"83c08c08",
X"fc055483",
X"c08c08ff",
X"bc050853",
X"83c08c08",
X"e0050852",
X"83c08c08",
X"c0050cb8",
X"e23f83c0",
X"800881ff",
X"0683c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"089c9238",
X"83c08c08",
X"ffbc0508",
X"87053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e80d538",
X"83c08c08",
X"ffbc0508",
X"86053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050882",
X"2e098106",
X"b33883c0",
X"8c08fc05",
X"2283c08c",
X"08ffa405",
X"0c870b83",
X"c08c08ff",
X"a4050827",
X"973883c0",
X"8c08c005",
X"08820552",
X"83c08c08",
X"c0050833",
X"51d7b43f",
X"83c08c08",
X"ffbc0508",
X"86053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050883",
X"2e098106",
X"9afb3883",
X"c08c08ff",
X"bc050892",
X"0583c08c",
X"08ffbc05",
X"08890533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"c4050c83",
X"c08c08ff",
X"a4050883",
X"2eb63883",
X"c08c08c4",
X"05088205",
X"3383c08c",
X"08fc0522",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa80508",
X"83c08c08",
X"ffac0508",
X"269a9638",
X"800b83c0",
X"8c08e405",
X"0c800b83",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a4050883",
X"2e098106",
X"88c13883",
X"c08c08c0",
X"05083383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"b005082e",
X"09810687",
X"fa3883c0",
X"8c08c005",
X"08810533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"942e0981",
X"0687d838",
X"83c08c08",
X"c0050882",
X"05337081",
X"0683c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffb005",
X"082e8a38",
X"880b83c0",
X"8c08e405",
X"0c83c08c",
X"08ffa805",
X"08812a70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e913883",
X"c08c08e4",
X"05088407",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"a8050882",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e91",
X"3883c08c",
X"08e40508",
X"820783c0",
X"8c08e405",
X"0c83c08c",
X"08ffa805",
X"08832a70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e913883",
X"c08c08e4",
X"05088107",
X"83c08c08",
X"e4050c83",
X"c08c08c0",
X"05088305",
X"3370982b",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa40508",
X"80259138",
X"83c08c08",
X"e4050890",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"ffa80508",
X"81ff0670",
X"852a7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"913883c0",
X"8c08e405",
X"08a00783",
X"c08c08e4",
X"050c83c0",
X"8c08ffa8",
X"0508842a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9238",
X"83c08c08",
X"e4050880",
X"c00783c0",
X"8c08e405",
X"0c83c08c",
X"08ffa805",
X"08862a70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e923883",
X"c08c08e4",
X"05088180",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"ffa80508",
X"810683c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"923883c0",
X"8c08e405",
X"08828007",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"a8050881",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e92",
X"3883c08c",
X"08e40508",
X"84800783",
X"c08c08e4",
X"050c83c0",
X"8c08c005",
X"08840533",
X"70982b83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a4050880",
X"25923883",
X"c08c08e4",
X"05088880",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"c0050885",
X"05337098",
X"2b83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"08802592",
X"3883c08c",
X"08e40508",
X"90800783",
X"c08c08e4",
X"050c83c0",
X"8c08c005",
X"08820533",
X"7081ff06",
X"70852a70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a4050880",
X"2e923883",
X"c08c08e4",
X"0508a080",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"ffa80508",
X"842a7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"933883c0",
X"8c08e405",
X"0880c080",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"ffa80508",
X"862a7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"933883c0",
X"8c08e405",
X"08818080",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"ffac0508",
X"982b83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"05088025",
X"933883c0",
X"8c08e405",
X"08828080",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"c0050887",
X"05337098",
X"2b83c08c",
X"08c00508",
X"89053370",
X"982b7098",
X"2c73982c",
X"81800554",
X"515383c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050883c0",
X"8c08f805",
X"2380ff0b",
X"83c08c08",
X"ffa40508",
X"3183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08fa0523",
X"84d93980",
X"0b83c08c",
X"08e4050c",
X"81800b83",
X"c08c08f8",
X"05238180",
X"0b83c08c",
X"08fa0523",
X"84b93983",
X"c08c08ff",
X"b0050810",
X"83c08c08",
X"05f80583",
X"c08c08ff",
X"b0050884",
X"2983c08c",
X"08ffb005",
X"08100583",
X"c08c08c4",
X"05080570",
X"84057033",
X"83c08c08",
X"c0050805",
X"703383c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffb8",
X"05082383",
X"c08c08ff",
X"a8050881",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508902e",
X"098106be",
X"3883c08c",
X"08ffa805",
X"083383c0",
X"8c08c005",
X"08058105",
X"70337082",
X"802983c0",
X"8c08ffb4",
X"05080551",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffb805",
X"082383c0",
X"8c08ffac",
X"05088605",
X"2283c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa805",
X"08a23883",
X"c08c08ff",
X"ac050888",
X"052283c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"050881ff",
X"2e80e538",
X"83c08c08",
X"ffb80508",
X"227083c0",
X"8c08ffa8",
X"05083170",
X"82802971",
X"3183c08c",
X"08ffac05",
X"08880522",
X"7083c08c",
X"08ffa805",
X"08317073",
X"355383c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c5183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"b8050823",
X"83c08c08",
X"ffb00508",
X"81057081",
X"ff0683c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa4",
X"050c810b",
X"83c08c08",
X"ffb00508",
X"27fce038",
X"800b83c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffb0",
X"05081083",
X"c08c08c4",
X"05080570",
X"90057033",
X"83c08c08",
X"c0050805",
X"70337281",
X"05337072",
X"06515351",
X"83c08c08",
X"ffa8050c",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e9b",
X"38900b83",
X"c08c08ff",
X"b005082b",
X"83c08c08",
X"e4050807",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"b0050881",
X"057081ff",
X"0683c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa405",
X"0c970b83",
X"c08c08ff",
X"b0050827",
X"fef43883",
X"c08c08f8",
X"052283c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508bf26",
X"913883c0",
X"8c08e405",
X"08820783",
X"c08c08e4",
X"050c81c0",
X"0b83c08c",
X"08ffa405",
X"08279138",
X"83c08c08",
X"e4050881",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"fa052283",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a40508bf",
X"26913883",
X"c08c08e4",
X"05088807",
X"83c08c08",
X"e4050c81",
X"c00b83c0",
X"8c08ffa4",
X"05082791",
X"3883c08c",
X"08e40508",
X"840783c0",
X"8c08e405",
X"0c83c08c",
X"08ffbc05",
X"08900533",
X"83c08c08",
X"e4050883",
X"c08c08ff",
X"a4050c83",
X"c08c08c4",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffbc",
X"05088c05",
X"082e85e0",
X"3883c08c",
X"08ffa405",
X"0883c08c",
X"08ffbc05",
X"088c050c",
X"83c08c08",
X"ffbc0508",
X"89053383",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a8050880",
X"2e859a38",
X"83c08c08",
X"e40583c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffa4",
X"05088f06",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"b0050c83",
X"c08c08d0",
X"050c83c0",
X"8c08ffa8",
X"0508822e",
X"09810681",
X"c238800b",
X"83c08c08",
X"ffa40508",
X"862a7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffa8",
X"05082e8c",
X"3881c00b",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffb00508",
X"872a7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"943883c0",
X"8c08ffa8",
X"05088190",
X"3283c08c",
X"08ffa805",
X"0c83c08c",
X"08ffb005",
X"08842a70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e943883",
X"c08c08ff",
X"a8050880",
X"d03283c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffb0",
X"050883c0",
X"8c08ffa8",
X"05083283",
X"c08c08ff",
X"b0050c80",
X"0b83c08c",
X"08f0050c",
X"800b83c0",
X"8c08f405",
X"23800b81",
X"eec43383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"b805082e",
X"82d33883",
X"c08c08f0",
X"0581eec4",
X"0b83c08c",
X"08ffac05",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"ffac0508",
X"3383c08c",
X"08ffac05",
X"08810533",
X"81722b81",
X"722b0770",
X"83c08c08",
X"ffb00508",
X"065283c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffa8",
X"05082e09",
X"810681be",
X"3883c08c",
X"08ffb805",
X"08852680",
X"f63883c0",
X"8c08ffac",
X"05088205",
X"337081ff",
X"0683c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"08802e80",
X"ca3883c0",
X"8c08ffb8",
X"050883c0",
X"8c08ffb8",
X"05088105",
X"7081ff06",
X"83c08c08",
X"c8050873",
X"055383c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffa4",
X"05083483",
X"c08c08ff",
X"ac050883",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"9d38810b",
X"83c08c08",
X"ffa40508",
X"2b83c08c",
X"08d00508",
X"080783c0",
X"8c08d005",
X"080c83c0",
X"8c08ffac",
X"05088405",
X"703383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa4",
X"0508fdc8",
X"3883c08c",
X"08f00552",
X"8051c1fb",
X"3f83c08c",
X"08e40508",
X"5283c08c",
X"08c40508",
X"51c3b63f",
X"83c08c08",
X"fb053370",
X"81800a29",
X"810a0570",
X"982c5583",
X"c08c08ff",
X"a4050c83",
X"c08c08f9",
X"05337081",
X"800a2981",
X"0a057098",
X"2c5583c0",
X"8c08ffa4",
X"050c83c0",
X"8c08c405",
X"085383c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa8",
X"050cc38e",
X"3f83c08c",
X"08ffbc05",
X"08880533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e84e1",
X"3883c08c",
X"08ffbc05",
X"08900533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"812684c1",
X"38807081",
X"ef840b81",
X"ef840b81",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffb4",
X"05082e81",
X"ae3883c0",
X"8c08ffac",
X"05088429",
X"83c08c08",
X"ffa80508",
X"05703383",
X"c08c08c0",
X"05080570",
X"33728105",
X"33707206",
X"51535183",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2eaa3881",
X"0b83c08c",
X"08ffac05",
X"082b83c0",
X"8c08ffb4",
X"05080770",
X"83ffff06",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffac0508",
X"81057081",
X"ff0681ef",
X"84718429",
X"71057081",
X"05335153",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"fed43883",
X"c08c08ff",
X"bc05088a",
X"052283c0",
X"8c08c005",
X"0c83c08c",
X"08ffb405",
X"0883c08c",
X"08c00508",
X"2e82ae38",
X"800b83c0",
X"8c08e805",
X"0c800b83",
X"c08c08ec",
X"05238070",
X"83c08c08",
X"e80583c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffb0",
X"050c81af",
X"3983c08c",
X"08ffb405",
X"0883c08c",
X"08ffac05",
X"082c7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"80e73883",
X"c08c08ff",
X"b0050883",
X"c08c08ff",
X"b0050881",
X"057081ff",
X"0683c08c",
X"08ffb805",
X"08730583",
X"c08c08ff",
X"bc050890",
X"053383c0",
X"8c08ffac",
X"05088429",
X"05535383",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a8050881",
X"ef860533",
X"83c08c08",
X"ffa40508",
X"3483c08c",
X"08ffac05",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a4050c8f",
X"0b83c08c",
X"08ffac05",
X"082783c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb0",
X"05088526",
X"8c3883c0",
X"8c08ffa4",
X"0508fea9",
X"3883c08c",
X"08e80552",
X"8051ffbc",
X"aa3f83c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffbc",
X"05088a05",
X"2383c08c",
X"08ffbc05",
X"0880d205",
X"3383c08c",
X"08ffbc05",
X"0880d405",
X"080583c0",
X"8c08ffbc",
X"050880d4",
X"050c83c0",
X"8c08d805",
X"080d83c0",
X"8c08d405",
X"0881800a",
X"2981800a",
X"0570982c",
X"83c08c08",
X"cc050881",
X"053383c0",
X"8c08ffa8",
X"050c5183",
X"c08c08d4",
X"050c83c0",
X"8c08ffa8",
X"050883c0",
X"8c08d405",
X"0824e1ae",
X"38800b83",
X"c08c08ff",
X"a8050c83",
X"c08c08dc",
X"05080d83",
X"c08c08ff",
X"a8050883",
X"c0800c9c",
X"3d0d83c0",
X"8c0c04f3",
X"3d0d02bf",
X"05330284",
X"0580c305",
X"3383cb90",
X"335a5b59",
X"79802e8d",
X"38787806",
X"5776802e",
X"8e38818a",
X"39787806",
X"5776802e",
X"81803883",
X"cb903370",
X"7a075858",
X"79883878",
X"09707906",
X"51577683",
X"cb903492",
X"983f83c0",
X"80085e80",
X"5c8f5d7d",
X"1c871133",
X"58587680",
X"2e80c238",
X"770881ec",
X"c82e0981",
X"06b73880",
X"5b815a7d",
X"1c701c9a",
X"11335959",
X"5976822e",
X"09810695",
X"3883cb90",
X"56815580",
X"54765397",
X"18335278",
X"51ffbd81",
X"3fff1a80",
X"d81c5c5a",
X"798025cf",
X"38ff1d81",
X"c41d5d5d",
X"7c8025ff",
X"a6388f3d",
X"0d04e93d",
X"0d696c02",
X"880580ea",
X"05225c5a",
X"5b807071",
X"415e58ff",
X"78797a7b",
X"7c7d464c",
X"4a45405d",
X"4362993d",
X"34620284",
X"0580dd05",
X"34777922",
X"80ffff06",
X"54457279",
X"2379782e",
X"8887387a",
X"7081055c",
X"3370842a",
X"718c0670",
X"822a5a56",
X"568306ff",
X"1b7083ff",
X"ff065c54",
X"56805475",
X"742e9138",
X"7a708105",
X"5c33ff1b",
X"7083ffff",
X"065c5454",
X"8176279b",
X"387381ff",
X"067b7081",
X"055d3355",
X"74828029",
X"05ff1b70",
X"83ffff06",
X"5c545482",
X"7627aa38",
X"7383ffff",
X"067b7081",
X"055d3370",
X"902b7207",
X"7d708105",
X"5f337098",
X"2b7207fe",
X"1f7083ff",
X"ff064052",
X"52525254",
X"547e802e",
X"80c43876",
X"86f73874",
X"8a2e0981",
X"06943881",
X"1f7081ff",
X"06811e70",
X"81ff065f",
X"52405386",
X"dc39748c",
X"2e098106",
X"86d338ff",
X"1f7081ff",
X"06ff1e70",
X"81ff065f",
X"5240537b",
X"632586bd",
X"38ff4386",
X"b8397681",
X"2e83bb38",
X"76812489",
X"3876802e",
X"8d3886a5",
X"3976822e",
X"84a63886",
X"9c39f815",
X"53728426",
X"84953872",
X"842981ef",
X"c4055372",
X"08046480",
X"2e80cd38",
X"78228380",
X"80065372",
X"8380802e",
X"098106bc",
X"38805675",
X"6427a438",
X"751e7083",
X"ffff0677",
X"101b9011",
X"72832a58",
X"51575153",
X"73753472",
X"87068171",
X"2b515372",
X"81163481",
X"167081ff",
X"06575397",
X"7627cc38",
X"7f840740",
X"800b993d",
X"43566116",
X"70337098",
X"2b70982c",
X"51515153",
X"80732480",
X"fb386073",
X"291e7083",
X"ffff067a",
X"22838080",
X"06525853",
X"72838080",
X"2e098106",
X"80de3860",
X"88327030",
X"70720780",
X"25639032",
X"70307072",
X"07802573",
X"07535458",
X"51555373",
X"802ebd38",
X"76870653",
X"72b63875",
X"84297610",
X"05791184",
X"1179832a",
X"57575153",
X"73753460",
X"81163465",
X"86142366",
X"88142375",
X"87387f81",
X"07408d39",
X"75812e09",
X"81068538",
X"7f820740",
X"81167081",
X"ff065753",
X"817627fe",
X"e5386361",
X"291e7083",
X"ffff065f",
X"53807046",
X"42ff0284",
X"0580dd05",
X"34ff0b99",
X"3d3483f5",
X"39811c70",
X"81ff065d",
X"53804273",
X"812e0981",
X"068e3877",
X"81800a29",
X"81800a05",
X"5880d339",
X"73802e89",
X"3873822e",
X"0981068d",
X"387c8180",
X"0a298180",
X"0a055da4",
X"39815f83",
X"b839ff1c",
X"7081ff06",
X"5d537b63",
X"258338ff",
X"437c802e",
X"92387c81",
X"800a2981",
X"ff0a055d",
X"7c982c5d",
X"83933977",
X"802e9238",
X"7781800a",
X"2981ff0a",
X"05587798",
X"2c5882fd",
X"39775383",
X"9e397489",
X"2680f438",
X"74842981",
X"efd80553",
X"72080473",
X"872e82e1",
X"3873852e",
X"82db3873",
X"882e82d5",
X"38738c2e",
X"82cf3873",
X"892e0981",
X"06863881",
X"4582c239",
X"73812e09",
X"810682b9",
X"38628025",
X"82b3387b",
X"982b7098",
X"2c514382",
X"a8397383",
X"ffff0646",
X"829f3973",
X"83ffff06",
X"47829639",
X"7381ff06",
X"41828e39",
X"73811a34",
X"82873973",
X"81ff0644",
X"81ff397e",
X"5382a039",
X"74812e81",
X"e3387481",
X"24893874",
X"802e8d38",
X"81e73974",
X"822e81d8",
X"3881de39",
X"74567b83",
X"38815674",
X"5373862e",
X"09810697",
X"38758106",
X"5372802e",
X"8e387822",
X"82ffff06",
X"fe808007",
X"53b6397b",
X"83388153",
X"73822e09",
X"81069738",
X"72810653",
X"72802e8e",
X"38782281",
X"ffff0681",
X"80800753",
X"93397b96",
X"38fc1453",
X"7281268e",
X"387822ff",
X"80800753",
X"72792380",
X"e5398055",
X"73812e09",
X"81068338",
X"73557753",
X"77802e89",
X"38748106",
X"537280ca",
X"3872d015",
X"54557281",
X"26833881",
X"5577802e",
X"b9387481",
X"06537280",
X"2eb03878",
X"22838080",
X"06537283",
X"80802e09",
X"81069f38",
X"73b02e09",
X"81068738",
X"61993d34",
X"913973b1",
X"2e098106",
X"89386102",
X"840580dd",
X"05346181",
X"05538c39",
X"61743181",
X"05538439",
X"61145372",
X"83ffff06",
X"4279f7fb",
X"387d832a",
X"5372821a",
X"34782283",
X"80800653",
X"72838080",
X"2e098106",
X"88388153",
X"7f872e83",
X"38805372",
X"83c0800c",
X"993d0d04",
X"fd3d0d75",
X"83113382",
X"12337198",
X"2b71902b",
X"07811433",
X"70882b72",
X"07753371",
X"0783c080",
X"0c525354",
X"56545285",
X"3d0d04f6",
X"3d0d02b7",
X"05330284",
X"05bb0533",
X"028805bf",
X"05335b5b",
X"5b805880",
X"5778882b",
X"7a075680",
X"557a5481",
X"53a3527c",
X"5192cc3f",
X"83c08008",
X"81ff0683",
X"c0800c8c",
X"3d0d04f6",
X"3d0d02b7",
X"05330284",
X"05bb0533",
X"028805bf",
X"05335b5b",
X"5b805880",
X"5778882b",
X"7a075680",
X"557a5483",
X"53a3527c",
X"5192903f",
X"83c08008",
X"81ff0683",
X"c0800c8c",
X"3d0d04f7",
X"3d0d02b3",
X"05330284",
X"05b60522",
X"605a5856",
X"80558054",
X"805381a3",
X"527b5191",
X"e23f83c0",
X"800881ff",
X"0683c080",
X"0c8b3d0d",
X"04ee3d0d",
X"6490115c",
X"5c807b34",
X"800b841c",
X"0c800b88",
X"1c34810b",
X"891c3488",
X"0b8a1c34",
X"800b8b1c",
X"34881b08",
X"c1068107",
X"881c0c8f",
X"3d70545d",
X"88527b51",
X"9c923f83",
X"c0800881",
X"ff06705b",
X"597881a9",
X"38903d33",
X"5e81db5a",
X"7d892e09",
X"81068199",
X"387c5392",
X"527b519b",
X"eb3f83c0",
X"800881ff",
X"06705b59",
X"78818238",
X"7c588857",
X"7856a955",
X"78548653",
X"81a0527b",
X"5190d03f",
X"83c08008",
X"81ff0670",
X"5b597880",
X"e03802ba",
X"05337b34",
X"7c547853",
X"7d527b51",
X"9bd33f83",
X"c0800881",
X"ff06705b",
X"597880c1",
X"3802bd05",
X"33527b51",
X"9beb3f83",
X"c0800881",
X"ff06705b",
X"5978aa38",
X"817b335a",
X"5a797926",
X"99388054",
X"79538852",
X"7b51fdbb",
X"3f811a70",
X"81ff067c",
X"33525b59",
X"e439810b",
X"881c3480",
X"5a7983c0",
X"800c943d",
X"0d04800b",
X"83c0800c",
X"04f93d0d",
X"79028405",
X"ab05338e",
X"3d705458",
X"5858ffaf",
X"ec3f8a3d",
X"8a0551ff",
X"afe33f75",
X"51fc8d3f",
X"83c08008",
X"8486812e",
X"be3883c0",
X"80088486",
X"81269938",
X"83c08008",
X"8482802e",
X"80e63883",
X"c0800884",
X"82812e9f",
X"3881b439",
X"83c08008",
X"80c08283",
X"2e80f438",
X"83c08008",
X"80c08683",
X"2e80e838",
X"81993983",
X"c09c3355",
X"80567476",
X"2e098106",
X"818b3874",
X"54765391",
X"527751fb",
X"d63f7454",
X"76539052",
X"7751fbcb",
X"3f745476",
X"53845277",
X"51fbfc3f",
X"810b83c0",
X"9c3481b1",
X"5680de39",
X"80547653",
X"91527751",
X"fba93f80",
X"54765390",
X"527751fb",
X"9e3f800b",
X"83c09c34",
X"76528718",
X"33519796",
X"3fb53980",
X"54765394",
X"527751fb",
X"823f8054",
X"76539052",
X"7751faf7",
X"3f7551ff",
X"ae973f83",
X"c0800889",
X"2a810653",
X"76528718",
X"335190cd",
X"3f800b83",
X"c09c3480",
X"567583c0",
X"800c893d",
X"0d04f23d",
X"0d609011",
X"5a58800b",
X"881a3371",
X"59565674",
X"762e82a5",
X"3882ac3f",
X"84190883",
X"c0800826",
X"82953878",
X"335a810b",
X"8e3d2390",
X"3df81155",
X"f4055399",
X"18527751",
X"8ae53f83",
X"c0800881",
X"ff067057",
X"5574772e",
X"09810681",
X"d9388639",
X"745681d2",
X"39815682",
X"578e3d33",
X"77065574",
X"802ebb38",
X"800b8d3d",
X"34903df0",
X"05548453",
X"75527751",
X"facd3f83",
X"c0800881",
X"ff065574",
X"9d387b53",
X"75527751",
X"fce73f83",
X"c0800881",
X"ff065574",
X"81b12e81",
X"8b3874ff",
X"b3387610",
X"81fc0681",
X"177081ff",
X"06585657",
X"877627ff",
X"a8388156",
X"757a2680",
X"eb38800b",
X"8d3d348c",
X"3d705557",
X"84537552",
X"7751f9f7",
X"3f83c080",
X"0881ff06",
X"557480c1",
X"387651ff",
X"ac933f83",
X"c0800882",
X"87065574",
X"82812e09",
X"8106aa38",
X"02ae0533",
X"81075574",
X"028405ae",
X"05347b53",
X"75527751",
X"fbeb3f83",
X"c0800881",
X"ff065574",
X"81b12e90",
X"3874feb8",
X"38811670",
X"81ff0657",
X"55ff9139",
X"80567581",
X"ff065697",
X"3f83c080",
X"088fd005",
X"841a0c75",
X"577683c0",
X"800c903d",
X"0d040490",
X"80a00883",
X"c0800c04",
X"ff3d0d73",
X"87e82951",
X"fefdaf3f",
X"833d0d04",
X"0483cb94",
X"0b83c080",
X"0c04fd3d",
X"0d757754",
X"54800b83",
X"caf43472",
X"8a389090",
X"800b8415",
X"0c903972",
X"812e0981",
X"06883890",
X"98800b84",
X"150c8414",
X"0883cb8c",
X"0c800b88",
X"150c800b",
X"8c150c83",
X"cb8c0853",
X"820b8780",
X"14348151",
X"ff9e3f83",
X"cb8c0853",
X"800b8814",
X"3483cb8c",
X"0853810b",
X"87801434",
X"83cb8c08",
X"53800b8c",
X"143483cb",
X"8c085380",
X"0ba41434",
X"91743480",
X"0b83c0a0",
X"34800b83",
X"c0a43480",
X"0b83c0a8",
X"34805473",
X"81c42983",
X"cb980553",
X"800b8314",
X"34811470",
X"81ff0655",
X"538f7427",
X"e638853d",
X"0d04fe3d",
X"0d747682",
X"113370bf",
X"0681712b",
X"ff055651",
X"51525390",
X"71278338",
X"ff527651",
X"71712383",
X"cb8c0851",
X"87133390",
X"1234800b",
X"83c0a434",
X"800b83c0",
X"a8348813",
X"338a1433",
X"52527180",
X"2eaa3870",
X"81ff0651",
X"84527083",
X"38705271",
X"83c0a434",
X"8a133370",
X"30708025",
X"842b7088",
X"07515152",
X"537083c0",
X"a8349039",
X"7081ff06",
X"51708338",
X"98527183",
X"c0a83480",
X"0b83c080",
X"0c843d0d",
X"04f13d0d",
X"61656802",
X"8c0580cb",
X"05330290",
X"0580ce05",
X"22029405",
X"80d60522",
X"4240415a",
X"4040fd8b",
X"3f83c080",
X"08a78805",
X"5b807071",
X"5b5b5283",
X"943983cb",
X"8c08517d",
X"94123483",
X"c0a43381",
X"07558070",
X"54567f86",
X"2680ea38",
X"7f842981",
X"f08c0583",
X"cb8c0853",
X"51700804",
X"800b8413",
X"34a13977",
X"33703070",
X"80258371",
X"31515152",
X"53708413",
X"348d3981",
X"0b841334",
X"b839830b",
X"84133481",
X"705456ad",
X"39810b84",
X"1334a239",
X"77337030",
X"70802583",
X"71315151",
X"52537084",
X"13348078",
X"33525270",
X"83388152",
X"71783481",
X"53748807",
X"5583c0a8",
X"3383cb8c",
X"08525781",
X"0b81d012",
X"3483cb8c",
X"0851810b",
X"81901234",
X"7e802eae",
X"3872802e",
X"a9387eff",
X"1e525470",
X"83ffff06",
X"537283ff",
X"ff2e9738",
X"73708105",
X"553383cb",
X"8c085351",
X"7081c013",
X"34ff1351",
X"de3983cb",
X"8c08a811",
X"33535176",
X"88123483",
X"cb8c0851",
X"74713481",
X"ff529139",
X"83cb8c08",
X"a0113370",
X"81065152",
X"53708f38",
X"fafd3f7a",
X"83c08008",
X"26e63881",
X"8839810b",
X"a0143483",
X"cb8c08a8",
X"113380ff",
X"06707807",
X"52535170",
X"802e80ed",
X"3871862a",
X"70810651",
X"5170802e",
X"91388078",
X"33525370",
X"83388153",
X"72783480",
X"e0397184",
X"2a708106",
X"51517080",
X"2e9b3881",
X"197083ff",
X"ff067d30",
X"709f2a51",
X"525a5178",
X"7c2e0981",
X"06af38a4",
X"3971832a",
X"70810651",
X"5170802e",
X"9338811a",
X"7081ff06",
X"5b517983",
X"2e098106",
X"90388a39",
X"71a30651",
X"70802e85",
X"38715192",
X"39f9e43f",
X"7a83c080",
X"0826fce2",
X"387181bf",
X"06517083",
X"c0800c91",
X"3d0d04f6",
X"3d0d02b3",
X"05330284",
X"05b70533",
X"028805ba",
X"05225959",
X"59800b8c",
X"3d348c3d",
X"fc055680",
X"55805476",
X"53775278",
X"51fbf23f",
X"83c08008",
X"81ff0683",
X"c0800c8c",
X"3d0d04f3",
X"3d0d7f62",
X"64028c05",
X"80c20522",
X"72228115",
X"33425f41",
X"5e595980",
X"78237d53",
X"78335281",
X"51ffa03f",
X"83c08008",
X"81ff0656",
X"75802e86",
X"38755481",
X"ad3983cb",
X"8c08a811",
X"33821b33",
X"70862a70",
X"81067398",
X"2b535157",
X"5c565779",
X"80258338",
X"81567376",
X"2e873881",
X"f0548182",
X"39818c17",
X"337081ff",
X"0679227d",
X"7131902b",
X"70902c70",
X"09709f2c",
X"72067052",
X"52535153",
X"57575475",
X"74248338",
X"75557484",
X"808029fc",
X"80800570",
X"902c5155",
X"74ff2e94",
X"3883cb8c",
X"08818011",
X"33515473",
X"7c708105",
X"5e34db39",
X"77227605",
X"54737823",
X"7909709f",
X"2a708106",
X"821c3381",
X"bf067186",
X"2b075151",
X"51547382",
X"1a347c76",
X"268a3877",
X"22547a74",
X"26febb38",
X"80547383",
X"c0800c8f",
X"3d0d04f9",
X"3d0d7a57",
X"800b893d",
X"23893dfc",
X"05537652",
X"7951f8da",
X"3f83c080",
X"0881ff06",
X"70575574",
X"96387c54",
X"7b53883d",
X"22527651",
X"fde53f83",
X"c0800881",
X"ff065675",
X"83c0800c",
X"893d0d04",
X"f03d0d62",
X"66028805",
X"80ce0522",
X"415d5e80",
X"02840580",
X"d205227f",
X"810533ff",
X"115a5d5a",
X"5d81da58",
X"76bf2680",
X"e9387880",
X"2e80e138",
X"7a58787b",
X"27833878",
X"58821e33",
X"70872a58",
X"5a76923d",
X"34923dfc",
X"05567755",
X"7b547e53",
X"7d335282",
X"51f8de3f",
X"83c08008",
X"81ff065d",
X"800b923d",
X"33585a76",
X"802e8338",
X"815a821e",
X"3380ff06",
X"7a872b07",
X"5776821f",
X"347c9138",
X"78783170",
X"83ffff06",
X"791e5e5a",
X"57ff9b39",
X"7c587783",
X"c0800c92",
X"3d0d04f8",
X"3d0d7b02",
X"8405b205",
X"22585880",
X"0b8a3d23",
X"8a3dfc05",
X"5377527a",
X"51f6f73f",
X"83c08008",
X"81ff0670",
X"57557496",
X"387d5476",
X"53893d22",
X"527751fe",
X"af3f83c0",
X"800881ff",
X"06567583",
X"c0800c8a",
X"3d0d04ec",
X"3d0d666e",
X"02880580",
X"df053302",
X"8c0580e3",
X"05330290",
X"0580e705",
X"33029405",
X"80eb0533",
X"02980580",
X"ee052241",
X"43415f5c",
X"40570280",
X"f2052296",
X"3d23963d",
X"f0055384",
X"17705377",
X"5259f686",
X"3f83c080",
X"0881ff06",
X"587781e5",
X"38777a81",
X"80065840",
X"80772583",
X"38814079",
X"943d347b",
X"02840580",
X"c905347c",
X"02840580",
X"ca05347d",
X"02840580",
X"cb05347a",
X"953d347a",
X"882a5776",
X"02840580",
X"cd053495",
X"3d225776",
X"02840580",
X"ce053476",
X"882a5776",
X"02840580",
X"cf053477",
X"923d3496",
X"3dec1157",
X"578855f4",
X"1754923d",
X"22537752",
X"7751f695",
X"3f83c080",
X"0881ff06",
X"587780ed",
X"387e802e",
X"80cb3892",
X"3d227908",
X"58587f80",
X"2e9c3876",
X"81808007",
X"790c7e54",
X"963dfc05",
X"537783ff",
X"ff065278",
X"51f9fc3f",
X"99397682",
X"80800779",
X"0c7e5495",
X"3d225377",
X"83ffff06",
X"527851fc",
X"8f3f83c0",
X"800881ff",
X"0658779d",
X"38923d22",
X"5380527f",
X"30708025",
X"84713153",
X"5157f987",
X"3f83c080",
X"0881ff06",
X"587783c0",
X"800c963d",
X"0d04f63d",
X"0d7c0284",
X"05b70533",
X"5b5b8058",
X"80578056",
X"80557954",
X"85538052",
X"7a51fda3",
X"3f83c080",
X"0881ff06",
X"59788538",
X"79871c34",
X"7883c080",
X"0c8c3d0d",
X"04f93d0d",
X"02a70533",
X"028405ab",
X"05330288",
X"05af0533",
X"58595780",
X"0b83cb9b",
X"33545472",
X"742e9f38",
X"81147081",
X"ff065553",
X"738f2681",
X"b6387381",
X"c42983cb",
X"98058311",
X"33515372",
X"e3387381",
X"c42983cb",
X"94055580",
X"0b871634",
X"76881634",
X"758a1634",
X"77891634",
X"80750c83",
X"cb8c088c",
X"160c800b",
X"84163488",
X"0b851634",
X"800b8616",
X"34841508",
X"ffa1ff06",
X"a0800784",
X"160c8114",
X"7081ff06",
X"53537451",
X"febc3f83",
X"c0800881",
X"ff067055",
X"537280cd",
X"388a3973",
X"08750c72",
X"5480c239",
X"7281f7ac",
X"555681f7",
X"ac08802e",
X"b2387584",
X"29147008",
X"76537008",
X"51545472",
X"2d83c080",
X"0881ff06",
X"5372802e",
X"ce388116",
X"7081ff06",
X"81f7ac71",
X"84291153",
X"56575372",
X"08d03880",
X"547383c0",
X"800c893d",
X"0d04f93d",
X"0d795780",
X"0b841808",
X"83cb8c0c",
X"58f0883f",
X"88170883",
X"c0800827",
X"83ed38ef",
X"fa3f83c0",
X"80088105",
X"88180c83",
X"cb8c08b8",
X"11337081",
X"ff065151",
X"5473812e",
X"a4387381",
X"24883873",
X"782e8a38",
X"b8397382",
X"2e9538b1",
X"39763381",
X"f0065473",
X"902ea638",
X"917734a1",
X"39735876",
X"3381f006",
X"5473902e",
X"09810691",
X"38efa83f",
X"83c08008",
X"81c8058c",
X"180ca077",
X"34805675",
X"81c42983",
X"cb9b1133",
X"55557380",
X"2eaa3883",
X"cb941570",
X"08565474",
X"802e9d38",
X"88150880",
X"2e96388c",
X"140883cb",
X"8c082e09",
X"81068938",
X"73518815",
X"0854732d",
X"81167081",
X"ff065754",
X"8f7627ff",
X"ba387633",
X"5473b02e",
X"81993873",
X"b0248f38",
X"73912eab",
X"3873a02e",
X"80f53882",
X"a6397380",
X"d02e81e4",
X"387380d0",
X"248b3873",
X"80c02e81",
X"9938828f",
X"39738180",
X"2e81fb38",
X"82853980",
X"567581c4",
X"2983cb98",
X"11831133",
X"56595573",
X"802ea838",
X"83cb9415",
X"70085654",
X"74802e9b",
X"388c1408",
X"83cb8c08",
X"2e098106",
X"8e387351",
X"84150854",
X"732d800b",
X"83193481",
X"167081ff",
X"0657548f",
X"7627ffb9",
X"38927734",
X"81b539ed",
X"c23f8c17",
X"0883c080",
X"082781a7",
X"38b07734",
X"81a13983",
X"cb8c0854",
X"800b8c15",
X"3483cb8c",
X"0854840b",
X"88153480",
X"c07734ed",
X"963f83c0",
X"8008b205",
X"8c180c80",
X"fa39ed87",
X"3f8c1708",
X"83c08008",
X"2780ec38",
X"83cb8c08",
X"54810b8c",
X"153483cb",
X"8c085480",
X"0b881534",
X"83cb8c08",
X"54880ba0",
X"1534ecdb",
X"3f83c080",
X"0894058c",
X"180c80d0",
X"7734bc39",
X"83cb8c08",
X"a0113370",
X"832a7081",
X"06515155",
X"5573802e",
X"a638880b",
X"a01634ec",
X"ae3f8c17",
X"0883c080",
X"08279438",
X"ff807734",
X"8e397753",
X"80528051",
X"fa8b3fff",
X"90773483",
X"cb8c08a0",
X"11337083",
X"2a708106",
X"51515555",
X"73802e86",
X"38880ba0",
X"1634893d",
X"0d04f43d",
X"0d02bb05",
X"33028405",
X"bf05335d",
X"5d800b83",
X"cb980b83",
X"cb940b8c",
X"11727188",
X"14755c5a",
X"5b5f5c59",
X"5b588315",
X"33537280",
X"2e818838",
X"7333537c",
X"732e0981",
X"0680fc38",
X"81143353",
X"7b732e09",
X"810680ef",
X"38750883",
X"cb8c082e",
X"09810680",
X"e2388056",
X"7581c429",
X"83cb9c11",
X"7033831e",
X"335b5755",
X"5374782e",
X"09810697",
X"3883cba0",
X"13087908",
X"2e098106",
X"8a388114",
X"33527451",
X"fef83f81",
X"167081ff",
X"0657538f",
X"7627c538",
X"80770854",
X"5472742e",
X"91387651",
X"84130853",
X"722d83c0",
X"800881ff",
X"0654800b",
X"831b3473",
X"53a93981",
X"1881c416",
X"81c41681",
X"c41981c4",
X"1f81c41e",
X"81c41d60",
X"81c40541",
X"5d5e5f59",
X"5656588f",
X"7825feca",
X"38805372",
X"83c0800c",
X"8e3d0d04",
X"f83d0d02",
X"ae05227d",
X"59578056",
X"81558054",
X"86538180",
X"527a51f4",
X"ee3f83c0",
X"800881ff",
X"0683c080",
X"0c8a3d0d",
X"04f73d0d",
X"02b20522",
X"028405b7",
X"0533605a",
X"5b578056",
X"82557954",
X"86538180",
X"527b51f4",
X"be3f83c0",
X"800881ff",
X"0683c080",
X"0c8b3d0d",
X"04f83d0d",
X"02af0533",
X"59805880",
X"57805680",
X"55785489",
X"5380527a",
X"51f4943f",
X"83c08008",
X"81ff0683",
X"c0800c8a",
X"3d0d04ff",
X"b83d0d80",
X"cb3d0870",
X"5381f3e8",
X"5256feaa",
X"c93f83c0",
X"800880f3",
X"387551fe",
X"a4b43f83",
X"ffff0b83",
X"c0800825",
X"80e13875",
X"51fea4b3",
X"3f83c080",
X"085583c0",
X"800880cf",
X"38828053",
X"83c08008",
X"528a3d70",
X"5257fee6",
X"8a3f7452",
X"7551fea3",
X"c43f8059",
X"80ca3dfd",
X"fc055482",
X"80537652",
X"7551fea1",
X"cb3f8115",
X"55748880",
X"2e098106",
X"e1388052",
X"7551fea3",
X"9c3f800b",
X"83e3d80c",
X"7583e3d4",
X"0c873980",
X"0b83e3d4",
X"0c80ca3d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04ffb8",
X"3d0d80cb",
X"3d707084",
X"05520858",
X"5683e3d4",
X"08802e80",
X"fa388a3d",
X"705a7655",
X"775481e9",
X"de5380cb",
X"3dfdfc05",
X"5255fecf",
X"da3f8052",
X"80ca3dfd",
X"fc0551ff",
X"ad3f83e3",
X"d8085283",
X"e3d40851",
X"fea2a23f",
X"80587451",
X"fecda03f",
X"80ca3dfd",
X"f8055483",
X"c0800853",
X"745283e3",
X"d40851fe",
X"a09e3f83",
X"e3d80818",
X"83e3d80c",
X"80ca3dfd",
X"f8055481",
X"5381f3f4",
X"5283e3d4",
X"0851fe9f",
X"ff3f83e3",
X"d8081883",
X"e3d80c80",
X"ca3d0d04",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002d46",
X"00002d87",
X"00002da9",
X"00002dcb",
X"00002df1",
X"00002df1",
X"00002df1",
X"00002df1",
X"00002e62",
X"00002eb3",
X"00002ebd",
X"000044a5",
X"00004ec5",
X"00004f8e",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3f00",
X"0c0c4000",
X"0a0a4100",
X"0b0b4100",
X"07074100",
X"0a0b4300",
X"080b4200",
X"06060004",
X"04044500",
X"05054400",
X"0e0f2900",
X"08080004",
X"09090004",
X"0a0f4300",
X"090f4200",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"00006172",
X"00006479",
X"00006285",
X"00006479",
X"000062c2",
X"00006313",
X"00006352",
X"0000635b",
X"00006479",
X"00006479",
X"00006479",
X"00006479",
X"00006364",
X"0000636c",
X"00006373",
X"00006579",
X"00006672",
X"00006786",
X"00006a7c",
X"00006a97",
X"00006a83",
X"00006a97",
X"00006a9e",
X"00006aa9",
X"00006ab0",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"25782e48",
X"75622e20",
X"25642070",
X"6f727473",
X"00000000",
X"25782e48",
X"49440000",
X"204d6f75",
X"73650000",
X"204b6579",
X"626f6172",
X"64000000",
X"204a6f79",
X"73746963",
X"6b3a2564",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"43505520",
X"54757262",
X"6f3a2564",
X"78000000",
X"44726976",
X"65205475",
X"72626f3a",
X"25730000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"526f7461",
X"74652055",
X"5342206a",
X"6f797374",
X"69636b73",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"66726565",
X"7a65722e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"4d454d00",
X"5374616e",
X"64617264",
X"00000000",
X"46617374",
X"28362900",
X"46617374",
X"28352900",
X"46617374",
X"28342900",
X"46617374",
X"28332900",
X"46617374",
X"28322900",
X"46617374",
X"28312900",
X"46617374",
X"28302900",
X"2f757362",
X"2e6c6f67",
X"00000000",
X"0a000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"000078a8",
X"000078ac",
X"000078b4",
X"000078c0",
X"000078cc",
X"000078d8",
X"000078e4",
X"000078e8",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00000028",
X"00000006",
X"00000005",
X"00000004",
X"00000003",
X"00000002",
X"00000001",
X"00000000",
X"000079a4",
X"000079b0",
X"000079b8",
X"000079c0",
X"000079c8",
X"000079d0",
X"000079d8",
X"000079e0",
X"00007800",
X"00007648",
X"00000000",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
