
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80de",
X"c4738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80e1",
X"a40c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580d8",
X"f22d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580d786",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"96bf0480",
X"3d0d80e2",
X"cc087008",
X"810683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d80e2",
X"cc087008",
X"70fe0676",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80e2cc08",
X"70087081",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80e2cc08",
X"700870fd",
X"06761007",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"e2cc0870",
X"0870822c",
X"bf0683e0",
X"800c5151",
X"823d0d04",
X"ff3d0d80",
X"e2cc0870",
X"0870fe83",
X"0676822b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80e2cc08",
X"70087088",
X"2c870683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80e2cc08",
X"700870f1",
X"ff067688",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d80e2cc",
X"08700870",
X"8b2cbf06",
X"83e0800c",
X"5151823d",
X"0d04ff3d",
X"0d80e2cc",
X"08700870",
X"f88fff06",
X"768b2b07",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"e2dc0870",
X"0870882c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"e2dc0870",
X"0870892c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"e2dc0870",
X"08708a2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"e2dc0870",
X"08708b2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"fd3d0d75",
X"81e62987",
X"2a80e2bc",
X"0854730c",
X"853d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d818080",
X"53805288",
X"800a51ff",
X"b33fa080",
X"53805282",
X"800a51c7",
X"3f843d0d",
X"04803d0d",
X"8151fccf",
X"3f72802e",
X"8338d33f",
X"8151fcf1",
X"3f8051fc",
X"ec3f8051",
X"fcb93f82",
X"3d0d04fd",
X"3d0d7552",
X"805480ff",
X"72258838",
X"810bff80",
X"135354ff",
X"bf125170",
X"99268638",
X"e012529e",
X"39ff9f12",
X"51997127",
X"9538d012",
X"e0137054",
X"54518971",
X"2788388f",
X"73278338",
X"80527380",
X"2e853881",
X"80125271",
X"81ff0683",
X"e0800c85",
X"3d0d0480",
X"3d0d84d8",
X"c0518071",
X"70810553",
X"347084e0",
X"c02e0981",
X"06f03882",
X"3d0d04fe",
X"3d0d0297",
X"053351ff",
X"863f83e0",
X"800881ff",
X"0683e09c",
X"08545280",
X"73249b38",
X"83e0b808",
X"137283e0",
X"bc080753",
X"53717334",
X"83e09c08",
X"810583e0",
X"9c0c843d",
X"0d04fa3d",
X"0d82800a",
X"1b558057",
X"883dfc05",
X"54795374",
X"527851a2",
X"cf3f883d",
X"0d04fe3d",
X"0d83e0b0",
X"08527451",
X"a9e33f83",
X"e080088c",
X"38765375",
X"5283e0b0",
X"0851c73f",
X"843d0d04",
X"fe3d0d83",
X"e0b00853",
X"75527451",
X"a3f13f83",
X"e080088d",
X"38775376",
X"5283e0b0",
X"0851ffa2",
X"3f843d0d",
X"04fd3d0d",
X"83e0b408",
X"51a2e53f",
X"83e08008",
X"90802e09",
X"8106ad38",
X"805483c1",
X"80805383",
X"e0800852",
X"83e0b408",
X"51fef33f",
X"87c18080",
X"143387c1",
X"90801534",
X"81145473",
X"90802e09",
X"8106e938",
X"853d0d04",
X"0b0b80df",
X"940b83e0",
X"800c04f7",
X"3d0d805a",
X"80598058",
X"80705757",
X"fde53f80",
X"0b83e09c",
X"0c800b83",
X"e0bc0c0b",
X"0b80df98",
X"519dc73f",
X"81800b83",
X"e0bc0c0b",
X"0b80df9c",
X"519db73f",
X"80d00b83",
X"e09c0c75",
X"30707707",
X"80257087",
X"2b83e0bc",
X"0c5154f9",
X"cb3f83e0",
X"8008520b",
X"0b80dfa4",
X"519d8f3f",
X"80f80b83",
X"e09c0c75",
X"81327030",
X"70720780",
X"2570872b",
X"83e0bc0c",
X"515555fe",
X"fb3f83e0",
X"8008520b",
X"0b80dfb0",
X"519ce33f",
X"81a00b83",
X"e09c0c75",
X"82327030",
X"70720780",
X"2570872b",
X"83e0bc0c",
X"515583e0",
X"b4085255",
X"9dfd3f83",
X"e0800852",
X"0b0b80df",
X"b8519cb2",
X"3f81c80b",
X"83e09c0c",
X"75833270",
X"30707207",
X"80257087",
X"2b83e0bc",
X"0c51550b",
X"0b80dfc0",
X"52559c8e",
X"3f81f00b",
X"83e09c0c",
X"75843270",
X"30707207",
X"80257087",
X"2b83e0bc",
X"0c51550b",
X"0b80dfd0",
X"52559bea",
X"3f82980b",
X"83e09c0c",
X"75853270",
X"30707207",
X"80257087",
X"2b83e0bc",
X"0c51550b",
X"0b80dfe8",
X"52559bc6",
X"3f82c00b",
X"83e09c0c",
X"75863270",
X"30707207",
X"80257087",
X"2b83e0bc",
X"0c51550b",
X"0b80e080",
X"52559ba2",
X"3f868da0",
X"51f9bd3f",
X"8052883d",
X"7052548a",
X"ef3f8352",
X"73518ae8",
X"3f781656",
X"75802585",
X"38805690",
X"39867625",
X"85388656",
X"87397586",
X"2682c938",
X"75842980",
X"ded40554",
X"730804f7",
X"8f3f83e0",
X"80087856",
X"5474812e",
X"09810689",
X"3883e080",
X"08105490",
X"3974ff2e",
X"09810688",
X"3883e080",
X"08812c54",
X"90742585",
X"38905488",
X"39738024",
X"83388154",
X"7351f6ec",
X"3f81fd39",
X"f6ff3f83",
X"e0800818",
X"54738025",
X"85388054",
X"88398774",
X"25833887",
X"547351f6",
X"fc3f81dc",
X"39778738",
X"79802e81",
X"d3389fbf",
X"0b83e0d0",
X"0c83e0b4",
X"08518cad",
X"3ffbaa3f",
X"81be3979",
X"802e81b8",
X"389ff00b",
X"83e0d00c",
X"83e0b008",
X"518c923f",
X"75832e09",
X"81069438",
X"81808053",
X"82808052",
X"83e0b008",
X"51fa973f",
X"81873975",
X"842e0981",
X"06af3882",
X"80805381",
X"80805283",
X"e0b00851",
X"f9fc3f80",
X"54848280",
X"80143384",
X"81808015",
X"34811454",
X"73818080",
X"2e098106",
X"e83880d1",
X"3975852e",
X"09810680",
X"c8388054",
X"81808053",
X"80c08052",
X"83e0b008",
X"51f9c33f",
X"82808053",
X"80c08052",
X"83e0b008",
X"51f9b33f",
X"84818080",
X"14338481",
X"c0801534",
X"84828080",
X"14338482",
X"c0801534",
X"81145473",
X"80c0802e",
X"098106dc",
X"3881548c",
X"39798738",
X"76802efa",
X"c3388054",
X"7383e080",
X"0c8b3d0d",
X"04ff3d0d",
X"f5d23f83",
X"e0800880",
X"2e863880",
X"5180dd39",
X"f5da3f83",
X"e0800880",
X"d138f680",
X"3f83e080",
X"08802eaa",
X"388151f3",
X"d23f82f7",
X"3f800b83",
X"e09c0cf9",
X"f23f83e0",
X"800852ff",
X"0b83e09c",
X"0c85963f",
X"71a43871",
X"51f3b03f",
X"a239f5b4",
X"3f83e080",
X"08802e97",
X"388151f3",
X"9e3f82c3",
X"3fff0b83",
X"e09c0c84",
X"f03f8151",
X"f6b73f83",
X"3d0d0483",
X"e08c0802",
X"83e08c0c",
X"fa3d0d80",
X"0b83e0a0",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"f8050c9b",
X"d03f83e0",
X"80088605",
X"fc0683e0",
X"8c08f405",
X"0c0283e0",
X"8c08f405",
X"08310d85",
X"3d7083e0",
X"8c08fc05",
X"08708405",
X"83e08c08",
X"fc050c0c",
X"51989a3f",
X"83e08c08",
X"f8050881",
X"0583e08c",
X"08f8050c",
X"83e08c08",
X"f8050886",
X"2e098106",
X"ffad3886",
X"94808051",
X"819f3fff",
X"0b83e09c",
X"0c800b83",
X"e0bc0c84",
X"d8c00b83",
X"e0b80c81",
X"51f1f43f",
X"8151f29d",
X"3f8051f2",
X"983f8151",
X"f2c23f81",
X"51f39f3f",
X"8251f2e9",
X"3f8e8352",
X"805195df",
X"3f908080",
X"52868480",
X"80519bb9",
X"3f83e080",
X"0880c838",
X"80e2e051",
X"a0ad3f83",
X"e0800883",
X"e0b40854",
X"0b0b80e0",
X"8c5383e0",
X"80085283",
X"e08c08f4",
X"050c9acf",
X"3f83e080",
X"088438f6",
X"ec3f8180",
X"80548280",
X"80530b0b",
X"80e08852",
X"83e08c08",
X"f4050851",
X"f6ae3f81",
X"51f49e3f",
X"fcf33ffc",
X"397183e0",
X"c40c8880",
X"800b83e0",
X"c00c8480",
X"800b83e0",
X"c80c04f0",
X"3d0d8380",
X"805683e0",
X"c4081683",
X"e0c00817",
X"56547433",
X"743483e0",
X"c8081654",
X"80743481",
X"16567583",
X"80a02e09",
X"8106db38",
X"83d08056",
X"83e0c408",
X"1683e0c0",
X"08175654",
X"74337434",
X"83e0c808",
X"16548074",
X"34811656",
X"7583d0a0",
X"2e098106",
X"db3883a8",
X"805683e0",
X"c4081683",
X"e0c00817",
X"56547433",
X"743483e0",
X"c8081654",
X"80743481",
X"16567583",
X"a8902e09",
X"8106db38",
X"805683e0",
X"c4081683",
X"e0c80817",
X"55557333",
X"75348116",
X"56758180",
X"802e0981",
X"06e438f3",
X"d63f893d",
X"58a25380",
X"def05277",
X"5180c387",
X"3f80578c",
X"805683e0",
X"c8081677",
X"19555573",
X"33753481",
X"16811858",
X"5676a22e",
X"098106e6",
X"3880e1bc",
X"08548674",
X"3480e1c0",
X"08548074",
X"3480e1f0",
X"08548074",
X"3480e1e0",
X"0854af74",
X"3480e1ec",
X"0854bf74",
X"3480e1e8",
X"08548074",
X"3480e1e4",
X"08549f74",
X"3480e1dc",
X"08548074",
X"3480e1cc",
X"0854f874",
X"3480e1c4",
X"08547674",
X"3480e1b4",
X"08548274",
X"3480e1c8",
X"08548274",
X"34923d0d",
X"04fe3d0d",
X"805383e0",
X"c8081383",
X"e0c40814",
X"52527033",
X"72348113",
X"53728180",
X"802e0981",
X"06e43883",
X"80805383",
X"e0c80813",
X"83e0c408",
X"14525270",
X"33723481",
X"13537283",
X"80a02e09",
X"8106e438",
X"83d08053",
X"83e0c808",
X"1383e0c4",
X"08145252",
X"70337234",
X"81135372",
X"83d0a02e",
X"098106e4",
X"3883a880",
X"5383e0c8",
X"081383e0",
X"c4081452",
X"52703372",
X"34811353",
X"7283a890",
X"2e098106",
X"e438843d",
X"0d04fd3d",
X"0d755480",
X"740c800b",
X"84150c80",
X"0b88150c",
X"80e1b008",
X"703380e1",
X"b4087033",
X"70822a70",
X"81067030",
X"70720770",
X"09709f2c",
X"78069e06",
X"54515154",
X"51515552",
X"54518072",
X"98065253",
X"70882e09",
X"81068338",
X"81537098",
X"32703070",
X"80257571",
X"3184180c",
X"51515180",
X"72860652",
X"5370822e",
X"09810683",
X"38815370",
X"86327030",
X"70802575",
X"7131770c",
X"51515171",
X"94327030",
X"70802588",
X"170c5151",
X"853d0d04",
X"fe3d0d74",
X"76545271",
X"51fee73f",
X"72812ea2",
X"38817326",
X"8d387282",
X"2eab3872",
X"832e9f38",
X"e6397108",
X"e2388412",
X"08dd3888",
X"1208d838",
X"a0398812",
X"08812e09",
X"8106cc38",
X"94398812",
X"08812e8d",
X"38710889",
X"38841208",
X"802effb7",
X"38843d0d",
X"04fc3d0d",
X"76705255",
X"b5d73f83",
X"e0800815",
X"ff055473",
X"752e8e38",
X"73335372",
X"ae2e8638",
X"ff1454ef",
X"39775281",
X"1451b4ef",
X"3f83e080",
X"08307083",
X"e0800807",
X"802583e0",
X"800c5386",
X"3d0d04fb",
X"3d0d7770",
X"52569acd",
X"3f83e080",
X"08558154",
X"83e08008",
X"80cc3875",
X"519a903f",
X"83e08008",
X"80e0a453",
X"83e08008",
X"5254ff91",
X"3f83e080",
X"08a13880",
X"e0a85273",
X"51ff823f",
X"83e08008",
X"923880e0",
X"ac527351",
X"fef33f83",
X"e0800880",
X"2e833881",
X"55745373",
X"5280e0b0",
X"518eab3f",
X"74547383",
X"e0800c87",
X"3d0d04fd",
X"3d0d7570",
X"525499e1",
X"3f815383",
X"e0800897",
X"38735199",
X"aa3f80e0",
X"c45283e0",
X"800851fe",
X"b03f83e0",
X"80085372",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"70525499",
X"b03f8153",
X"83e08008",
X"97387351",
X"98f93f80",
X"e0c85283",
X"e0800851",
X"fdff3f83",
X"e0800853",
X"7283e080",
X"0c853d0d",
X"04e03d0d",
X"a33d0870",
X"525e8eef",
X"3f83e080",
X"0833943d",
X"56547394",
X"3880e2f0",
X"52745184",
X"b2397d52",
X"785191f1",
X"3f84bc39",
X"7d518ed7",
X"3f83e080",
X"08527451",
X"8e873f83",
X"e0d00852",
X"933d7052",
X"5d94e13f",
X"83e08008",
X"59800b83",
X"e0800855",
X"5b83e080",
X"087b2e94",
X"38811b74",
X"525b9894",
X"3f83e080",
X"085483e0",
X"8008ee38",
X"805aff7a",
X"437a427a",
X"415f7909",
X"709f2c7b",
X"065b547a",
X"7a248438",
X"ff1b5af6",
X"1a700970",
X"9f2c7206",
X"7bff125a",
X"5a525555",
X"80752595",
X"38765197",
X"d33f83e0",
X"800876ff",
X"18585557",
X"738024ed",
X"38747f2e",
X"8638ec8b",
X"3f745f78",
X"ff1b7058",
X"5d58807a",
X"25953877",
X"5197a93f",
X"83e08008",
X"76ff1858",
X"55587380",
X"24ed3880",
X"0b83e09c",
X"0c800b83",
X"e0bc0c80",
X"e0cc518b",
X"cd3f8180",
X"0b83e0bc",
X"0c80e0d4",
X"518bbf3f",
X"a80b83e0",
X"9c0c7680",
X"2e80e438",
X"83e09c08",
X"77793270",
X"30707207",
X"80257087",
X"2b83e0bc",
X"0c515678",
X"53565696",
X"e03f83e0",
X"8008802e",
X"883880e0",
X"dc518b86",
X"3f765196",
X"a23f83e0",
X"80085280",
X"dfb4518a",
X"f53f7651",
X"96aa3f83",
X"e0800883",
X"e09c0855",
X"57757425",
X"8638a816",
X"56f73975",
X"83e09c0c",
X"86f07624",
X"ff983887",
X"980b83e0",
X"9c0c7780",
X"2eb13877",
X"5195e03f",
X"83e08008",
X"78525596",
X"803f80e0",
X"e45483e0",
X"80088d38",
X"87398076",
X"34fda039",
X"80e0f854",
X"74537352",
X"80e09851",
X"8a943f80",
X"5480e1a0",
X"518a8b3f",
X"81145473",
X"a82e0981",
X"06ef3886",
X"8da051e8",
X"9b3f8052",
X"903d7052",
X"54f9cd3f",
X"83527351",
X"f9c63f61",
X"802e80fd",
X"387b5473",
X"ff2e9638",
X"78802e80",
X"fe387851",
X"958a3f83",
X"e08008ff",
X"155559e7",
X"3978802e",
X"80e93878",
X"5195863f",
X"83e08008",
X"802efc96",
X"38785194",
X"ce3f83e0",
X"80085280",
X"e0a051ad",
X"f13f83e0",
X"8008a438",
X"7c51afa9",
X"3f83e080",
X"085574ff",
X"16565480",
X"7425fc83",
X"38741d70",
X"33555673",
X"af2efed2",
X"38e83978",
X"51948e3f",
X"83e08008",
X"527c51ae",
X"e03ffbe3",
X"397f8829",
X"6010057a",
X"0561055a",
X"fc9439a2",
X"3d0d04fe",
X"3d0d80e1",
X"f8087033",
X"7081ff06",
X"70842a81",
X"32810655",
X"51525371",
X"802e8c38",
X"a8733480",
X"e1f80851",
X"b8713471",
X"83e0800c",
X"843d0d04",
X"fe3d0d80",
X"e1f80870",
X"337081ff",
X"0670852a",
X"81328106",
X"55515253",
X"71802e8c",
X"38987334",
X"80e1f808",
X"51b87134",
X"7183e080",
X"0c843d0d",
X"04803d0d",
X"80e1f408",
X"51937134",
X"80e28008",
X"51ff7134",
X"823d0d04",
X"fe3d0d02",
X"93053380",
X"e1f40853",
X"53807234",
X"8a51e5e8",
X"3fd33f80",
X"e2840852",
X"80f87234",
X"80e29c08",
X"52807234",
X"fa1380e2",
X"a4085353",
X"72723480",
X"e28c0852",
X"80723480",
X"e2940852",
X"72723480",
X"e1f80852",
X"80723480",
X"e1f80852",
X"b8723484",
X"3d0d04ff",
X"3d0d028f",
X"053380e1",
X"fc085252",
X"717134fe",
X"9e3f83e0",
X"8008802e",
X"f638833d",
X"0d04803d",
X"0d8439ee",
X"c83ffeb8",
X"3f83e080",
X"08802ef3",
X"3880e1fc",
X"08703370",
X"81ff0683",
X"e0800c51",
X"51823d0d",
X"04803d0d",
X"80e1f408",
X"51a37134",
X"80e28008",
X"51ff7134",
X"80e1f808",
X"51a87134",
X"80e1f808",
X"51b87134",
X"823d0d04",
X"803d0d80",
X"e1f40870",
X"337081c0",
X"06703070",
X"802583e0",
X"800c5151",
X"5151823d",
X"0d04ff3d",
X"0d80e1f8",
X"08703370",
X"81ff0670",
X"832a8132",
X"70810651",
X"51515252",
X"70802ee5",
X"38b07234",
X"80e1f808",
X"51b87134",
X"833d0d04",
X"803d0d80",
X"e2b00870",
X"08810683",
X"e0800c51",
X"823d0d04",
X"fd3d0d75",
X"77545480",
X"73259438",
X"73708105",
X"55335280",
X"e0e85185",
X"9d3fff13",
X"53e93985",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"adba3f83",
X"e080087a",
X"27ee3874",
X"802e80dd",
X"38745275",
X"51ada53f",
X"83e08008",
X"75537652",
X"54adcc3f",
X"83e08008",
X"7a537552",
X"56ad8d3f",
X"83e08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"e08008c5",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9f",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fc813f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd53f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbb13f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83e0900c",
X"7183e094",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383e090",
X"085283e0",
X"940851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"adfe5351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fd3d",
X"0d757052",
X"54a5b63f",
X"83e08008",
X"14537274",
X"2e9238ff",
X"13703353",
X"5371af2e",
X"098106ee",
X"38811353",
X"7283e080",
X"0c853d0d",
X"04fd3d0d",
X"75777053",
X"5454c73f",
X"83e08008",
X"732ea138",
X"83e08008",
X"733152ff",
X"125271ff",
X"2e8f3872",
X"70810554",
X"33747081",
X"055634eb",
X"39ff1454",
X"80743485",
X"3d0d0480",
X"3d0d7251",
X"ff903f82",
X"3d0d0471",
X"83e0800c",
X"04803d0d",
X"72518071",
X"34810bbc",
X"120c800b",
X"80c0120c",
X"823d0d04",
X"800b83e2",
X"f808248a",
X"38a6a63f",
X"ff0b83e2",
X"f80c800b",
X"83e0800c",
X"04ff3d0d",
X"735283e0",
X"d408722e",
X"8d38d93f",
X"715197b7",
X"3f7183e0",
X"d40c833d",
X"0d04f43d",
X"0d7e6062",
X"5c5a5581",
X"54bc1508",
X"81913874",
X"51cf3f79",
X"58807a25",
X"80f73883",
X"e3a80870",
X"892a5783",
X"ff067884",
X"80723156",
X"56577378",
X"25833873",
X"557583e2",
X"f8082e84",
X"38ff893f",
X"83e2f808",
X"8025a638",
X"75892b51",
X"9aa33f83",
X"e3a8088f",
X"3dfc1155",
X"5c548152",
X"f81b5198",
X"883f7614",
X"83e3a80c",
X"7583e2f8",
X"0c745376",
X"527851a4",
X"b93f83e0",
X"800883e3",
X"a8081683",
X"e3a80c78",
X"7631761b",
X"5b595677",
X"8024ff8b",
X"38617a71",
X"0c547554",
X"75802e83",
X"38815473",
X"83e0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"9b3f7651",
X"feaf3f86",
X"3dfc0553",
X"02a20522",
X"52775197",
X"a83f7986",
X"3d22710c",
X"5483e080",
X"085483e0",
X"8008802e",
X"83388154",
X"7383e080",
X"0c863d0d",
X"04fd3d0d",
X"7683e2f8",
X"08535380",
X"72248938",
X"71732e84",
X"38fdd13f",
X"7551fde5",
X"3f725198",
X"f03f7352",
X"73802e83",
X"38815271",
X"83e0800c",
X"853d0d04",
X"803d0d72",
X"80c01108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"72bc1108",
X"83e0800c",
X"51823d0d",
X"0480c40b",
X"83e0800c",
X"04fd3d0d",
X"75777154",
X"70535553",
X"a18f3f82",
X"c81308bc",
X"150c82c0",
X"130880c0",
X"150cfcec",
X"3f735194",
X"ca3f7383",
X"e0d40c83",
X"e0800853",
X"83e08008",
X"802e8338",
X"81537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"5553fcc0",
X"3f72802e",
X"a538bc13",
X"08527351",
X"a0993f83",
X"e080088f",
X"38775272",
X"51ff9a3f",
X"83e08008",
X"538a3982",
X"cc130853",
X"d8398153",
X"7283e080",
X"0c853d0d",
X"04fe3d0d",
X"ff0b83e2",
X"f80c7483",
X"e0d80c75",
X"83e2f40c",
X"a0fe3f83",
X"e0800881",
X"ff065281",
X"53719938",
X"83e39051",
X"8fc23f83",
X"e0800852",
X"83e08008",
X"802e8338",
X"72527153",
X"7283e080",
X"0c843d0d",
X"04fa3d0d",
X"787a82c4",
X"120882c4",
X"12087072",
X"24595656",
X"57577373",
X"2e098106",
X"913880c0",
X"165280c0",
X"17519e8a",
X"3f83e080",
X"08557483",
X"e0800c88",
X"3d0d04f6",
X"3d0d7c5b",
X"807b715c",
X"54577a77",
X"2e8c3881",
X"1a82cc14",
X"08545a72",
X"f6388059",
X"80d9397a",
X"54815780",
X"707b7b31",
X"5a5755ff",
X"18537473",
X"2580c138",
X"82cc1408",
X"527351ff",
X"8c3f800b",
X"83e08008",
X"25a13882",
X"cc140882",
X"cc110882",
X"cc160c74",
X"82cc120c",
X"5375802e",
X"86387282",
X"cc170c72",
X"54805773",
X"82cc1508",
X"81175755",
X"56ffb839",
X"81195980",
X"0bff1b54",
X"54787325",
X"83388154",
X"76813270",
X"75065153",
X"72ff9038",
X"8c3d0d04",
X"f53d0d7d",
X"7f5c5c82",
X"d05283e2",
X"f40851a0",
X"c73f83e0",
X"800859f9",
X"e33f80e0",
X"f051f7f6",
X"3f7b5283",
X"e2fc5196",
X"f23f83e0",
X"80085580",
X"5683e080",
X"08762e09",
X"810682ae",
X"3880e0fc",
X"51f7d33f",
X"83e0d808",
X"80e0a053",
X"7052579d",
X"bc3f80e0",
X"a05280c0",
X"17519db1",
X"3f76bc18",
X"0c7482c0",
X"180c810b",
X"82c4180c",
X"810b82c8",
X"180cff19",
X"75595981",
X"b83983e0",
X"e4337082",
X"2a708106",
X"51565674",
X"81a73875",
X"812a8106",
X"5a79819d",
X"3878802e",
X"81b13882",
X"d017ff1a",
X"77842a81",
X"0682c413",
X"0c83e0e4",
X"33810682",
X"c8130c83",
X"e0e55480",
X"e180535a",
X"58f6d73f",
X"7b527751",
X"9cc73f77",
X"519cde3f",
X"83e08008",
X"1855af75",
X"70810557",
X"3474bc19",
X"0c83e0e5",
X"5274519c",
X"a83f83e0",
X"dc0882c0",
X"190c83e0",
X"f2528390",
X"17519c95",
X"3f7982cc",
X"190c7a80",
X"2e8d3877",
X"517a2d83",
X"e0800880",
X"2ea33876",
X"802e8638",
X"7782cc18",
X"0c7782cc",
X"19085582",
X"c0190854",
X"83e0dc08",
X"5380e184",
X"5257f5e6",
X"3f83e0dc",
X"5283e2fc",
X"5195ee3f",
X"83e08008",
X"8a3883e0",
X"e5335574",
X"feb03880",
X"e19051f5",
X"c53f800b",
X"82cc190c",
X"7a802e89",
X"3883e0d8",
X"0851fc87",
X"3f83e0d8",
X"08567583",
X"e0800c8d",
X"3d0d04ff",
X"3d0d8052",
X"7351fd84",
X"3f833d0d",
X"04f03d0d",
X"62705254",
X"f5e03f83",
X"e0800874",
X"53873d70",
X"535555f6",
X"803ff6e0",
X"3f7351d3",
X"3f635374",
X"5283e080",
X"0851fa87",
X"3f923d0d",
X"047183e0",
X"800c0480",
X"c01283e0",
X"800c0480",
X"3d0d7282",
X"c0110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"82cc1108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"7282c411",
X"0883e080",
X"0c51823d",
X"0d04f63d",
X"0d7c83e0",
X"98085959",
X"81792782",
X"a9387888",
X"19082782",
X"a1387733",
X"5675822e",
X"819b3875",
X"82248938",
X"75812e8d",
X"38828b39",
X"75832e81",
X"b7388282",
X"397883ff",
X"ff067081",
X"2a117083",
X"ffff0670",
X"83ff0671",
X"892a903d",
X"5f525a51",
X"51557683",
X"ff2e8e38",
X"82547653",
X"8c180815",
X"527951a9",
X"39755476",
X"538c1808",
X"15527951",
X"9ab33f83",
X"e0800881",
X"bd387554",
X"83e08008",
X"538c1808",
X"15810552",
X"8c3dfd05",
X"519a963f",
X"83e08008",
X"81a03802",
X"a905338c",
X"3d337188",
X"2b077a81",
X"0671842a",
X"53575856",
X"74863876",
X"9fff0656",
X"75558180",
X"39755478",
X"1083fe06",
X"5378882a",
X"8c190805",
X"528c3dfc",
X"055199d5",
X"3f83e080",
X"0880df38",
X"02a90533",
X"8c3d3371",
X"882b0756",
X"5780d139",
X"84547882",
X"2b83fc06",
X"5378872a",
X"8c190805",
X"528c3dfc",
X"055199a5",
X"3f83e080",
X"08b03802",
X"ab053302",
X"8405aa05",
X"3371982b",
X"71902b07",
X"028c05a9",
X"05337088",
X"2b720790",
X"3d337180",
X"fffffe80",
X"06075152",
X"53575856",
X"83398155",
X"7483e080",
X"0c8c3d0d",
X"04fb3d0d",
X"83e09808",
X"fe198812",
X"08fe0555",
X"56548056",
X"7473278d",
X"38821433",
X"75712994",
X"16080557",
X"537583e0",
X"800c873d",
X"0d04fc3d",
X"0d7683e0",
X"98085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"ff933f83",
X"e0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183e080",
X"0c863d0d",
X"04fa3d0d",
X"7883e098",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fbdb3f",
X"81527183",
X"e0800827",
X"a8388352",
X"83e08008",
X"88170827",
X"9c3883e0",
X"80088c16",
X"0c83e080",
X"0851fdf9",
X"3f83e080",
X"0890160c",
X"73752380",
X"527183e0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585d5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"a0269138",
X"7a51fdd2",
X"3f83e080",
X"0856807c",
X"3483a839",
X"933d841c",
X"0870585a",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"38807059",
X"5d887f08",
X"5f5a7c81",
X"1e7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535f57",
X"557480d8",
X"3876ae2e",
X"09810683",
X"38815577",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675ac",
X"3888588b",
X"5affab39",
X"ff9f1755",
X"74992689",
X"38e01770",
X"81ff0658",
X"55778119",
X"7081ff06",
X"721c535a",
X"57557675",
X"34ff8739",
X"7c1e7f0c",
X"805576a0",
X"26833881",
X"55748b1a",
X"347a51fc",
X"913f83e0",
X"800880f5",
X"38a0547a",
X"2270852b",
X"83e00654",
X"55901b08",
X"527b5194",
X"ac3f83e0",
X"80085783",
X"e0800881",
X"82387b33",
X"5574802e",
X"80f5388b",
X"1c337083",
X"2a708106",
X"51565674",
X"b4388b7c",
X"841d0883",
X"e0800859",
X"5b5b58ff",
X"185877ff",
X"2e9a3879",
X"7081055b",
X"33797081",
X"055b3371",
X"71315256",
X"5675802e",
X"e2388639",
X"75802ebc",
X"387a51fb",
X"f43fff86",
X"3983e080",
X"085683e0",
X"8008802e",
X"a93883e0",
X"8008832e",
X"09810680",
X"de38841b",
X"088b1133",
X"51557480",
X"d2388456",
X"80cd3983",
X"56ec3981",
X"5680c439",
X"7656841b",
X"088b1133",
X"515574b7",
X"388b1c33",
X"70842a70",
X"81065156",
X"5774802e",
X"d538951c",
X"33941d33",
X"71982b71",
X"902b079b",
X"1f337f9a",
X"05337188",
X"2b077207",
X"7f88050c",
X"5a585658",
X"fcda3975",
X"83e0800c",
X"903d0d04",
X"f83d0d7a",
X"7c595782",
X"5483fe53",
X"77527651",
X"92bb3f83",
X"5683e080",
X"0880ec38",
X"81173377",
X"3371882b",
X"07565682",
X"567482d4",
X"d52e0981",
X"0680d438",
X"7554b653",
X"77527651",
X"928f3f83",
X"e0800898",
X"38811733",
X"77337188",
X"2b0783e0",
X"80085256",
X"56748182",
X"c62eac38",
X"825480d2",
X"53775276",
X"5191e63f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62e83",
X"38815675",
X"83e0800c",
X"8a3d0d04",
X"ec3d0d66",
X"59800b83",
X"e0980c78",
X"5678802e",
X"83e83891",
X"933f83e0",
X"80088106",
X"55825674",
X"83d83874",
X"75538e3d",
X"70535858",
X"fec23f83",
X"e0800881",
X"ff065675",
X"812e0981",
X"0680d438",
X"905483be",
X"53745276",
X"5190f23f",
X"83e08008",
X"80c9388e",
X"3d335574",
X"802e80c9",
X"3802bb05",
X"33028405",
X"ba053371",
X"982b7190",
X"2b07028c",
X"05b90533",
X"70882b72",
X"07943d33",
X"71077058",
X"7c575452",
X"5d575956",
X"fde63f83",
X"e0800881",
X"ff065675",
X"832e0981",
X"06863881",
X"5682db39",
X"75802e86",
X"38875682",
X"d139a454",
X"8d537752",
X"76519089",
X"3f815683",
X"e0800882",
X"bd3802ba",
X"05330284",
X"05b90533",
X"71882b07",
X"585c76ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"0754525d",
X"57585602",
X"b3053377",
X"71290288",
X"05b20533",
X"028c05b1",
X"05337188",
X"2b07701c",
X"708c1f0c",
X"5e595758",
X"5c8d3d33",
X"821a3402",
X"b505338f",
X"3d337188",
X"2b07595b",
X"77841a23",
X"02b70533",
X"028405b6",
X"05337188",
X"2b07565b",
X"74ab3802",
X"80c60533",
X"02840580",
X"c5053371",
X"982b7190",
X"2b07953d",
X"3370882b",
X"72070294",
X"0580c305",
X"33710751",
X"5253575d",
X"5b747631",
X"77317884",
X"2a8f3d33",
X"54717131",
X"5356568f",
X"f73f83e0",
X"80088205",
X"70881b0c",
X"709ff626",
X"81055755",
X"83fff675",
X"27833883",
X"56757934",
X"75832e09",
X"8106af38",
X"0280d205",
X"33028405",
X"80d10533",
X"71982b71",
X"902b0798",
X"3d337088",
X"2b720702",
X"940580cf",
X"05337107",
X"901f0c52",
X"5d575956",
X"8639761a",
X"901a0c84",
X"19228c1a",
X"08187184",
X"2a05941b",
X"0c5c800b",
X"811a3478",
X"83e0980c",
X"80567583",
X"e0800c96",
X"3d0d04e9",
X"3d0d83e0",
X"98085686",
X"5475802e",
X"81a63880",
X"0b811734",
X"993de011",
X"466a54c0",
X"1153ec05",
X"51f6cf3f",
X"83e08008",
X"5483e080",
X"08818538",
X"893d3354",
X"73802e93",
X"3802ab05",
X"3370842a",
X"70810651",
X"55557380",
X"2e863883",
X"5480e539",
X"02b50533",
X"8f3d3371",
X"982b7190",
X"2b07028c",
X"05bb0533",
X"029005ba",
X"05337188",
X"2b077207",
X"a01b0c02",
X"9005bf05",
X"33029405",
X"be053371",
X"982b7190",
X"2b07029c",
X"05bd0533",
X"70882b72",
X"07993d33",
X"71077f9c",
X"050c5283",
X"e0800898",
X"1f0c565a",
X"52525357",
X"5957810b",
X"81173483",
X"e0800854",
X"7383e080",
X"0c993d0d",
X"04f53d0d",
X"7d600288",
X"05ba0522",
X"7283e098",
X"085b5d5a",
X"5c5c807b",
X"23865676",
X"802e81e0",
X"38811733",
X"81065585",
X"5674802e",
X"81d2389c",
X"17089818",
X"08315574",
X"78278738",
X"7483ffff",
X"06587780",
X"2e81ae38",
X"98170870",
X"83ff0656",
X"567480ca",
X"38821733",
X"ff057689",
X"2a067081",
X"ff065a55",
X"78a03875",
X"8738a017",
X"08558d39",
X"a4170851",
X"efe03f83",
X"e0800855",
X"81752780",
X"f83874a4",
X"180ca417",
X"0851f28d",
X"3f83e080",
X"08802e80",
X"e43883e0",
X"800819a8",
X"180c9817",
X"0883ff06",
X"84807131",
X"7083ffff",
X"06585155",
X"77762783",
X"38775675",
X"54981708",
X"83ff0653",
X"a8170852",
X"79557b83",
X"387b5574",
X"518aae3f",
X"83e08008",
X"a4389817",
X"08169818",
X"0c751a78",
X"77317083",
X"ffff067d",
X"22790552",
X"5a565a74",
X"7b23fece",
X"39805688",
X"39800b81",
X"18348156",
X"7583e080",
X"0c8d3d0d",
X"04fa3d0d",
X"7883e098",
X"08555686",
X"5573802e",
X"81dc3881",
X"14338106",
X"53855572",
X"802e81ce",
X"389c1408",
X"53727627",
X"83387256",
X"98140857",
X"800b9815",
X"0c75802e",
X"81a93882",
X"14337089",
X"2b565376",
X"802eb538",
X"7452ff16",
X"518ae53f",
X"83e08008",
X"ff187654",
X"70535853",
X"8ad63f83",
X"e0800873",
X"26963874",
X"30707806",
X"7098170c",
X"777131a4",
X"17085258",
X"51538939",
X"a0140870",
X"a4160c53",
X"747627b4",
X"387251ed",
X"c13f83e0",
X"80085381",
X"0b83e080",
X"082780cb",
X"3883e080",
X"08881508",
X"2780c038",
X"83e08008",
X"a4150c98",
X"14081598",
X"150c7575",
X"3156c939",
X"98140816",
X"7098160c",
X"735256ef",
X"c83f83e0",
X"8008802e",
X"96388214",
X"33ff0576",
X"892a0683",
X"e0800805",
X"a8150c80",
X"55883980",
X"0b811534",
X"81557483",
X"e0800c88",
X"3d0d04ee",
X"3d0d6456",
X"865583e0",
X"9808802e",
X"80f63894",
X"3df41184",
X"180c6654",
X"d4055275",
X"51f1973f",
X"83e08008",
X"5583e080",
X"0880cf38",
X"893d3354",
X"73802ebc",
X"3802ab05",
X"3370842a",
X"70810651",
X"55558455",
X"73802ebc",
X"3802b505",
X"338f3d33",
X"71982b71",
X"902b0702",
X"8c05bb05",
X"33029005",
X"ba053371",
X"882b0772",
X"07881b0c",
X"53575957",
X"7551eed2",
X"3f83e080",
X"08557483",
X"2e098106",
X"83388455",
X"7483e080",
X"0c943d0d",
X"04e43d0d",
X"6ea13d08",
X"405d8656",
X"83e09808",
X"802e8491",
X"389e3df4",
X"05841e0c",
X"7e98387c",
X"51ee973f",
X"83e08008",
X"5683fa39",
X"814181f6",
X"39834181",
X"f139933d",
X"7f960541",
X"59807f82",
X"95055f56",
X"756081ff",
X"05348341",
X"901d0876",
X"2e81d338",
X"a0547c22",
X"70852b83",
X"e0065458",
X"901d0852",
X"78518689",
X"3f83e080",
X"084183e0",
X"8008ffb8",
X"3878335c",
X"7b802eff",
X"b4388b19",
X"3370bf06",
X"71810652",
X"43557480",
X"2e80de38",
X"7b81bf06",
X"55748f24",
X"80d3389a",
X"19335574",
X"80cb38f3",
X"1e70585e",
X"8156758b",
X"2e098106",
X"85388e56",
X"8b39759a",
X"2e098106",
X"83389c56",
X"75197070",
X"81055233",
X"7133811a",
X"821a5f5b",
X"525b5574",
X"86387977",
X"34853980",
X"df773477",
X"7b57577a",
X"a02e0981",
X"06c03881",
X"567b81e5",
X"32703070",
X"9f2a5151",
X"557bae2e",
X"93387480",
X"2e8e3861",
X"832a7081",
X"06515574",
X"802e9738",
X"7c51ed81",
X"3f83e080",
X"084183e0",
X"80088738",
X"901d08fe",
X"af388060",
X"3475802e",
X"88387d52",
X"7f5183b1",
X"3f60802e",
X"8638800b",
X"901e0c60",
X"5660832e",
X"09810688",
X"38800b90",
X"1e0c8539",
X"6081d238",
X"891f5790",
X"1d08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347c51eb",
X"883f83e0",
X"80085683",
X"e0800883",
X"2e098106",
X"8838800b",
X"901e0c80",
X"56961f33",
X"55748a38",
X"891f5296",
X"1f5181b1",
X"3f7583e0",
X"800c9e3d",
X"0d04fd3d",
X"0d757753",
X"54733351",
X"70893871",
X"33517080",
X"2ea13873",
X"33723352",
X"53727127",
X"8538ff51",
X"94397073",
X"27853881",
X"518b3981",
X"14811353",
X"54d33980",
X"517083e0",
X"800c853d",
X"0d04fd3d",
X"0d757754",
X"54723370",
X"81ff0652",
X"5270802e",
X"a3387181",
X"ff068114",
X"ffbf1253",
X"54527099",
X"268938a0",
X"127081ff",
X"06535171",
X"74708105",
X"5634d239",
X"80743485",
X"3d0d04ff",
X"bd3d0d80",
X"c63d0852",
X"a53d7052",
X"54ffb33f",
X"80c73d08",
X"52853d70",
X"5253ffa6",
X"3f725273",
X"51fedf3f",
X"80c53d0d",
X"04fe3d0d",
X"74765353",
X"71708105",
X"53335170",
X"73708105",
X"553470f0",
X"38843d0d",
X"04fe3d0d",
X"74528072",
X"33525370",
X"732e8d38",
X"81128114",
X"71335354",
X"5270f538",
X"7283e080",
X"0c843d0d",
X"04fd3d0d",
X"75547383",
X"e3c0082e",
X"a73880e2",
X"c00874a0",
X"0a07710c",
X"80e2d008",
X"53537108",
X"5170802e",
X"f9388073",
X"0c710851",
X"70fb3873",
X"83e3c00c",
X"853d0d04",
X"ff0b83e3",
X"c00c8180",
X"800b83e3",
X"bc0c800b",
X"83e0800c",
X"04fc3d0d",
X"76028405",
X"a2052202",
X"8805a605",
X"227a5455",
X"5555ff9d",
X"3f72802e",
X"a33883e3",
X"bc081452",
X"71337570",
X"81055734",
X"81147083",
X"ffff06ff",
X"157083ff",
X"ff065652",
X"5552da39",
X"800b83e0",
X"800c863d",
X"0d04f73d",
X"0d7b7d7f",
X"11585559",
X"80557376",
X"2eb13883",
X"e3bc088b",
X"3d595774",
X"19703375",
X"fc061970",
X"085d7683",
X"067b0753",
X"54545172",
X"71347972",
X"0c811481",
X"16565473",
X"762e0981",
X"06d93880",
X"0b83e080",
X"0c8b3d0d",
X"04fe3d0d",
X"80e2c008",
X"83e3c008",
X"900a0771",
X"0c80e2d0",
X"08535371",
X"08517080",
X"2ef93880",
X"730c7108",
X"5170fb38",
X"843d0d04",
X"83e08c08",
X"0283e08c",
X"0cfd3d0d",
X"805383e0",
X"8c088c05",
X"085283e0",
X"8c088805",
X"085183d4",
X"3f83e080",
X"087083e0",
X"800c5485",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"fd3d0d81",
X"5383e08c",
X"088c0508",
X"5283e08c",
X"08880508",
X"5183a13f",
X"83e08008",
X"7083e080",
X"0c54853d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cf9",
X"3d0d800b",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"05088025",
X"b93883e0",
X"8c088805",
X"083083e0",
X"8c088805",
X"0c800b83",
X"e08c08f4",
X"050c83e0",
X"8c08fc05",
X"088a3881",
X"0b83e08c",
X"08f4050c",
X"83e08c08",
X"f4050883",
X"e08c08fc",
X"050c83e0",
X"8c088c05",
X"088025b9",
X"3883e08c",
X"088c0508",
X"3083e08c",
X"088c050c",
X"800b83e0",
X"8c08f005",
X"0c83e08c",
X"08fc0508",
X"8a38810b",
X"83e08c08",
X"f0050c83",
X"e08c08f0",
X"050883e0",
X"8c08fc05",
X"0c805383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"05085181",
X"df3f83e0",
X"80087083",
X"e08c08f8",
X"050c5483",
X"e08c08fc",
X"0508802e",
X"903883e0",
X"8c08f805",
X"083083e0",
X"8c08f805",
X"0c83e08c",
X"08f80508",
X"7083e080",
X"0c54893d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cfb",
X"3d0d800b",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"05088025",
X"993883e0",
X"8c088805",
X"083083e0",
X"8c088805",
X"0c810b83",
X"e08c08fc",
X"050c83e0",
X"8c088c05",
X"08802590",
X"3883e08c",
X"088c0508",
X"3083e08c",
X"088c050c",
X"815383e0",
X"8c088c05",
X"085283e0",
X"8c088805",
X"0851bd3f",
X"83e08008",
X"7083e08c",
X"08f8050c",
X"5483e08c",
X"08fc0508",
X"802e9038",
X"83e08c08",
X"f8050830",
X"83e08c08",
X"f8050c83",
X"e08c08f8",
X"05087083",
X"e0800c54",
X"873d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cfd3d0d",
X"810b83e0",
X"8c08fc05",
X"0c800b83",
X"e08c08f8",
X"050c83e0",
X"8c088c05",
X"0883e08c",
X"08880508",
X"27b93883",
X"e08c08fc",
X"0508802e",
X"ae38800b",
X"83e08c08",
X"8c050824",
X"a23883e0",
X"8c088c05",
X"081083e0",
X"8c088c05",
X"0c83e08c",
X"08fc0508",
X"1083e08c",
X"08fc050c",
X"ffb83983",
X"e08c08fc",
X"0508802e",
X"80e13883",
X"e08c088c",
X"050883e0",
X"8c088805",
X"0826ad38",
X"83e08c08",
X"88050883",
X"e08c088c",
X"05083183",
X"e08c0888",
X"050c83e0",
X"8c08f805",
X"0883e08c",
X"08fc0508",
X"0783e08c",
X"08f8050c",
X"83e08c08",
X"fc050881",
X"2a83e08c",
X"08fc050c",
X"83e08c08",
X"8c050881",
X"2a83e08c",
X"088c050c",
X"ff953983",
X"e08c0890",
X"0508802e",
X"933883e0",
X"8c088805",
X"087083e0",
X"8c08f405",
X"0c519139",
X"83e08c08",
X"f8050870",
X"83e08c08",
X"f4050c51",
X"83e08c08",
X"f4050883",
X"e0800c85",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"ff3d0d80",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"88050881",
X"06ff1170",
X"097083e0",
X"8c088c05",
X"080683e0",
X"8c08fc05",
X"081183e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"812a83e0",
X"8c088805",
X"0c83e08c",
X"088c0508",
X"1083e08c",
X"088c050c",
X"51515151",
X"83e08c08",
X"88050880",
X"2e8438ff",
X"ab3983e0",
X"8c08fc05",
X"087083e0",
X"800c5183",
X"3d0d83e0",
X"8c0c04fc",
X"3d0d7670",
X"797b5555",
X"55558f72",
X"278c3872",
X"75078306",
X"5170802e",
X"a938ff12",
X"5271ff2e",
X"98387270",
X"81055433",
X"74708105",
X"5634ff12",
X"5271ff2e",
X"098106ea",
X"387483e0",
X"800c863d",
X"0d047451",
X"72708405",
X"54087170",
X"8405530c",
X"72708405",
X"54087170",
X"8405530c",
X"72708405",
X"54087170",
X"8405530c",
X"72708405",
X"54087170",
X"8405530c",
X"f0125271",
X"8f26c938",
X"83722795",
X"38727084",
X"05540871",
X"70840553",
X"0cfc1252",
X"718326ed",
X"387054ff",
X"81390000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"0000097b",
X"000009bc",
X"000009dd",
X"000009fb",
X"000009fb",
X"000009fb",
X"00000ab5",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"31364b00",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"43617274",
X"72696467",
X"65203332",
X"6b000000",
X"43617274",
X"72696467",
X"65203136",
X"6b206f6e",
X"65206368",
X"69700000",
X"43617274",
X"72696467",
X"65203136",
X"6b207477",
X"6f206368",
X"69700000",
X"45786974",
X"00000000",
X"61636964",
X"35323030",
X"2e726f6d",
X"00000000",
X"25732025",
X"73000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"66696c74",
X"65725f64",
X"69736b73",
X"3a25733a",
X"25640a00",
X"524f4d00",
X"42494e00",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"6f70656e",
X"64697220",
X"00000000",
X"4f4b2000",
X"25732000",
X"6e202564",
X"20256420",
X"25782000",
X"6469725f",
X"656e7472",
X"69657320",
X"646f6e65",
X"20000000",
X"00000000",
X"00000000",
X"0001e80a",
X"0001e809",
X"0001e80f",
X"0001d40e",
X"0001d403",
X"0001d402",
X"0001d400",
X"0001d401",
X"0001d409",
X"0001d301",
X"0001d300",
X"0001c010",
X"0001c01b",
X"0001c016",
X"0001c019",
X"0001c018",
X"0001c017",
X"0001c01a",
X"0004007c",
X"00040078",
X"00040074",
X"00040068",
X"00040060",
X"0004005c",
X"00040058",
X"00040054",
X"00040050",
X"0004004c",
X"00040048",
X"00040044",
X"00040040",
X"00040034",
X"00040030",
X"0004002c",
X"00040028",
X"00040024",
X"00040020",
X"0004001c",
X"00040018",
X"00040014",
X"00040010",
X"0004000c",
X"00040008",
X"00040004",
X"00040000",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
