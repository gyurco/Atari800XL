
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80ef",
X"f4738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80f3",
X"ac0c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580eb",
X"bf2d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580e9d3",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80d1ae04",
X"f23d0d60",
X"913dec11",
X"56565990",
X"53f01552",
X"7851948a",
X"3f83e080",
X"0880e538",
X"7a902e09",
X"810680dc",
X"3802b305",
X"3380f3b4",
X"0b80f3b4",
X"33575757",
X"8c397477",
X"2e8a3884",
X"16703356",
X"5674f338",
X"75337058",
X"5574802e",
X"80cf3880",
X"0b821722",
X"70832a57",
X"58587775",
X"27bb3896",
X"800a5790",
X"3dec0554",
X"80c08053",
X"76527851",
X"93ac3f83",
X"e0800888",
X"387a80c0",
X"802e8538",
X"80579a39",
X"811880c0",
X"80188218",
X"2270832a",
X"585c5858",
X"747826cb",
X"38811633",
X"577683e0",
X"800c903d",
X"0d04fc3d",
X"0d767052",
X"55b3cc3f",
X"83e08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"811451b2",
X"e43f83e0",
X"80083070",
X"83e08008",
X"07802583",
X"e0800c53",
X"863d0d04",
X"fc3d0d76",
X"7052559a",
X"833f83e0",
X"80085481",
X"5383e080",
X"0880c738",
X"745199c6",
X"3f83e080",
X"080b0b80",
X"f1b45383",
X"e0800852",
X"53ff8f3f",
X"83e08008",
X"a5380b0b",
X"80f1b852",
X"7251fefe",
X"3f83e080",
X"0894380b",
X"0b80f1bc",
X"527251fe",
X"ed3f83e0",
X"8008802e",
X"83388154",
X"73537283",
X"e0800c86",
X"3d0d04fd",
X"3d0d7570",
X"5254999c",
X"3f815383",
X"e0800898",
X"38735198",
X"e53f83e0",
X"a0085283",
X"e0800851",
X"feb43f83",
X"e0800853",
X"7283e080",
X"0c853d0d",
X"04e03d0d",
X"a33d0870",
X"525e8f87",
X"3f83e080",
X"0833943d",
X"56547394",
X"3880f7e0",
X"52745184",
X"c6397d52",
X"7851928c",
X"3f84d039",
X"7d518eef",
X"3f83e080",
X"08527451",
X"8e9f3f83",
X"e0a80852",
X"933d7052",
X"5d94fd3f",
X"83e08008",
X"59800b83",
X"e0800855",
X"5b83e080",
X"087b2e94",
X"38811b74",
X"525b97ff",
X"3f83e080",
X"085483e0",
X"8008ee38",
X"805aff7a",
X"437a427a",
X"415f7909",
X"709f2c7b",
X"065b547a",
X"7a248438",
X"ff1b5af6",
X"1a700970",
X"9f2c7206",
X"7bff125a",
X"5a525555",
X"80752595",
X"38765197",
X"be3f83e0",
X"800876ff",
X"18585557",
X"738024ed",
X"38747f2e",
X"8638b99e",
X"3f745f78",
X"ff1b7058",
X"5d58807a",
X"25953877",
X"5197943f",
X"83e08008",
X"76ff1858",
X"55587380",
X"24ed3880",
X"0b83e3a8",
X"0c800b83",
X"e3c80c0b",
X"0b80f1c0",
X"518be33f",
X"81800b83",
X"e3c80c0b",
X"0b80f1c8",
X"518bd33f",
X"a80b83e3",
X"a80c7680",
X"2e80e838",
X"83e3a808",
X"77793270",
X"30707207",
X"80257087",
X"2b83e3c8",
X"0c515678",
X"53565696",
X"c73f83e0",
X"8008802e",
X"8a380b0b",
X"80f1d051",
X"8b983f76",
X"5196873f",
X"83e08008",
X"520b0b80",
X"f2dc518b",
X"853f7651",
X"968d3f83",
X"e0800883",
X"e3a80855",
X"57757425",
X"8638a816",
X"56f73975",
X"83e3a80c",
X"86f07624",
X"ff943887",
X"980b83e3",
X"a80c7780",
X"2eb73877",
X"5195c33f",
X"83e08008",
X"78525595",
X"e33f0b0b",
X"80f1d854",
X"83e08008",
X"8f388739",
X"807634fd",
X"96390b0b",
X"80f1d454",
X"74537352",
X"0b0b80f1",
X"a8518a9e",
X"3f80540b",
X"0b80f3a8",
X"518a933f",
X"81145473",
X"a82e0981",
X"06ed3886",
X"8da051b5",
X"9d3f8052",
X"903d7052",
X"5480d5f9",
X"3f835273",
X"5180d5f1",
X"3f61802e",
X"80ff387b",
X"5473ff2e",
X"96387880",
X"2e818038",
X"785194e3",
X"3f83e080",
X"08ff1555",
X"59e73978",
X"802e80eb",
X"38785194",
X"df3f83e0",
X"8008802e",
X"fc843878",
X"5194a73f",
X"83e08008",
X"520b0b80",
X"f1b051ac",
X"873f83e0",
X"8008a438",
X"7c51adbf",
X"3f83e080",
X"085574ff",
X"16565480",
X"7425fbef",
X"38741d70",
X"33555673",
X"af2efec8",
X"38e83978",
X"5193e53f",
X"83e08008",
X"527c51ac",
X"f63ffbcf",
X"397f8829",
X"6010057a",
X"0561055a",
X"fc8039a2",
X"3d0d04fe",
X"3d0d80f6",
X"e8087033",
X"7081ff06",
X"70842a81",
X"32810655",
X"51525371",
X"802e8c38",
X"a8733480",
X"f6e80851",
X"b8713471",
X"83e0800c",
X"843d0d04",
X"fe3d0d80",
X"f6e80870",
X"337081ff",
X"0670852a",
X"81328106",
X"55515253",
X"71802e8c",
X"38987334",
X"80f6e808",
X"51b87134",
X"7183e080",
X"0c843d0d",
X"04803d0d",
X"80f6e408",
X"51937134",
X"80f6f008",
X"51ff7134",
X"823d0d04",
X"fe3d0d02",
X"93053380",
X"f6e40853",
X"53807234",
X"8a51b2e6",
X"3fd33f80",
X"f6f40852",
X"80f87234",
X"80f78c08",
X"52807234",
X"fa1380f7",
X"94085353",
X"72723480",
X"f6fc0852",
X"80723480",
X"f7840852",
X"72723480",
X"f6e80852",
X"80723480",
X"f6e80852",
X"b8723484",
X"3d0d04ff",
X"3d0d028f",
X"053380f6",
X"ec085252",
X"717134fe",
X"9e3f83e0",
X"8008802e",
X"f638833d",
X"0d04803d",
X"0d8439bc",
X"933ffeb8",
X"3f83e080",
X"08802ef3",
X"3880f6ec",
X"08703370",
X"81ff0683",
X"e0800c51",
X"51823d0d",
X"04803d0d",
X"80f6e408",
X"51a37134",
X"80f6f008",
X"51ff7134",
X"80f6e808",
X"51a87134",
X"80f6e808",
X"51b87134",
X"823d0d04",
X"803d0d80",
X"f6e40870",
X"337081c0",
X"06703070",
X"802583e0",
X"800c5151",
X"5151823d",
X"0d04ff3d",
X"0d80f6e8",
X"08703370",
X"81ff0670",
X"832a8132",
X"70810651",
X"51515252",
X"70802ee5",
X"38b07234",
X"80f6e808",
X"51b87134",
X"833d0d04",
X"803d0d80",
X"f7a00870",
X"08810683",
X"e0800c51",
X"823d0d04",
X"fd3d0d75",
X"77545480",
X"73259438",
X"73708105",
X"55335280",
X"f1dc5185",
X"a13fff13",
X"53e93985",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"80d3de3f",
X"83e08008",
X"7a27ed38",
X"74802e80",
X"e0387452",
X"755180d3",
X"c83f83e0",
X"80087553",
X"76525480",
X"d3ee3f83",
X"e080087a",
X"53755256",
X"80d3ae3f",
X"83e08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"e08008c2",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9c",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fbfd3f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd13f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbad3f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83e0900c",
X"7183e094",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383e090",
X"085283e0",
X"940851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"9aaa5351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fd3d",
X"0d757052",
X"54a3c83f",
X"83e08008",
X"14537274",
X"2e9238ff",
X"13703353",
X"5371af2e",
X"098106ee",
X"38811353",
X"7283e080",
X"0c853d0d",
X"04fd3d0d",
X"75777053",
X"5454c73f",
X"83e08008",
X"732ea138",
X"83e08008",
X"733152ff",
X"125271ff",
X"2e8f3872",
X"70810554",
X"33747081",
X"055634eb",
X"39ff1454",
X"80743485",
X"3d0d0480",
X"3d0d7251",
X"ff903f82",
X"3d0d0471",
X"83e0800c",
X"04803d0d",
X"72518071",
X"34810bbc",
X"120c800b",
X"80c0120c",
X"823d0d04",
X"800b83e2",
X"d408248b",
X"3880ccc6",
X"3fff0b83",
X"e2d40c80",
X"0b83e080",
X"0c04ff3d",
X"0d735283",
X"e0b00872",
X"2e8d38d8",
X"3f715196",
X"9c3f7183",
X"e0b00c83",
X"3d0d04f4",
X"3d0d7e60",
X"625c5a55",
X"8154bc15",
X"08819238",
X"7451cf3f",
X"7958807a",
X"2580f838",
X"83e38408",
X"70892a57",
X"83ff0678",
X"84807231",
X"56565773",
X"78258338",
X"73557583",
X"e2d4082e",
X"8438ff88",
X"3f83e2d4",
X"088025a6",
X"3875892b",
X"5198df3f",
X"83e38408",
X"8f3dfc11",
X"555c5481",
X"52f81b51",
X"96c93f76",
X"1483e384",
X"0c7583e2",
X"d40c7453",
X"76527851",
X"80cad83f",
X"83e08008",
X"83e38408",
X"1683e384",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8a3861",
X"7a710c54",
X"75547580",
X"2e833881",
X"547383e0",
X"800c8e3d",
X"0d04fc3d",
X"0dfe993f",
X"7651feae",
X"3f863dfc",
X"05537852",
X"775195eb",
X"3f797571",
X"0c5483e0",
X"80085483",
X"e0800880",
X"2e833881",
X"547383e0",
X"800c863d",
X"0d04fe3d",
X"0d7583e2",
X"d4085353",
X"80722489",
X"3871732e",
X"8438fdd4",
X"3f7451fd",
X"e93f7251",
X"97b03f83",
X"e0800852",
X"83e08008",
X"802e8338",
X"81527183",
X"e0800c84",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"e0800c51",
X"823d0d04",
X"80c40b83",
X"e0800c04",
X"fd3d0d75",
X"77715470",
X"5355539f",
X"9e3f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfce93f",
X"735193ad",
X"3f7383e0",
X"b00c83e0",
X"80085383",
X"e0800880",
X"2e833881",
X"537283e0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcbd3f",
X"72802ea5",
X"38bc1308",
X"5273519e",
X"a83f83e0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"e0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83e0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83e2d4",
X"0c7483e0",
X"b40c7583",
X"e2d00c80",
X"c79b3f83",
X"e0800881",
X"ff065281",
X"53719938",
X"83e2ec51",
X"8e963f83",
X"e0800852",
X"83e08008",
X"802e8338",
X"72527153",
X"7283e080",
X"0c843d0d",
X"04fa3d0d",
X"787a82c4",
X"120882c4",
X"12087072",
X"24595656",
X"57577373",
X"2e098106",
X"913880c0",
X"165280c0",
X"17519c98",
X"3f83e080",
X"08557483",
X"e0800c88",
X"3d0d04f6",
X"3d0d7c5b",
X"807b715c",
X"54577a77",
X"2e8c3881",
X"1a82cc14",
X"08545a72",
X"f6388059",
X"80d9397a",
X"54815780",
X"707b7b31",
X"5a5755ff",
X"18537473",
X"2580c138",
X"82cc1408",
X"527351ff",
X"8c3f800b",
X"83e08008",
X"25a13882",
X"cc140882",
X"cc110882",
X"cc160c74",
X"82cc120c",
X"5375802e",
X"86387282",
X"cc170c72",
X"54805773",
X"82cc1508",
X"81175755",
X"56ffb839",
X"81195980",
X"0bff1b54",
X"54787325",
X"83388154",
X"76813270",
X"75065153",
X"72ff9038",
X"8c3d0d04",
X"f73d0d7b",
X"7d5a5a82",
X"d05283e2",
X"d0085180",
X"c6e33f83",
X"e0800857",
X"f9de3f79",
X"5283e2d8",
X"5195b63f",
X"83e08008",
X"54805383",
X"e0800873",
X"2e098106",
X"82833883",
X"e0b4080b",
X"0b80f1b0",
X"53705256",
X"9bd53f0b",
X"0b80f1b0",
X"5280c016",
X"519bc83f",
X"75bc170c",
X"7382c017",
X"0c810b82",
X"c4170c81",
X"0b82c817",
X"0c7382cc",
X"170cff17",
X"82d01755",
X"57819139",
X"83e0c033",
X"70822a70",
X"81065154",
X"55728180",
X"3874812a",
X"81065877",
X"80f63874",
X"842a8106",
X"82c4150c",
X"83e0c033",
X"810682c8",
X"150c7952",
X"73519aef",
X"3f73519b",
X"863f83e0",
X"80081453",
X"af737081",
X"05553472",
X"bc150c83",
X"e0c15272",
X"519ad03f",
X"83e0b808",
X"82c0150c",
X"83e0ce52",
X"80c01451",
X"9abd3f78",
X"802e8d38",
X"7351782d",
X"83e08008",
X"802e9938",
X"7782cc15",
X"0c75802e",
X"86387382",
X"cc170c73",
X"82d015ff",
X"19595556",
X"76802e9b",
X"3883e0b8",
X"5283e2d8",
X"5194ac3f",
X"83e08008",
X"8a3883e0",
X"c1335372",
X"fed23878",
X"802e8938",
X"83e0b408",
X"51fcb83f",
X"83e0b408",
X"537283e0",
X"800c8b3d",
X"0d04ff3d",
X"0d805273",
X"51fdb53f",
X"833d0d04",
X"f03d0d62",
X"705254f6",
X"8d3f83e0",
X"80087453",
X"873d7053",
X"5555f6ad",
X"3ff78d3f",
X"7351d33f",
X"63537452",
X"83e08008",
X"51fab73f",
X"923d0d04",
X"7183e080",
X"0c0480c0",
X"1283e080",
X"0c04803d",
X"0d7282c0",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"cc110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"82c41108",
X"83e0800c",
X"51823d0d",
X"04f93d0d",
X"7983e098",
X"08575781",
X"77278198",
X"38768817",
X"08278190",
X"38753355",
X"74822e89",
X"3874832e",
X"b4388180",
X"39745476",
X"1083fe06",
X"5376882a",
X"8c170805",
X"52893dfc",
X"055180c1",
X"b53f83e0",
X"800880e0",
X"38029d05",
X"33893d33",
X"71882b07",
X"565680d2",
X"39845476",
X"822b83fc",
X"06537687",
X"2a8c1708",
X"0552893d",
X"fc055180",
X"c1843f83",
X"e08008b0",
X"38029f05",
X"33028405",
X"9e053371",
X"982b7190",
X"2b07028c",
X"059d0533",
X"70882b72",
X"078d3d33",
X"7180ffff",
X"fe800607",
X"51525357",
X"58568339",
X"81557483",
X"e0800c89",
X"3d0d04fb",
X"3d0d83e0",
X"9808fe19",
X"881208fe",
X"05555654",
X"80567473",
X"278d3882",
X"14337571",
X"29941608",
X"05575375",
X"83e0800c",
X"873d0d04",
X"fc3d0d76",
X"52800b83",
X"e0980870",
X"33515253",
X"70832e09",
X"81069138",
X"95123394",
X"13337198",
X"2b71902b",
X"07555551",
X"9b12339a",
X"13337188",
X"2b077407",
X"83e0800c",
X"55863d0d",
X"04fc3d0d",
X"7683e098",
X"08555580",
X"75238815",
X"08537281",
X"2e883888",
X"14087326",
X"85388152",
X"b2397290",
X"38733352",
X"71832e09",
X"81068538",
X"90140853",
X"728c160c",
X"72802e8d",
X"387251fe",
X"d63f83e0",
X"80085285",
X"39901408",
X"52719016",
X"0c805271",
X"83e0800c",
X"863d0d04",
X"fa3d0d78",
X"83e09808",
X"71228105",
X"7083ffff",
X"06575457",
X"5573802e",
X"88389015",
X"08537286",
X"38835280",
X"e739738f",
X"06527180",
X"da388113",
X"90160c8c",
X"15085372",
X"9038830b",
X"84172257",
X"52737627",
X"80c638bf",
X"39821633",
X"ff057484",
X"2a065271",
X"b2387251",
X"fcaf3f81",
X"527183e0",
X"800827a8",
X"38835283",
X"e0800888",
X"1708279c",
X"3883e080",
X"088c160c",
X"83e08008",
X"51fdbc3f",
X"83e08008",
X"90160c73",
X"75238052",
X"7183e080",
X"0c883d0d",
X"04f23d0d",
X"60626458",
X"5e5b7533",
X"5574a02e",
X"09810688",
X"38811670",
X"4456ef39",
X"62703356",
X"5674af2e",
X"09810684",
X"38811643",
X"800b881c",
X"0c627033",
X"5155749f",
X"2691387a",
X"51fdd23f",
X"83e08008",
X"56807d34",
X"83813993",
X"3d841c08",
X"7058595f",
X"8a55a076",
X"70810558",
X"34ff1555",
X"74ff2e09",
X"8106ef38",
X"80705a5c",
X"887f085f",
X"5a7b811d",
X"7081ff06",
X"60137033",
X"70af3270",
X"30a07327",
X"71802507",
X"5151525b",
X"535e5755",
X"7480e738",
X"76ae2e09",
X"81068338",
X"8155787a",
X"27750755",
X"74802e9f",
X"38798832",
X"703078ae",
X"32703070",
X"73079f2a",
X"53515751",
X"5675bb38",
X"88598b5a",
X"ffab3976",
X"982b5574",
X"80258738",
X"80ef8417",
X"3357ff9f",
X"17557499",
X"268938e0",
X"177081ff",
X"06585578",
X"811a7081",
X"ff06721b",
X"535b5755",
X"767534fe",
X"f8397b1e",
X"7f0c8055",
X"76a02683",
X"38815574",
X"8b19347a",
X"51fc823f",
X"83e08008",
X"80f538a0",
X"547a2270",
X"852b83e0",
X"06545590",
X"1b08527c",
X"51bbbf3f",
X"83e08008",
X"5783e080",
X"08818138",
X"7c335574",
X"802e80f4",
X"388b1d33",
X"70832a70",
X"81065156",
X"5674b438",
X"8b7d841d",
X"0883e080",
X"08595b5b",
X"58ff1858",
X"77ff2e9a",
X"38797081",
X"055b3379",
X"7081055b",
X"33717131",
X"52565675",
X"802ee238",
X"86397580",
X"2e96387a",
X"51fbe53f",
X"ff863983",
X"e0800856",
X"83e08008",
X"b6388339",
X"7656841b",
X"088b1133",
X"515574a7",
X"388b1d33",
X"70842a70",
X"81065156",
X"56748938",
X"83569439",
X"81569039",
X"7c51fa94",
X"3f83e080",
X"08881c0c",
X"fd813975",
X"83e0800c",
X"903d0d04",
X"f83d0d7a",
X"7c595782",
X"5483fe53",
X"77527651",
X"ba843f83",
X"5683e080",
X"0880ec38",
X"81173377",
X"3371882b",
X"07565682",
X"567482d4",
X"d52e0981",
X"0680d438",
X"7554b653",
X"77527651",
X"b9d83f83",
X"e0800898",
X"38811733",
X"77337188",
X"2b0783e0",
X"80085256",
X"56748182",
X"c62eac38",
X"825480d2",
X"53775276",
X"51b9af3f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62e83",
X"38815675",
X"83e0800c",
X"8a3d0d04",
X"eb3d0d67",
X"5a800b83",
X"e0980cb8",
X"e43f83e0",
X"80088106",
X"55825674",
X"83ee3874",
X"75538f3d",
X"70535759",
X"feca3f83",
X"e0800881",
X"ff065776",
X"812e0981",
X"0680d438",
X"905483be",
X"53745275",
X"51b8c33f",
X"83e08008",
X"80c9388f",
X"3d335574",
X"802e80c9",
X"3802bf05",
X"33028405",
X"be053371",
X"982b7190",
X"2b07028c",
X"05bd0533",
X"70882b72",
X"07953d33",
X"71077058",
X"7b575e52",
X"5e575957",
X"fdee3f83",
X"e0800881",
X"ff065776",
X"832e0981",
X"06863881",
X"5682f139",
X"76802e86",
X"38865682",
X"e739a454",
X"8d537852",
X"7551b7da",
X"3f815683",
X"e0800882",
X"d33802be",
X"05330284",
X"05bd0533",
X"71882b07",
X"595d77ab",
X"380280ce",
X"05330284",
X"0580cd05",
X"3371982b",
X"71902b07",
X"973d3370",
X"882b7207",
X"02940580",
X"cb053371",
X"0754525e",
X"57595602",
X"b7053378",
X"71290288",
X"05b60533",
X"028c05b5",
X"05337188",
X"2b07701d",
X"707f8c05",
X"0c5f5957",
X"595d8e3d",
X"33821b34",
X"02b90533",
X"903d3371",
X"882b075a",
X"5c78841b",
X"2302bb05",
X"33028405",
X"ba053371",
X"882b0756",
X"5c74ab38",
X"0280ca05",
X"33028405",
X"80c90533",
X"71982b71",
X"902b0796",
X"3d337088",
X"2b720702",
X"940580c7",
X"05337107",
X"51525357",
X"5e5c7476",
X"31783179",
X"842a903d",
X"33547171",
X"31535656",
X"b7c73f83",
X"e0800882",
X"0570881c",
X"0c83e080",
X"08e08a05",
X"56567483",
X"dffe2683",
X"38825783",
X"fff67627",
X"85388357",
X"89398656",
X"76802e80",
X"db38767a",
X"3476832e",
X"098106b0",
X"380280d6",
X"05330284",
X"0580d505",
X"3371982b",
X"71902b07",
X"993d3370",
X"882b7207",
X"02940580",
X"d3053371",
X"077f9005",
X"0c525e57",
X"58568639",
X"771b901b",
X"0c841a22",
X"8c1b0819",
X"71842a05",
X"941c0c5d",
X"800b811b",
X"347983e0",
X"980c8056",
X"7583e080",
X"0c973d0d",
X"04e93d0d",
X"83e09808",
X"56855475",
X"802e8182",
X"38800b81",
X"1734993d",
X"e011466a",
X"548a3d70",
X"5458ec05",
X"51f6e63f",
X"83e08008",
X"5483e080",
X"0880df38",
X"893d3354",
X"73802e91",
X"3802ab05",
X"3370842a",
X"81065155",
X"74802e86",
X"38835480",
X"c1397651",
X"f48a3f83",
X"e08008a0",
X"170c02bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"3371079c",
X"1c0c5278",
X"981b0c53",
X"56595781",
X"0b811734",
X"74547383",
X"e0800c99",
X"3d0d04f5",
X"3d0d7d7f",
X"617283e0",
X"98085a5d",
X"5d595c80",
X"7b0c8557",
X"75802e81",
X"e0388116",
X"33810655",
X"84577480",
X"2e81d238",
X"91397481",
X"17348639",
X"800b8117",
X"34815781",
X"c0399c16",
X"08981708",
X"31557478",
X"27833874",
X"5877802e",
X"81a93898",
X"16087083",
X"ff065657",
X"7480cf38",
X"821633ff",
X"0577892a",
X"067081ff",
X"065a5578",
X"a0387687",
X"38a01608",
X"558d39a4",
X"160851f0",
X"e83f83e0",
X"80085581",
X"7527ffa8",
X"3874a417",
X"0ca41608",
X"51f2843f",
X"83e08008",
X"5583e080",
X"08802eff",
X"893883e0",
X"800819a8",
X"170c9816",
X"0883ff06",
X"84807131",
X"51557775",
X"27833877",
X"557483ff",
X"ff065498",
X"160883ff",
X"0653a816",
X"08527957",
X"7b83387b",
X"577651b2",
X"813f83e0",
X"8008fed0",
X"38981608",
X"1598170c",
X"741a7876",
X"317c0817",
X"7d0c595a",
X"fed33980",
X"577683e0",
X"800c8d3d",
X"0d04fa3d",
X"0d7883e0",
X"98085556",
X"85557380",
X"2e81e138",
X"81143381",
X"06538455",
X"72802e81",
X"d3389c14",
X"08537276",
X"27833872",
X"56981408",
X"57800b98",
X"150c7580",
X"2e81b738",
X"82143370",
X"892b5653",
X"76802eb5",
X"387452ff",
X"1651b2c9",
X"3f83e080",
X"08ff1876",
X"54705358",
X"53b2ba3f",
X"83e08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed73f83",
X"e0800853",
X"810b83e0",
X"8008278b",
X"38881408",
X"83e08008",
X"26883880",
X"0b811534",
X"b03983e0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc83f",
X"83e08008",
X"8c3883e0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683e0",
X"800805a8",
X"150c8055",
X"7483e080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83e09808",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1d23f",
X"83e08008",
X"5583e080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef8",
X"3f83e080",
X"0888170c",
X"7551efa9",
X"3f83e080",
X"08557483",
X"e0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683e0",
X"9808802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f83f83e0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"ae8c3f83",
X"e0800841",
X"83e08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"ede23f83",
X"e0800841",
X"83e08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"83a53f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f33f83e0",
X"80088332",
X"70307072",
X"079f2c83",
X"e0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"81b13f75",
X"83e0800c",
X"9e3d0d04",
X"fd3d0d75",
X"77535473",
X"33517089",
X"38713351",
X"70802ea1",
X"38733372",
X"33525372",
X"71278538",
X"ff519439",
X"70732785",
X"3881518b",
X"39811481",
X"135354d3",
X"39805170",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"77545472",
X"337081ff",
X"06525270",
X"802ea338",
X"7181ff06",
X"8114ffbf",
X"12535452",
X"70992689",
X"38a01270",
X"81ff0653",
X"51717470",
X"81055634",
X"d2398074",
X"34853d0d",
X"04ffbd3d",
X"0d80c63d",
X"0852a53d",
X"705254ff",
X"b33f80c7",
X"3d085285",
X"3d705253",
X"ffa63f72",
X"527351fe",
X"df3f80c5",
X"3d0d04fe",
X"3d0d7476",
X"53537170",
X"81055333",
X"51707370",
X"81055534",
X"70f03884",
X"3d0d04fe",
X"3d0d7452",
X"80723352",
X"5370732e",
X"8d388112",
X"81147133",
X"53545270",
X"f5387283",
X"e0800c84",
X"3d0d0471",
X"83e39c0c",
X"8880800b",
X"83e3980c",
X"8480800b",
X"83e3a00c",
X"04fd3d0d",
X"77701755",
X"7705ff1a",
X"535371ff",
X"2e943873",
X"70810555",
X"33517073",
X"70810555",
X"34ff1252",
X"e939853d",
X"0d04fc3d",
X"0d80f6b4",
X"08557433",
X"83e3a434",
X"a05483a0",
X"805383e3",
X"9c085283",
X"e3980851",
X"ffb73fa0",
X"5483a480",
X"5383e39c",
X"085283e3",
X"980851ff",
X"a43f9054",
X"83a88053",
X"83e39c08",
X"5283e398",
X"0851ff91",
X"3fa05380",
X"5283e3a0",
X"0883a080",
X"055185d2",
X"3fa05380",
X"5283e3a0",
X"0883a480",
X"055185c2",
X"3f905380",
X"5283e3a0",
X"0883a880",
X"055185b2",
X"3f80f6b4",
X"0855ff75",
X"3483a080",
X"54805383",
X"e39c0852",
X"83e3a008",
X"51fec63f",
X"80d08054",
X"83b08053",
X"83e39c08",
X"5283e3a0",
X"0851feb1",
X"3f86d33f",
X"a2548053",
X"83e3a008",
X"8c800552",
X"80f4a851",
X"fe9b3f80",
X"f6d80855",
X"86753480",
X"f6dc0855",
X"80753480",
X"f6d40855",
X"80753480",
X"f6c40855",
X"af753480",
X"f6d00855",
X"bf753480",
X"f6cc0855",
X"80753480",
X"f6c80855",
X"9f753480",
X"f6c00855",
X"80753480",
X"f6ac0855",
X"e0753480",
X"f6a40855",
X"a2753480",
X"f6a00855",
X"83753480",
X"f6a80855",
X"82753486",
X"3d0d04fc",
X"3d0d83a0",
X"80548053",
X"83e3a008",
X"5283e39c",
X"0851fda1",
X"3f80d080",
X"5483b080",
X"5383e3a0",
X"085283e3",
X"9c0851fd",
X"8c3fa054",
X"83a08053",
X"83e3a008",
X"5283e39c",
X"0851fcf9",
X"3fa05483",
X"a4805383",
X"e3a00852",
X"83e39c08",
X"51fce63f",
X"905483a8",
X"805383e3",
X"a0085283",
X"e39c0851",
X"fcd33f80",
X"f6b40855",
X"83e3a433",
X"7534863d",
X"0d04803d",
X"0d80f7bc",
X"08700881",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d80f7bc",
X"08700870",
X"fe067607",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"f7bc0870",
X"0870812c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"ff3d0d80",
X"f7bc0870",
X"0870fd06",
X"76100772",
X"0c525283",
X"3d0d0480",
X"3d0d80f7",
X"bc087008",
X"70822cbf",
X"0683e080",
X"0c515182",
X"3d0d04ff",
X"3d0d80f7",
X"bc087008",
X"70fe8306",
X"76822b07",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"f7bc0870",
X"0870882c",
X"870683e0",
X"800c5151",
X"823d0d04",
X"ff3d0d80",
X"f7bc0870",
X"0870f1ff",
X"0676882b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80f7bc08",
X"7008708b",
X"2cbf0683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80f7bc08",
X"700870f8",
X"8fff0676",
X"8b2b0772",
X"0c525283",
X"3d0d0480",
X"3d0d80f7",
X"bc087008",
X"70912cbf",
X"0683e080",
X"0c515182",
X"3d0d04ff",
X"3d0d80f7",
X"bc087008",
X"70fc87ff",
X"ff067691",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d80f7cc",
X"08700870",
X"882c8106",
X"83e0800c",
X"5151823d",
X"0d04803d",
X"0d80f7cc",
X"08700870",
X"892c8106",
X"83e0800c",
X"5151823d",
X"0d04803d",
X"0d80f7cc",
X"08700870",
X"8a2c8106",
X"83e0800c",
X"5151823d",
X"0d04803d",
X"0d80f7cc",
X"08700870",
X"8b2c8106",
X"83e0800c",
X"5151823d",
X"0d04fd3d",
X"0d7581e6",
X"29872a80",
X"f7ac0854",
X"730c853d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"81055434",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727084",
X"05540cff",
X"1151f039",
X"843d0d04",
X"fe3d0d84",
X"80805380",
X"5288800a",
X"51ffb33f",
X"81808053",
X"80528280",
X"0a51c63f",
X"843d0d04",
X"803d0d81",
X"51fc9b3f",
X"72802e83",
X"38d23f81",
X"51fcbd3f",
X"8051fcb8",
X"3f8051fc",
X"853f823d",
X"0d04fd3d",
X"0d755280",
X"5480ff72",
X"25883881",
X"0bff8013",
X"5354ffbf",
X"12517099",
X"268638e0",
X"12529e39",
X"ff9f1251",
X"99712795",
X"38d012e0",
X"13705454",
X"51897127",
X"88388f73",
X"27833880",
X"5273802e",
X"85388180",
X"12527181",
X"ff0683e0",
X"800c853d",
X"0d04803d",
X"0d84d8c0",
X"51807170",
X"81055334",
X"7084e0c0",
X"2e098106",
X"f038823d",
X"0d04fe3d",
X"0d029705",
X"3351ff86",
X"3f83e080",
X"0881ff06",
X"83e3a808",
X"54528073",
X"249b3883",
X"e3c40813",
X"7283e3c8",
X"08075353",
X"71733483",
X"e3a80881",
X"0583e3a8",
X"0c843d0d",
X"04fa3d0d",
X"82800a1b",
X"55805788",
X"3dfc0554",
X"79537452",
X"7851d5d6",
X"3f883d0d",
X"04fe3d0d",
X"83e3c008",
X"527451dc",
X"bb3f83e0",
X"80088c38",
X"76537552",
X"83e3c008",
X"51c73f84",
X"3d0d04fe",
X"3d0d83e3",
X"c0085375",
X"527451d6",
X"f93f83e0",
X"80088d38",
X"77537652",
X"83e3c008",
X"51ffa23f",
X"843d0d04",
X"fe3d0d83",
X"e3c00851",
X"d5ed3f83",
X"e0800881",
X"80802e09",
X"81068838",
X"83c18080",
X"539b3983",
X"e3c00851",
X"d5d13f83",
X"e0800880",
X"d0802e09",
X"81069338",
X"83c1b080",
X"5383e080",
X"085283e3",
X"c00851fe",
X"d83f843d",
X"0d04803d",
X"0dfa993f",
X"83e08008",
X"842980f4",
X"cc057008",
X"83e0800c",
X"51823d0d",
X"04ee3d0d",
X"80438042",
X"80418070",
X"5a5bfdd2",
X"3f800b83",
X"e3a80c80",
X"0b83e3c8",
X"0c80f2a8",
X"51d0bb3f",
X"81800b83",
X"e3c80c80",
X"f2ac51d0",
X"ad3f80d0",
X"0b83e3a8",
X"0c783070",
X"7a078025",
X"70872b83",
X"e3c80c51",
X"55f9883f",
X"83e08008",
X"5280f2b4",
X"51d0873f",
X"80f80b83",
X"e3a80c78",
X"81327030",
X"70720780",
X"2570872b",
X"83e3c80c",
X"515656fe",
X"f13f83e0",
X"80085280",
X"f2c051cf",
X"dd3f81a0",
X"0b83e3a8",
X"0c788232",
X"70307072",
X"07802570",
X"872b83e3",
X"c80c5156",
X"83e3c008",
X"5256d0f7",
X"3f83e080",
X"085280f2",
X"c851cfae",
X"3f81f00b",
X"83e3a80c",
X"810b83e3",
X"ac5b5883",
X"e3a80882",
X"197a3270",
X"30707207",
X"80257087",
X"2b83e3c8",
X"0c51578e",
X"3d7055ff",
X"1b545757",
X"5799873f",
X"79708405",
X"5b0851d0",
X"ae3f7454",
X"83e08008",
X"53775280",
X"f2d051ce",
X"e13fa817",
X"83e3a80c",
X"81185877",
X"852e0981",
X"06ffb038",
X"83900b83",
X"e3a80c78",
X"87327030",
X"70720780",
X"2570872b",
X"83e3c80c",
X"515656f8",
X"ba3f80f2",
X"e05583e0",
X"8008802e",
X"8e3883e3",
X"bc0851cf",
X"da3f83e0",
X"80085574",
X"5280f2e8",
X"51ce8f3f",
X"83e00b83",
X"e3a80c78",
X"88327030",
X"70720780",
X"2570872b",
X"83e3c80c",
X"515780f2",
X"f45255cd",
X"ed3f868d",
X"a051f982",
X"3f805291",
X"3d705255",
X"99df3f83",
X"52745199",
X"d83f6119",
X"59788025",
X"85388059",
X"90398879",
X"25853888",
X"59873978",
X"882682db",
X"3878822b",
X"5580f184",
X"150804f6",
X"a23f83e0",
X"80086157",
X"5575812e",
X"09810689",
X"3883e080",
X"08105590",
X"3975ff2e",
X"09810688",
X"3883e080",
X"08812c55",
X"90752585",
X"38905588",
X"39748024",
X"83388155",
X"7451f5ff",
X"3f829039",
X"f6923f83",
X"e0800861",
X"05557480",
X"25853880",
X"55883987",
X"75258338",
X"87557451",
X"f68e3f81",
X"ee396087",
X"3862802e",
X"81e53883",
X"e0a40883",
X"e0a00c8c",
X"830b83e0",
X"a80c83e3",
X"c00851ff",
X"bed73ffa",
X"e73f81c7",
X"39605680",
X"76259938",
X"8b9c0b83",
X"e0a80c83",
X"e3a01570",
X"085255ff",
X"beb73f74",
X"08529139",
X"75802591",
X"3883e3a0",
X"150851cd",
X"c83f8052",
X"fd1951b8",
X"3962802e",
X"818d3883",
X"e3a01570",
X"0883e3ac",
X"08720c83",
X"e3ac0cfd",
X"1a705351",
X"558af83f",
X"83e08008",
X"5680518a",
X"ee3f83e0",
X"80085274",
X"51878c3f",
X"75528051",
X"87853f80",
X"d6396055",
X"807525b8",
X"3883e0ac",
X"0883e0a0",
X"0c8c830b",
X"83e0a80c",
X"83e3bc08",
X"51ffbdc1",
X"3f83e3bc",
X"0851ffba",
X"b73f83e0",
X"800881ff",
X"06705255",
X"f5a13f74",
X"802e9c38",
X"8155a039",
X"74802593",
X"3883e3bc",
X"0851ccb9",
X"3f8051f5",
X"863f8439",
X"6287387a",
X"802efa8a",
X"38805574",
X"83e0800c",
X"943d0d04",
X"fe3d0df5",
X"853f83e0",
X"8008802e",
X"86388051",
X"80f739f5",
X"8d3f83e0",
X"800880eb",
X"38f5b33f",
X"83e08008",
X"802eaa38",
X"8151f2d2",
X"3fefa73f",
X"800b83e3",
X"a80cf9b9",
X"3f83e080",
X"0853ff0b",
X"83e3a80c",
X"f1b13f72",
X"be387251",
X"f2b03fbc",
X"39f4e73f",
X"83e08008",
X"802eb138",
X"8151f29e",
X"3feef33f",
X"8b9c0b83",
X"e0a80c83",
X"e3ac0851",
X"ffbc863f",
X"ff0b83e3",
X"a80cf0fb",
X"3f83e3ac",
X"08528051",
X"85953f81",
X"51f5d13f",
X"843d0d04",
X"fc3d0d90",
X"80805286",
X"84808051",
X"cf8e3f83",
X"e0800880",
X"c33888e0",
X"3f80f7d0",
X"51d3cf3f",
X"83e08008",
X"559c800a",
X"5480c080",
X"5380f2fc",
X"5283e080",
X"0851f79f",
X"3f83e3c0",
X"085380f3",
X"8c527451",
X"ce983f83",
X"e0800884",
X"38f7ad3f",
X"8151f4f8",
X"3f92eb3f",
X"8151f4f0",
X"3ffe913f",
X"fc3983e0",
X"8c080283",
X"e08c0cfb",
X"3d0d0280",
X"f3980b83",
X"e0a40c80",
X"f39c0b83",
X"e09c0c80",
X"f3a00b83",
X"e0ac0c83",
X"e08c08fc",
X"050c800b",
X"83e3ac0b",
X"83e08c08",
X"f8050c83",
X"e08c08f4",
X"050cccf0",
X"3f83e080",
X"088605fc",
X"0683e08c",
X"08f0050c",
X"0283e08c",
X"08f00508",
X"310d833d",
X"7083e08c",
X"08f80508",
X"70840583",
X"e08c08f8",
X"050c0c51",
X"c9b73f83",
X"e08c08f4",
X"05088105",
X"83e08c08",
X"f4050c83",
X"e08c08f4",
X"0508862e",
X"098106ff",
X"ad388694",
X"808051ec",
X"8a3fff0b",
X"83e3a80c",
X"800b83e3",
X"c80c84d8",
X"c00b83e3",
X"c40c8151",
X"efd83f81",
X"51f0813f",
X"8051effc",
X"3f8151f0",
X"a63f8151",
X"f1833f82",
X"51f0cd3f",
X"8051f1ab",
X"3f80c7aa",
X"528051c6",
X"f63ffdc0",
X"3f83e08c",
X"08fc0508",
X"0d800b83",
X"e0800c87",
X"3d0d83e0",
X"8c0c0480",
X"3d0d81ff",
X"51800b83",
X"e3d41234",
X"ff115170",
X"f438823d",
X"0d04ff3d",
X"0d737033",
X"53518111",
X"33713471",
X"81123483",
X"3d0d04fb",
X"3d0d7779",
X"56568070",
X"71555552",
X"717525ac",
X"38721670",
X"33701470",
X"81ff0655",
X"51515171",
X"74278938",
X"81127081",
X"ff065351",
X"71811470",
X"83ffff06",
X"55525474",
X"7324d638",
X"7183e080",
X"0c873d0d",
X"04fc3d0d",
X"7655c0a0",
X"3f83e080",
X"08802ef6",
X"3883e5f0",
X"08860570",
X"81ff0652",
X"53ffbdf8",
X"3f8439fb",
X"833fc080",
X"3f83e080",
X"08812ef3",
X"38805473",
X"1553ffbe",
X"d53f83e0",
X"80087334",
X"81145473",
X"852e0981",
X"06e93884",
X"39fad93f",
X"ffbfd53f",
X"83e08008",
X"802ef238",
X"743383e3",
X"d4348115",
X"3383e3d5",
X"34821533",
X"83e3d634",
X"83153383",
X"e3d73484",
X"5283e3d4",
X"51febc3f",
X"83e08008",
X"81ff0684",
X"16335653",
X"72752e09",
X"81068d38",
X"ffbec53f",
X"83e08008",
X"802e9a38",
X"83e5f008",
X"a82e0981",
X"06893886",
X"0b83e5f0",
X"0c8739a8",
X"0b83e5f0",
X"0c80e451",
X"efd43f86",
X"3d0d04f4",
X"3d0d7e60",
X"5955805d",
X"8075822b",
X"7183e5f4",
X"120c83e6",
X"88175b5b",
X"57767934",
X"77772e83",
X"b2387652",
X"7751c886",
X"3f8e3dfc",
X"05549053",
X"83e5dc52",
X"7751c7c2",
X"3f7c5675",
X"902e0981",
X"06839038",
X"83e5dc51",
X"fd983f83",
X"e5de51fd",
X"913f83e5",
X"e051fd8a",
X"3f7683e5",
X"ec0c7751",
X"c58d3f80",
X"f1b85283",
X"e0800851",
X"ffb4933f",
X"83e08008",
X"812e0981",
X"0680d338",
X"7683e684",
X"0c820b83",
X"e5dc34ff",
X"960b83e5",
X"dd347751",
X"c7d53f83",
X"e0800855",
X"83e08008",
X"77258838",
X"83e08008",
X"8f055574",
X"842c7083",
X"ffff0670",
X"882a5851",
X"557583e5",
X"de347483",
X"e5df3476",
X"83e5e034",
X"ff800b83",
X"e5e13481",
X"8f3983e5",
X"dc3383e5",
X"dd337188",
X"2b07565b",
X"7483ffff",
X"2e098106",
X"80e738fe",
X"800b83e6",
X"840c810b",
X"83e5ec0c",
X"ff0b83e5",
X"dc34ff0b",
X"83e5dd34",
X"7751c6e3",
X"3f83e080",
X"0883e68c",
X"0c83e080",
X"085583e0",
X"80088025",
X"883883e0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83e5de34",
X"7483e5df",
X"347683e5",
X"e034ff80",
X"0b83e5e1",
X"34810b83",
X"e5eb34a4",
X"39748596",
X"2e098106",
X"80fd3875",
X"83e6840c",
X"7751c698",
X"3f83e5eb",
X"3383e080",
X"08075574",
X"83e5eb34",
X"83e5eb33",
X"81065574",
X"802e8338",
X"845783e5",
X"e03383e5",
X"e1337188",
X"2b07565c",
X"7481802e",
X"098106a1",
X"3883e5de",
X"3383e5df",
X"3371882b",
X"07565bad",
X"80752787",
X"38768207",
X"579c3976",
X"81075796",
X"39748280",
X"2e098106",
X"87387683",
X"07578739",
X"7481ff26",
X"8a387783",
X"e5f41b0c",
X"7679348e",
X"3d0d0480",
X"3d0d7284",
X"2983e5f4",
X"05700883",
X"e0800c51",
X"823d0d04",
X"fe3d0d80",
X"0b83e5d8",
X"0c800b83",
X"e5d40cff",
X"0b83e3d0",
X"0ca80b83",
X"e5f00cae",
X"51ffb8c8",
X"3f800b83",
X"e5f45452",
X"80737084",
X"05550c81",
X"12527184",
X"2e098106",
X"ef38843d",
X"0d04fe3d",
X"0d740284",
X"05960522",
X"53537180",
X"2e973872",
X"70810554",
X"3351ffb8",
X"e63fff12",
X"7083ffff",
X"065152e6",
X"39843d0d",
X"04fe3d0d",
X"02920522",
X"5382ac51",
X"eaec3f80",
X"c351ffb8",
X"c23f8196",
X"51eadf3f",
X"725283e3",
X"d451ffb2",
X"3f725283",
X"e3d451f8",
X"f63f83e0",
X"800881ff",
X"0651ffb8",
X"9e3f843d",
X"0d04ffb1",
X"3d0d80d1",
X"3df80551",
X"f99f3f83",
X"e5d80881",
X"0583e5d8",
X"0c80cf3d",
X"33cf1170",
X"81ff0651",
X"56567483",
X"2688ec38",
X"758f06ff",
X"05567583",
X"e3d0082e",
X"9b387583",
X"26963875",
X"83e3d00c",
X"75842983",
X"e5f40570",
X"08535575",
X"51fa9c3f",
X"80762488",
X"c8387584",
X"2983e5f4",
X"05557408",
X"802e88b9",
X"3883e3d0",
X"08842983",
X"e5f40570",
X"08028805",
X"82b90533",
X"525b5574",
X"80d22e84",
X"b0387480",
X"d2249038",
X"74bf2e9c",
X"387480d0",
X"2e81d738",
X"87f73974",
X"80d32e80",
X"d2387480",
X"d72e81c6",
X"3887e639",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"055656ff",
X"b79f3f80",
X"c151ffb6",
X"d23ff6ef",
X"3f860b83",
X"e3d43481",
X"5283e3d4",
X"51ffb88c",
X"3f8151fd",
X"e43f7489",
X"38860b83",
X"e5f00c87",
X"39a80b83",
X"e5f00cff",
X"b6eb3f80",
X"c151ffb6",
X"9e3ff6bb",
X"3f900b83",
X"e5eb3381",
X"06565674",
X"802e8338",
X"985683e5",
X"e03383e5",
X"e1337188",
X"2b075659",
X"7481802e",
X"0981069c",
X"3883e5de",
X"3383e5df",
X"3371882b",
X"075657ad",
X"8075278c",
X"38758180",
X"07568539",
X"75a00756",
X"7583e3d4",
X"34ff0b83",
X"e3d534e0",
X"0b83e3d6",
X"34800b83",
X"e3d73484",
X"5283e3d4",
X"51ffb780",
X"3f845186",
X"9d390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290556",
X"59ffb5dd",
X"3f7951c0",
X"df3f83e0",
X"8008802e",
X"8b3880ce",
X"51ffb583",
X"3f85f239",
X"80c151ff",
X"b4f93fff",
X"b6803fff",
X"b4833f83",
X"e6840858",
X"8375259b",
X"3883e5e0",
X"3383e5e1",
X"3371882b",
X"07fc1771",
X"297a0583",
X"80055a51",
X"578d3974",
X"81802918",
X"ff800558",
X"81805780",
X"5676762e",
X"9338ffb4",
X"d53f83e0",
X"800883e3",
X"d4173481",
X"1656ea39",
X"ffb4c33f",
X"83e08008",
X"81ff0677",
X"5383e3d4",
X"5256f4df",
X"3f83e080",
X"0881ff06",
X"5575752e",
X"09810681",
X"8a38ffb4",
X"c43f80c1",
X"51ffb3f7",
X"3fffb4fe",
X"3f775279",
X"51ffbeee",
X"3f805e80",
X"d13dfdf4",
X"05547653",
X"83e3d452",
X"7951ffbc",
X"fa3f0282",
X"b9053355",
X"81587480",
X"d72e0981",
X"06bd3880",
X"d13dfdf0",
X"05547653",
X"8f3d7053",
X"7a5259ff",
X"be803f80",
X"5676762e",
X"a2387519",
X"83e3d417",
X"33713370",
X"72327030",
X"70802570",
X"307e0681",
X"1d5d5e51",
X"5151525b",
X"55db3982",
X"ac51e5a6",
X"3f77802e",
X"863880c3",
X"51843980",
X"ce51ffb2",
X"f23fffb3",
X"f93fffb1",
X"fc3f83dd",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055955",
X"80705d59",
X"ffb3923f",
X"80c151ff",
X"b2c53f83",
X"e5ec0879",
X"2e82de38",
X"83e68c08",
X"80fc0555",
X"80fd5274",
X"5188963f",
X"83e08008",
X"5b778224",
X"b238ff18",
X"70872b83",
X"ffff8006",
X"80f4ec05",
X"83e3d459",
X"57558180",
X"55757081",
X"05573377",
X"70810559",
X"34ff1570",
X"81ff0651",
X"5574ea38",
X"828d3977",
X"82e82e81",
X"ab387782",
X"e92e0981",
X"0681b238",
X"80f3a451",
X"ffb8df3f",
X"78587787",
X"32703070",
X"72078025",
X"7a8a3270",
X"30707207",
X"80257307",
X"53545a51",
X"57557580",
X"2e973878",
X"78269238",
X"a00b83e3",
X"d41a3481",
X"197081ff",
X"065a55eb",
X"39811870",
X"81ff0659",
X"558a7827",
X"ffbc388f",
X"5883e3cf",
X"183383e3",
X"d41934ff",
X"187081ff",
X"06595577",
X"8426ea38",
X"9058800b",
X"83e3d419",
X"34811870",
X"81ff0670",
X"982b5259",
X"55748025",
X"e93880c6",
X"557a858f",
X"24843880",
X"c2557483",
X"e3d43480",
X"f10b83e3",
X"d734810b",
X"83e3d834",
X"7a83e3d5",
X"347a882c",
X"557483e3",
X"d63480cb",
X"3982f078",
X"2580c438",
X"7780fd29",
X"fd97d305",
X"527951ff",
X"bb9c3f80",
X"d13dfdec",
X"055480fd",
X"5383e3d4",
X"527951ff",
X"bad43f7b",
X"81195956",
X"7580fc24",
X"83387858",
X"77882c55",
X"7483e4d1",
X"347783e4",
X"d2347583",
X"e4d33481",
X"805980cc",
X"3983e684",
X"08578378",
X"259b3883",
X"e5e03383",
X"e5e13371",
X"882b07fc",
X"1a712979",
X"05838005",
X"5951598d",
X"39778180",
X"2917ff80",
X"05578180",
X"59765279",
X"51ffbaaa",
X"3f80d13d",
X"fdec0554",
X"785383e3",
X"d4527951",
X"ffb9e33f",
X"7851f6b9",
X"3fffb096",
X"3fffae99",
X"3f8b3983",
X"e5d40881",
X"0583e5d4",
X"0c80d13d",
X"0d04f6da",
X"3feba93f",
X"f939fc3d",
X"0d767871",
X"842983e5",
X"f4057008",
X"51535353",
X"709e3880",
X"ce723480",
X"cf0b8113",
X"3480ce0b",
X"82133480",
X"c50b8313",
X"34708413",
X"3480e739",
X"83e68813",
X"335480d2",
X"72347382",
X"2a708106",
X"515180cf",
X"53708438",
X"80d75372",
X"811334a0",
X"0b821334",
X"73830651",
X"70812e9e",
X"38708124",
X"88387080",
X"2e8f389f",
X"3970822e",
X"92387083",
X"2e923893",
X"3980d855",
X"8e3980d3",
X"55893980",
X"cd558439",
X"80c45574",
X"83133480",
X"c40b8413",
X"34800b85",
X"1334863d",
X"0d04fd3d",
X"0d755480",
X"740c800b",
X"84150c80",
X"0b88150c",
X"80f6b808",
X"70337081",
X"ff067081",
X"2a813271",
X"81327181",
X"06718106",
X"31841a0c",
X"56567083",
X"2a813271",
X"822a8132",
X"71810671",
X"81063179",
X"0c525551",
X"515180f6",
X"b0087033",
X"70098106",
X"88170c51",
X"51853d0d",
X"04fe3d0d",
X"74765452",
X"7151ff9a",
X"3f72812e",
X"a2388173",
X"268d3872",
X"822eab38",
X"72832e9f",
X"38e63971",
X"08e23884",
X"1208dd38",
X"881208d8",
X"38a03988",
X"1208812e",
X"098106cc",
X"38943988",
X"1208812e",
X"8d387108",
X"89388412",
X"08802eff",
X"b738843d",
X"0d04fd3d",
X"0d755473",
X"83e69408",
X"2ea73880",
X"f7b00874",
X"a00a0771",
X"0c80f7c0",
X"08535371",
X"08517080",
X"2ef93880",
X"730c7108",
X"5170fb38",
X"7383e694",
X"0c853d0d",
X"04ff0b83",
X"e6940c81",
X"80800b83",
X"e6900c80",
X"0b83e080",
X"0c04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"9d3f7280",
X"2ea33883",
X"e6900814",
X"52713375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552da",
X"39800b83",
X"e0800c86",
X"3d0d04f7",
X"3d0d7b7d",
X"7f115855",
X"59805573",
X"762eb138",
X"83e69008",
X"8b3d5957",
X"74197033",
X"75fc0619",
X"70085d76",
X"83067b07",
X"53545451",
X"72713479",
X"720c8114",
X"81165654",
X"73762e09",
X"8106d938",
X"800b83e0",
X"800c8b3d",
X"0d04fe3d",
X"0d80f7b0",
X"0883e694",
X"08900a07",
X"710c80f7",
X"c0085353",
X"71085170",
X"802ef938",
X"80730c71",
X"085170fb",
X"38843d0d",
X"0483e08c",
X"080283e0",
X"8c0cfd3d",
X"0d805383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"05085183",
X"d43f83e0",
X"80087083",
X"e0800c54",
X"853d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cfd3d0d",
X"815383e0",
X"8c088c05",
X"085283e0",
X"8c088805",
X"085183a1",
X"3f83e080",
X"087083e0",
X"800c5485",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"f93d0d80",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"88050880",
X"25b93883",
X"e08c0888",
X"05083083",
X"e08c0888",
X"050c800b",
X"83e08c08",
X"f4050c83",
X"e08c08fc",
X"05088a38",
X"810b83e0",
X"8c08f405",
X"0c83e08c",
X"08f40508",
X"83e08c08",
X"fc050c83",
X"e08c088c",
X"05088025",
X"b93883e0",
X"8c088c05",
X"083083e0",
X"8c088c05",
X"0c800b83",
X"e08c08f0",
X"050c83e0",
X"8c08fc05",
X"088a3881",
X"0b83e08c",
X"08f0050c",
X"83e08c08",
X"f0050883",
X"e08c08fc",
X"050c8053",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"81df3f83",
X"e0800870",
X"83e08c08",
X"f8050c54",
X"83e08c08",
X"fc050880",
X"2e903883",
X"e08c08f8",
X"05083083",
X"e08c08f8",
X"050c83e0",
X"8c08f805",
X"087083e0",
X"800c5489",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"fb3d0d80",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"88050880",
X"25993883",
X"e08c0888",
X"05083083",
X"e08c0888",
X"050c810b",
X"83e08c08",
X"fc050c83",
X"e08c088c",
X"05088025",
X"903883e0",
X"8c088c05",
X"083083e0",
X"8c088c05",
X"0c815383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"050851bd",
X"3f83e080",
X"087083e0",
X"8c08f805",
X"0c5483e0",
X"8c08fc05",
X"08802e90",
X"3883e08c",
X"08f80508",
X"3083e08c",
X"08f8050c",
X"83e08c08",
X"f8050870",
X"83e0800c",
X"54873d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cfd3d",
X"0d810b83",
X"e08c08fc",
X"050c800b",
X"83e08c08",
X"f8050c83",
X"e08c088c",
X"050883e0",
X"8c088805",
X"0827b938",
X"83e08c08",
X"fc050880",
X"2eae3880",
X"0b83e08c",
X"088c0508",
X"24a23883",
X"e08c088c",
X"05081083",
X"e08c088c",
X"050c83e0",
X"8c08fc05",
X"081083e0",
X"8c08fc05",
X"0cffb839",
X"83e08c08",
X"fc050880",
X"2e80e138",
X"83e08c08",
X"8c050883",
X"e08c0888",
X"050826ad",
X"3883e08c",
X"08880508",
X"83e08c08",
X"8c050831",
X"83e08c08",
X"88050c83",
X"e08c08f8",
X"050883e0",
X"8c08fc05",
X"080783e0",
X"8c08f805",
X"0c83e08c",
X"08fc0508",
X"812a83e0",
X"8c08fc05",
X"0c83e08c",
X"088c0508",
X"812a83e0",
X"8c088c05",
X"0cff9539",
X"83e08c08",
X"90050880",
X"2e933883",
X"e08c0888",
X"05087083",
X"e08c08f4",
X"050c5191",
X"3983e08c",
X"08f80508",
X"7083e08c",
X"08f4050c",
X"5183e08c",
X"08f40508",
X"83e0800c",
X"853d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cff3d0d",
X"800b83e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"8106ff11",
X"70097083",
X"e08c088c",
X"05080683",
X"e08c08fc",
X"05081183",
X"e08c08fc",
X"050c83e0",
X"8c088805",
X"08812a83",
X"e08c0888",
X"050c83e0",
X"8c088c05",
X"081083e0",
X"8c088c05",
X"0c515151",
X"5183e08c",
X"08880508",
X"802e8438",
X"ffab3983",
X"e08c08fc",
X"05087083",
X"e0800c51",
X"833d0d83",
X"e08c0c04",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"0000265b",
X"0000269c",
X"000026be",
X"000026e5",
X"000026e5",
X"000026e5",
X"000026e5",
X"00002756",
X"000027a8",
X"25732025",
X"73000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"6e616d65",
X"20000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"000038e4",
X"000038e8",
X"000038f0",
X"000038fc",
X"00003908",
X"00003914",
X"00003920",
X"00003924",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"0001d20f",
X"0001d400",
X"0001d401",
X"0001d409",
X"0001d010",
X"0001d301",
X"0001d300",
X"0001d20a",
X"0001d01b",
X"0001d016",
X"0001d019",
X"0001d018",
X"0001d017",
X"0001d01a",
X"0001d403",
X"0001d402",
X"0001d40e",
X"0004007c",
X"00040078",
X"00040074",
X"00040068",
X"00040060",
X"0004005c",
X"00040058",
X"00040054",
X"00040050",
X"0004004c",
X"00040048",
X"00040044",
X"00040040",
X"00040034",
X"00040030",
X"0004002c",
X"00040028",
X"00040024",
X"00040020",
X"0004001c",
X"00040018",
X"00040014",
X"00040010",
X"0004000c",
X"00040008",
X"00040004",
X"00040000",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
