
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81d4",
X"b4738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81dc",
X"a40c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757580f2",
X"952d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7580f1d4",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80dca004",
X"fd3d0d75",
X"705254ae",
X"a73f83c0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"c0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83c0",
X"8008732e",
X"a13883c0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183c0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83c2d008",
X"248a38b4",
X"f83fff0b",
X"83c2d00c",
X"800b83c0",
X"800c04ff",
X"3d0d7352",
X"83c0ac08",
X"722e8d38",
X"d93f7151",
X"96993f71",
X"83c0ac0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"558154bc",
X"15088191",
X"387451cf",
X"3f795880",
X"7a2580f7",
X"3883c380",
X"0870892a",
X"5783ff06",
X"78848072",
X"31565657",
X"73782583",
X"38735575",
X"83c2d008",
X"2e8438ff",
X"893f83c2",
X"d0088025",
X"a6387589",
X"2b5198dc",
X"3f83c380",
X"088f3dfc",
X"11555c54",
X"8152f81b",
X"5196c63f",
X"761483c3",
X"800c7583",
X"c2d00c74",
X"53765278",
X"51b3a93f",
X"83c08008",
X"83c38008",
X"1683c380",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8b3861",
X"7a710c54",
X"75547580",
X"2e833881",
X"547383c0",
X"800c8e3d",
X"0d04fc3d",
X"0dfe9b3f",
X"7651feaf",
X"3f863dfc",
X"05537852",
X"775195e9",
X"3f797571",
X"0c5483c0",
X"80085483",
X"c0800880",
X"2e833881",
X"547383c0",
X"800c863d",
X"0d04fe3d",
X"0d7583c2",
X"d0085353",
X"80722489",
X"3871732e",
X"8438fdd6",
X"3f7451fd",
X"ea3f7251",
X"97ae3f83",
X"c0800852",
X"83c08008",
X"802e8338",
X"81527183",
X"c0800c84",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"c0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"c0800c51",
X"823d0d04",
X"80c40b83",
X"c0800c04",
X"fd3d0d75",
X"77715470",
X"535553a9",
X"ff3f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfceb3f",
X"735193ab",
X"3f7383c0",
X"ac0c83c0",
X"80085383",
X"c0800880",
X"2e833881",
X"537283c0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcbf3f",
X"72802ea5",
X"38bc1308",
X"527351a9",
X"893f83c0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"c0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83c0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83c2d0",
X"0c7483c0",
X"b00c7583",
X"c2cc0caf",
X"dd3f83c0",
X"800881ff",
X"06528153",
X"71993883",
X"c2e8518e",
X"943f83c0",
X"80085283",
X"c0800880",
X"2e833872",
X"52715372",
X"83c0800c",
X"843d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"51a6fa3f",
X"83c08008",
X"557483c0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"c0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283c2cc",
X"085180e0",
X"d73f83c0",
X"800857f9",
X"e13f7952",
X"83c2d451",
X"95b73f83",
X"c0800854",
X"805383c0",
X"8008732e",
X"09810682",
X"833883c0",
X"b0080b0b",
X"81d9c053",
X"705256a6",
X"b73f0b0b",
X"81d9c052",
X"80c01651",
X"a6aa3f75",
X"bc170c73",
X"82c0170c",
X"810b82c4",
X"170c810b",
X"82c8170c",
X"7382cc17",
X"0cff1782",
X"d0175557",
X"81913983",
X"c0bc3370",
X"822a7081",
X"06515455",
X"72818038",
X"74812a81",
X"06587780",
X"f6387484",
X"2a810682",
X"c4150c83",
X"c0bc3381",
X"0682c815",
X"0c795273",
X"51a5d13f",
X"7351a5e8",
X"3f83c080",
X"081453af",
X"73708105",
X"553472bc",
X"150c83c0",
X"bd527251",
X"a5b23f83",
X"c0b40882",
X"c0150c83",
X"c0ca5280",
X"c01451a5",
X"9f3f7880",
X"2e8d3873",
X"51782d83",
X"c0800880",
X"2e993877",
X"82cc150c",
X"75802e86",
X"387382cc",
X"170c7382",
X"d015ff19",
X"59555676",
X"802e9b38",
X"83c0b452",
X"83c2d451",
X"94ad3f83",
X"c080088a",
X"3883c0bd",
X"335372fe",
X"d2387880",
X"2e893883",
X"c0b00851",
X"fcb83f83",
X"c0b00853",
X"7283c080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb53f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f690",
X"3f83c080",
X"08745387",
X"3d705355",
X"55f6b03f",
X"f7903f73",
X"51d33f63",
X"53745283",
X"c0800851",
X"fab83f92",
X"3d0d0471",
X"83c0800c",
X"0480c012",
X"83c0800c",
X"04803d0d",
X"7282c011",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"c0800c51",
X"823d0d04",
X"f93d0d79",
X"83c09008",
X"57578177",
X"27819638",
X"76881708",
X"27818e38",
X"75335574",
X"822e8938",
X"74832eb3",
X"3880fe39",
X"74547610",
X"83fe0653",
X"76882a8c",
X"17080552",
X"893dfc05",
X"51aa8b3f",
X"83c08008",
X"80df3802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d13984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"51a9db3f",
X"83c08008",
X"b038029f",
X"05330284",
X"059e0533",
X"71982b71",
X"902b0702",
X"8c059d05",
X"3370882b",
X"72078d3d",
X"337180ff",
X"fffe8006",
X"07515253",
X"57585683",
X"39815574",
X"83c0800c",
X"893d0d04",
X"fb3d0d83",
X"c09008fe",
X"19881208",
X"fe055556",
X"54805674",
X"73278d38",
X"82143375",
X"71299416",
X"08055753",
X"7583c080",
X"0c873d0d",
X"04fc3d0d",
X"7652800b",
X"83c09008",
X"70335152",
X"5370832e",
X"09810691",
X"38951233",
X"94133371",
X"982b7190",
X"2b075555",
X"519b1233",
X"9a133371",
X"882b0774",
X"0783c080",
X"0c55863d",
X"0d04fc3d",
X"0d7683c0",
X"90085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"fed63f83",
X"c0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183c080",
X"0c863d0d",
X"04fa3d0d",
X"7883c090",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fcb13f",
X"81527183",
X"c0800827",
X"a8388352",
X"83c08008",
X"88170827",
X"9c3883c0",
X"80088c16",
X"0c83c080",
X"0851fdbc",
X"3f83c080",
X"0890160c",
X"73752380",
X"527183c0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585e5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"9f269138",
X"7a51fdd2",
X"3f83c080",
X"0856807d",
X"34838139",
X"933d841c",
X"08705859",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"3880705a",
X"5c887f08",
X"5f5a7b81",
X"1d7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535e57",
X"557480e7",
X"3876ae2e",
X"09810683",
X"38815578",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675bb",
X"3888598b",
X"5affab39",
X"76982b55",
X"74802587",
X"3881d3c4",
X"173357ff",
X"9f175574",
X"99268938",
X"e0177081",
X"ff065855",
X"78811a70",
X"81ff0672",
X"1b535b57",
X"55767534",
X"fef8397b",
X"1e7f0c80",
X"5576a026",
X"83388155",
X"748b1934",
X"7a51fc82",
X"3f83c080",
X"0880f538",
X"a0547a22",
X"70852b83",
X"e0065455",
X"901b0852",
X"7c51a496",
X"3f83c080",
X"085783c0",
X"80088181",
X"387c3355",
X"74802e80",
X"f4388b1d",
X"3370832a",
X"70810651",
X"565674b4",
X"388b7d84",
X"1d0883c0",
X"8008595b",
X"5b58ff18",
X"5877ff2e",
X"9a387970",
X"81055b33",
X"79708105",
X"5b337171",
X"31525656",
X"75802ee2",
X"38863975",
X"802e9638",
X"7a51fbe5",
X"3fff8639",
X"83c08008",
X"5683c080",
X"08b63883",
X"39765684",
X"1b088b11",
X"33515574",
X"a7388b1d",
X"3370842a",
X"70810651",
X"56567489",
X"38835694",
X"39815690",
X"397c51fa",
X"943f83c0",
X"8008881c",
X"0cfd8139",
X"7583c080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"51a2db3f",
X"835683c0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"51a2af3f",
X"83c08008",
X"98388117",
X"33773371",
X"882b0783",
X"c0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"7651a286",
X"3f83c080",
X"08983881",
X"17337733",
X"71882b07",
X"83c08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583c080",
X"0c8a3d0d",
X"04eb3d0d",
X"675a800b",
X"83c0900c",
X"a1a83f83",
X"c0800881",
X"06558256",
X"7483ef38",
X"7475538f",
X"3d705357",
X"59feca3f",
X"83c08008",
X"81ff0657",
X"76812e09",
X"810680d4",
X"38905483",
X"be537452",
X"7551a19a",
X"3f83c080",
X"0880c938",
X"8f3d3355",
X"74802e80",
X"c93802bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"33710770",
X"587b575e",
X"525e5759",
X"57fdee3f",
X"83c08008",
X"81ff0657",
X"76832e09",
X"81068638",
X"815682f2",
X"3976802e",
X"86388656",
X"82e839a4",
X"548d5378",
X"527551a0",
X"b13f8156",
X"83c08008",
X"82d43802",
X"be053302",
X"8405bd05",
X"3371882b",
X"07595d77",
X"ab380280",
X"ce053302",
X"840580cd",
X"05337198",
X"2b71902b",
X"07973d33",
X"70882b72",
X"07029405",
X"80cb0533",
X"71075452",
X"5e575956",
X"02b70533",
X"78712902",
X"8805b605",
X"33028c05",
X"b5053371",
X"882b0770",
X"1d707f8c",
X"050c5f59",
X"57595d8e",
X"3d33821b",
X"3402b905",
X"33903d33",
X"71882b07",
X"5a5c7884",
X"1b2302bb",
X"05330284",
X"05ba0533",
X"71882b07",
X"565c74ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"07515253",
X"575e5c74",
X"76317831",
X"79842a90",
X"3d335471",
X"71315356",
X"5680d1bc",
X"3f83c080",
X"08820570",
X"881c0c83",
X"c08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83c0900c",
X"80567583",
X"c0800c97",
X"3d0d04e9",
X"3d0d83c0",
X"90085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e53f83c0",
X"80085483",
X"c0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f489",
X"3f83c080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383c080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83c09008",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0e93f",
X"83c08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"833f83c0",
X"80085583",
X"c0800880",
X"2eff8938",
X"83c08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"519ad73f",
X"83c08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83c0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83c09008",
X"55568555",
X"73802e81",
X"e3388114",
X"33810653",
X"84557280",
X"2e81d538",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b9388214",
X"3370892b",
X"56537680",
X"2eb73874",
X"52ff1651",
X"80ccbd3f",
X"83c08008",
X"ff187654",
X"70535853",
X"80ccad3f",
X"83c08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed63f83",
X"c0800853",
X"810b83c0",
X"8008278b",
X"38881408",
X"83c08008",
X"26883880",
X"0b811534",
X"b03983c0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc53f",
X"83c08008",
X"8c3883c0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683c0",
X"800805a8",
X"150c8055",
X"7483c080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83c09008",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1cf3f",
X"83c08008",
X"5583c080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef5",
X"3f83c080",
X"0888170c",
X"7551efa6",
X"3f83c080",
X"08557483",
X"c0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683c0",
X"9008802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f53f83c0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"96e03f83",
X"c0800841",
X"83c08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"eddf3f83",
X"c0800841",
X"83c08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"8e863f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f03f83c0",
X"80088332",
X"70307072",
X"079f2c83",
X"c0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"8c923f75",
X"83c0800c",
X"9e3d0d04",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"7751e0d2",
X"3f83c080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3381dcac",
X"0b81dcac",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"527751e0",
X"813f83c0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583c0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"558b993f",
X"83c08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"8114518a",
X"b13f83c0",
X"80083070",
X"83c08008",
X"07802583",
X"c0800c53",
X"863d0d04",
X"fc3d0d76",
X"705255e6",
X"ee3f83c0",
X"80085481",
X"5383c080",
X"0880c138",
X"7451e6b1",
X"3f83c080",
X"0881d9d0",
X"5383c080",
X"085253ff",
X"913f83c0",
X"8008a138",
X"81d9d452",
X"7251ff82",
X"3f83c080",
X"08923881",
X"d9d85272",
X"51fef33f",
X"83c08008",
X"802e8338",
X"81547353",
X"7283c080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"e68d3f81",
X"5383c080",
X"08983873",
X"51e5d63f",
X"83c39808",
X"5283c080",
X"0851feba",
X"3f83c080",
X"08537283",
X"c0800c85",
X"3d0d04df",
X"3d0da43d",
X"0870525e",
X"dbfb3f83",
X"c0800833",
X"953d5654",
X"73963881",
X"dffc5274",
X"5189913f",
X"9a397d52",
X"7851defc",
X"3f84d039",
X"7d51dbe1",
X"3f83c080",
X"08527451",
X"db913f80",
X"43804280",
X"41804083",
X"c3a00852",
X"943d7052",
X"5de1e43f",
X"83c08008",
X"59800b83",
X"c0800855",
X"5b83c080",
X"087b2e94",
X"38811b74",
X"525be4e6",
X"3f83c080",
X"085483c0",
X"8008ee38",
X"805aff5f",
X"7909709f",
X"2c7b065b",
X"547a7a24",
X"8438ff1b",
X"5af61a70",
X"09709f2c",
X"72067bff",
X"125a5a52",
X"55558075",
X"25953876",
X"51e4ab3f",
X"83c08008",
X"76ff1858",
X"55577380",
X"24ed3874",
X"7f2e8638",
X"a0bd3f74",
X"5f78ff1b",
X"70585d58",
X"807a2595",
X"387751e4",
X"813f83c0",
X"800876ff",
X"18585558",
X"738024ed",
X"38800b83",
X"c7d00c80",
X"0b83c894",
X"0c81d9dc",
X"518d903f",
X"81800b83",
X"c8940c81",
X"d9e4518d",
X"823fa80b",
X"83c7d00c",
X"76802e80",
X"e43883c7",
X"d0087779",
X"32703070",
X"72078025",
X"70872b83",
X"c8940c51",
X"56785356",
X"56e3b83f",
X"83c08008",
X"802e8838",
X"81d9ec51",
X"8cc93f76",
X"51e2fa3f",
X"83c08008",
X"5281db8c",
X"518cb83f",
X"7651e382",
X"3f83c080",
X"0883c7d0",
X"08555775",
X"74258638",
X"a81656f7",
X"397583c7",
X"d00c86f0",
X"7624ff98",
X"3887980b",
X"83c7d00c",
X"77802eb1",
X"387751e2",
X"b83f83c0",
X"80087852",
X"55e2d83f",
X"81d9f454",
X"83c08008",
X"8d388739",
X"80763481",
X"d03981d9",
X"f0547453",
X"735281d9",
X"c4518bd7",
X"3f805481",
X"d9cc518b",
X"ce3f8114",
X"5473a82e",
X"098106ef",
X"38868da0",
X"519cb03f",
X"8052903d",
X"70525780",
X"c29f3f83",
X"52765180",
X"c2973f62",
X"818f3861",
X"802e80fb",
X"387b5473",
X"ff2e9638",
X"78802e81",
X"8a387851",
X"e1dc3f83",
X"c08008ff",
X"155559e7",
X"3978802e",
X"80f53878",
X"51e1d83f",
X"83c08008",
X"802efc8e",
X"387851e1",
X"a03f83c0",
X"80085281",
X"d9c05183",
X"e43f83c0",
X"8008a338",
X"7c51859c",
X"3f83c080",
X"085574ff",
X"16565480",
X"7425ae38",
X"741d7033",
X"555673af",
X"2efecd38",
X"e9397851",
X"e0e13f83",
X"c0800852",
X"7c5184d4",
X"3f8f397f",
X"88296010",
X"057a0561",
X"055afc90",
X"3962802e",
X"fbd13880",
X"52765180",
X"c0f73fa3",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067084",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d38a8",
X"0b9088b8",
X"34b80b90",
X"88b83470",
X"83c0800c",
X"823d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"852a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"980b9088",
X"b834b80b",
X"9088b834",
X"7083c080",
X"0c823d0d",
X"04930b90",
X"88bc34ff",
X"0b9088a8",
X"3404ff3d",
X"0d028f05",
X"3352800b",
X"9088bc34",
X"8a5199f7",
X"3fdf3f80",
X"f80b9088",
X"a034800b",
X"90888834",
X"fa125271",
X"90888034",
X"800b9088",
X"98347190",
X"88903490",
X"88b85280",
X"7234b872",
X"34833d0d",
X"04803d0d",
X"028b0533",
X"51709088",
X"b434febf",
X"3f83c080",
X"08802ef6",
X"38823d0d",
X"04803d0d",
X"8439a4ae",
X"3ffed93f",
X"83c08008",
X"802ef338",
X"9088b433",
X"7081ff06",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"a30b9088",
X"bc34ff0b",
X"9088a834",
X"9088b851",
X"a87134b8",
X"7134823d",
X"0d04803d",
X"0d9088bc",
X"337081c0",
X"06703070",
X"802583c0",
X"800c5151",
X"51823d0d",
X"04803d0d",
X"9088b833",
X"7081ff06",
X"70832a81",
X"32708106",
X"51515151",
X"70802ee8",
X"38b00b90",
X"88b834b8",
X"0b9088b8",
X"34823d0d",
X"04803d0d",
X"9080ac08",
X"810683c0",
X"800c823d",
X"0d04fd3d",
X"0d757754",
X"54807325",
X"94387370",
X"81055533",
X"5281d9f8",
X"5187843f",
X"ff1353e9",
X"39853d0d",
X"04fd3d0d",
X"75775354",
X"73335170",
X"89387133",
X"5170802e",
X"a1387333",
X"72335253",
X"72712785",
X"38ff5194",
X"39707327",
X"85388151",
X"8b398114",
X"81135354",
X"d3398051",
X"7083c080",
X"0c853d0d",
X"04fd3d0d",
X"75775454",
X"72337081",
X"ff065252",
X"70802ea3",
X"387181ff",
X"068114ff",
X"bf125354",
X"52709926",
X"8938a012",
X"7081ff06",
X"53517174",
X"70810556",
X"34d23980",
X"7434853d",
X"0d04ffbd",
X"3d0d80c6",
X"3d0852a5",
X"3d705254",
X"ffb33f80",
X"c73d0852",
X"853d7052",
X"53ffa63f",
X"72527351",
X"fedf3f80",
X"c53d0d04",
X"fe3d0d74",
X"76535371",
X"70810553",
X"33517073",
X"70810555",
X"3470f038",
X"843d0d04",
X"fe3d0d74",
X"52807233",
X"52537073",
X"2e8d3881",
X"12811471",
X"33535452",
X"70f53872",
X"83c0800c",
X"843d0d04",
X"f63d0d7c",
X"7e60625a",
X"5d5b5680",
X"59815585",
X"39747a29",
X"55745275",
X"51b9913f",
X"83c08008",
X"7a27ee38",
X"74802e80",
X"dd387452",
X"7551b8fc",
X"3f83c080",
X"08755376",
X"5254b980",
X"3f83c080",
X"087a5375",
X"5256b8e4",
X"3f83c080",
X"08793070",
X"7b079f2a",
X"70778024",
X"07515154",
X"55728738",
X"83c08008",
X"c5387681",
X"18b01655",
X"58588974",
X"258b38b7",
X"14537a85",
X"3880d714",
X"53727834",
X"811959ff",
X"9f398077",
X"348c3d0d",
X"04f73d0d",
X"7b7d7f62",
X"029005bb",
X"05335759",
X"565a5ab0",
X"58728338",
X"a0587570",
X"70810552",
X"33715954",
X"55903980",
X"74258e38",
X"ff147770",
X"81055933",
X"545472ef",
X"3873ff15",
X"55538073",
X"25893877",
X"52795178",
X"2def3975",
X"33755753",
X"72802e90",
X"38725279",
X"51782d75",
X"70810557",
X"3353ed39",
X"8b3d0d04",
X"ee3d0d64",
X"66696970",
X"70810552",
X"335b4a5c",
X"5e5e7680",
X"2e82f938",
X"76a52e09",
X"810682e0",
X"38807041",
X"67707081",
X"05523371",
X"4a59575f",
X"76b02e09",
X"81068c38",
X"75708105",
X"57337648",
X"57815fd0",
X"17567589",
X"2680da38",
X"76675c59",
X"805c9339",
X"778a2480",
X"c3387b8a",
X"29187b70",
X"81055d33",
X"5a5cd019",
X"7081ff06",
X"58588977",
X"27a438ff",
X"9f197081",
X"ff06ffa9",
X"1b5a5156",
X"85762792",
X"38ffbf19",
X"7081ff06",
X"51567585",
X"268a38c9",
X"19587780",
X"25ffb938",
X"7a477b40",
X"7881ff06",
X"577680e4",
X"2e80e538",
X"7680e424",
X"a7387680",
X"d82e8186",
X"387680d8",
X"24903876",
X"802e81cc",
X"3876a52e",
X"81b63881",
X"b9397680",
X"e32e818c",
X"3881af39",
X"7680f52e",
X"9b387680",
X"f5248b38",
X"7680f32e",
X"81813881",
X"99397680",
X"f82e80ca",
X"38818f39",
X"913d7055",
X"5780538a",
X"5279841b",
X"7108535b",
X"56fc813f",
X"7655ab39",
X"79841b71",
X"08943d70",
X"5b5b525b",
X"56758025",
X"8c387530",
X"56ad7834",
X"0280c105",
X"57765480",
X"538a5275",
X"51fbd53f",
X"77557e54",
X"b839913d",
X"70557780",
X"d8327030",
X"70802556",
X"51585690",
X"5279841b",
X"7108535b",
X"57fbb13f",
X"7555db39",
X"79841b83",
X"1233545b",
X"56983979",
X"841b7108",
X"575b5680",
X"547f537c",
X"527d51fc",
X"9c3f8739",
X"76527d51",
X"7c2d6670",
X"33588105",
X"47fd8339",
X"943d0d04",
X"7283c094",
X"0c7183c0",
X"980c04fb",
X"3d0d883d",
X"70708405",
X"52085754",
X"755383c0",
X"94085283",
X"c0980851",
X"fcc63f87",
X"3d0d04ff",
X"3d0d7370",
X"08535102",
X"93053372",
X"34700881",
X"05710c83",
X"3d0d04fc",
X"3d0d873d",
X"88115578",
X"54bdbb53",
X"51fc993f",
X"8052873d",
X"51d13f86",
X"3d0d04fc",
X"3d0d7655",
X"7483c3a8",
X"082eaf38",
X"80537451",
X"87c13f83",
X"c0800881",
X"ff06ff14",
X"7081ff06",
X"7230709f",
X"2a515255",
X"53547280",
X"2e843871",
X"dd3873fe",
X"387483c3",
X"a80c863d",
X"0d04ff3d",
X"0dff0b83",
X"c3a80c84",
X"a53f8151",
X"87853f83",
X"c0800881",
X"ff065271",
X"ee3881d3",
X"3f7183c0",
X"800c833d",
X"0d04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"823f7280",
X"2ea03883",
X"c3bc1433",
X"75708105",
X"57348114",
X"7083ffff",
X"06ff1570",
X"83ffff06",
X"56525552",
X"dd39800b",
X"83c0800c",
X"863d0d04",
X"fc3d0d76",
X"787a1156",
X"53558053",
X"71742e93",
X"38721551",
X"703383c3",
X"bc133481",
X"12811454",
X"52ea3980",
X"0b83c080",
X"0c863d0d",
X"04fd3d0d",
X"905483c3",
X"a8085186",
X"f43f83c0",
X"800881ff",
X"06ff1571",
X"30713070",
X"73079f2a",
X"729f2a06",
X"52555255",
X"5372db38",
X"853d0d04",
X"803d0d83",
X"c3b40810",
X"83c3ac08",
X"079080a8",
X"0c823d0d",
X"04800b83",
X"c3b40ce4",
X"3f04810b",
X"83c3b40c",
X"db3f04ed",
X"3f047183",
X"c3b00c04",
X"803d0d80",
X"51f43f81",
X"0b83c3b4",
X"0c810b83",
X"c3ac0cff",
X"bb3f823d",
X"0d04803d",
X"0d723070",
X"74078025",
X"83c3ac0c",
X"51ffa53f",
X"823d0d04",
X"803d0d02",
X"8b053390",
X"80a40c90",
X"80a80870",
X"81065151",
X"70f53890",
X"80a40870",
X"81ff0683",
X"c0800c51",
X"823d0d04",
X"803d0d81",
X"ff51d13f",
X"83c08008",
X"81ff0683",
X"c0800c82",
X"3d0d0480",
X"3d0d7390",
X"2b730790",
X"80b40c82",
X"3d0d0404",
X"fb3d0d78",
X"0284059f",
X"05337098",
X"2b555755",
X"7280259b",
X"387580ff",
X"06568052",
X"80f751e0",
X"3f83c080",
X"0881ff06",
X"54738126",
X"80ff3880",
X"51fee73f",
X"ffa23f81",
X"51fedf3f",
X"ff9a3f75",
X"51feed3f",
X"74982a51",
X"fee63f74",
X"902a7081",
X"ff065253",
X"feda3f74",
X"882a7081",
X"ff065253",
X"fece3f74",
X"81ff0651",
X"fec63f81",
X"557580c0",
X"2e098106",
X"86388195",
X"558d3975",
X"80c82e09",
X"81068438",
X"81875574",
X"51fea53f",
X"8a55fec8",
X"3f83c080",
X"0881ff06",
X"70982b54",
X"54728025",
X"8c38ff15",
X"7081ff06",
X"565374e2",
X"387383c0",
X"800c873d",
X"0d04fa3d",
X"0dfdc53f",
X"8051fdda",
X"3f8a54fe",
X"933fff14",
X"7081ff06",
X"555373f3",
X"38737453",
X"5580c051",
X"fea63f83",
X"c0800881",
X"ff065473",
X"812e0981",
X"06829f38",
X"83aa5280",
X"c851fe8c",
X"3f83c080",
X"0881ff06",
X"5372812e",
X"09810681",
X"a8387454",
X"873d7411",
X"5456fdc8",
X"3f83c080",
X"08733481",
X"147081ff",
X"06555383",
X"7427e538",
X"029a0533",
X"5372812e",
X"09810681",
X"d938029b",
X"05335380",
X"ce905472",
X"81aa2e8d",
X"3881c739",
X"80e4518a",
X"9e3fff14",
X"5473802e",
X"81b83882",
X"0a5281e9",
X"51fda53f",
X"83c08008",
X"81ff0653",
X"72de3872",
X"5280fa51",
X"fd923f83",
X"c0800881",
X"ff065372",
X"81903872",
X"54731653",
X"fcd63f83",
X"c0800873",
X"34811470",
X"81ff0655",
X"53837427",
X"e838873d",
X"3370862a",
X"70810651",
X"54548c55",
X"7280e338",
X"845580de",
X"39745281",
X"e951fccc",
X"3f83c080",
X"0881ff06",
X"53825581",
X"e9568173",
X"27863873",
X"5580c156",
X"80ce9054",
X"8a3980e4",
X"5189903f",
X"ff145473",
X"802ea938",
X"80527551",
X"fc9a3f83",
X"c0800881",
X"ff065372",
X"e1388480",
X"5280d051",
X"fc863f83",
X"c0800881",
X"ff065372",
X"802e8338",
X"80557483",
X"c3b83480",
X"51fb873f",
X"fbc23f88",
X"3d0d04fb",
X"3d0d7754",
X"800b83c3",
X"b8337083",
X"2a708106",
X"51555755",
X"72752e09",
X"81068538",
X"73892b54",
X"735280d1",
X"51fbbd3f",
X"83c08008",
X"81ff0653",
X"72bd3882",
X"b8c054fb",
X"833f83c0",
X"800881ff",
X"06537281",
X"ff2e0981",
X"068938ff",
X"145473e7",
X"389f3972",
X"81fe2e09",
X"81069638",
X"83c7bc52",
X"83c3bc51",
X"faed3ffa",
X"d33ffad0",
X"3f833981",
X"558051fa",
X"893ffac4",
X"3f7481ff",
X"0683c080",
X"0c873d0d",
X"04fb3d0d",
X"7783c3bc",
X"56548151",
X"f9ec3f83",
X"c3b83370",
X"832a7081",
X"06515456",
X"72853873",
X"892b5473",
X"5280d851",
X"fab63f83",
X"c0800881",
X"ff065372",
X"80e43881",
X"ff51f9d4",
X"3f81fe51",
X"f9ce3f84",
X"80537470",
X"81055633",
X"51f9c13f",
X"ff137083",
X"ffff0651",
X"5372eb38",
X"7251f9b0",
X"3f7251f9",
X"ab3ff9d0",
X"3f83c080",
X"089f0653",
X"a7885472",
X"852e8c38",
X"993980e4",
X"5186c83f",
X"ff1454f9",
X"b33f83c0",
X"800881ff",
X"2e843873",
X"e9388051",
X"f8e43ff9",
X"9f3f800b",
X"83c0800c",
X"873d0d04",
X"7183c7c0",
X"0c888080",
X"0b83c7bc",
X"0c848080",
X"0b83c7c4",
X"0c04fd3d",
X"0d777017",
X"557705ff",
X"1a535371",
X"ff2e9438",
X"73708105",
X"55335170",
X"73708105",
X"5534ff12",
X"52e93985",
X"3d0d04fc",
X"3d0d87a6",
X"81557433",
X"83c7c834",
X"a05483a0",
X"805383c7",
X"c0085283",
X"c7bc0851",
X"ffb83fa0",
X"5483a480",
X"5383c7c0",
X"085283c7",
X"bc0851ff",
X"a53f9054",
X"83a88053",
X"83c7c008",
X"5283c7bc",
X"0851ff92",
X"3fa05380",
X"5283c7c4",
X"0883a080",
X"055185a0",
X"3fa05380",
X"5283c7c4",
X"0883a480",
X"05518590",
X"3f905380",
X"5283c7c4",
X"0883a880",
X"05518580",
X"3fff7534",
X"83a08054",
X"805383c7",
X"c0085283",
X"c7c40851",
X"fecc3f80",
X"d0805483",
X"b0805383",
X"c7c00852",
X"83c7c408",
X"51feb73f",
X"86c53fa2",
X"54805383",
X"c7c4088c",
X"80055281",
X"dda051fe",
X"a13f860b",
X"87a88334",
X"800b87a8",
X"8234800b",
X"87a09a34",
X"af0b87a0",
X"9634bf0b",
X"87a09734",
X"800b87a0",
X"98349f0b",
X"87a09934",
X"800b87a0",
X"9b34e00b",
X"87a88934",
X"a20b87a8",
X"8034830b",
X"87a48f34",
X"820b87a8",
X"8134863d",
X"0d04fd3d",
X"0d83a080",
X"54805383",
X"c7c40852",
X"83c7c008",
X"51fdbf3f",
X"80d08054",
X"83b08053",
X"83c7c408",
X"5283c7c0",
X"0851fdaa",
X"3fa05483",
X"a0805383",
X"c7c40852",
X"83c7c008",
X"51fd973f",
X"a05483a4",
X"805383c7",
X"c4085283",
X"c7c00851",
X"fd843f90",
X"5483a880",
X"5383c7c4",
X"085283c7",
X"c00851fc",
X"f13f83c7",
X"c83387a6",
X"8134853d",
X"0d04803d",
X"0d908090",
X"08810683",
X"c0800c82",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe067607",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"812c8106",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fd06",
X"76100772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087082",
X"2cbf0683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fe8306",
X"76822b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"882c8706",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f1ff",
X"0676882b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70912cbf",
X"0683c080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870fc",
X"87ffff06",
X"76912b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"992c8106",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870ffbf",
X"0a067699",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908080",
X"0870882c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"80087089",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8a2c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708b2c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708c2c",
X"bf0683c0",
X"800c5182",
X"3d0d04fe",
X"3d0d7481",
X"e629872a",
X"9080a00c",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d848080",
X"53805288",
X"800a51ff",
X"b33f8180",
X"80538052",
X"82800a51",
X"c63f843d",
X"0d04803d",
X"0d8151fc",
X"aa3f7280",
X"2e903880",
X"51fdfe3f",
X"cd3f83c7",
X"cc3351fd",
X"f43f8151",
X"fcbb3f80",
X"51fcb63f",
X"8051fc87",
X"3f823d0d",
X"04fd3d0d",
X"75528054",
X"80ff7225",
X"8838810b",
X"ff801353",
X"54ffbf12",
X"51709926",
X"8638e012",
X"52b039ff",
X"9f125199",
X"7127a738",
X"d012e013",
X"54517089",
X"26853872",
X"52983972",
X"8f268538",
X"72528f39",
X"71ba2e09",
X"81068538",
X"9a528339",
X"80527380",
X"2e853881",
X"80125271",
X"81ff0683",
X"c0800c85",
X"3d0d0480",
X"3d0d84d8",
X"c0518071",
X"70810553",
X"347084e0",
X"c02e0981",
X"06f03882",
X"3d0d04fe",
X"3d0d0297",
X"053351fe",
X"f43f83c0",
X"800881ff",
X"0683c7d0",
X"08545280",
X"73249b38",
X"83c89008",
X"137283c8",
X"94080753",
X"53717334",
X"83c7d008",
X"810583c7",
X"d00c843d",
X"0d04fa3d",
X"0d82800a",
X"1b558057",
X"883dfc05",
X"54795374",
X"527851ff",
X"bba43f88",
X"3d0d04fe",
X"3d0d83c7",
X"e8085274",
X"51c2883f",
X"83c08008",
X"8c387653",
X"755283c7",
X"e80851c6",
X"3f843d0d",
X"04fe3d0d",
X"83c7e808",
X"53755274",
X"51ffbcc6",
X"3f83c080",
X"088d3877",
X"53765283",
X"c7e80851",
X"ffa03f84",
X"3d0d04fe",
X"3d0d83c7",
X"e80851ff",
X"bbb93f83",
X"c0800881",
X"80802e09",
X"81068838",
X"83c18080",
X"539c3983",
X"c7e80851",
X"ffbb9c3f",
X"83c08008",
X"80d0802e",
X"09810693",
X"3883c1b0",
X"805383c0",
X"80085283",
X"c7e80851",
X"fed43f84",
X"3d0d0480",
X"3d0df9fc",
X"3f83c080",
X"08842981",
X"ddc40570",
X"0883c080",
X"0c51823d",
X"0d04ed3d",
X"0d804480",
X"43804280",
X"4180705a",
X"5bfdcc3f",
X"800b83c7",
X"d00c800b",
X"83c8940c",
X"81dac451",
X"eac13f81",
X"800b83c8",
X"940c81da",
X"c851eab3",
X"3f80d00b",
X"83c7d00c",
X"7830707a",
X"07802570",
X"872b83c8",
X"940c5155",
X"f8ed3f83",
X"c0800852",
X"81dad051",
X"ea8d3f80",
X"f80b83c7",
X"d00c7881",
X"32703070",
X"72078025",
X"70872b83",
X"c8940c51",
X"56569d9e",
X"3f83c080",
X"085281da",
X"e051e9e3",
X"3f81a00b",
X"83c7d00c",
X"78823270",
X"30707207",
X"80257087",
X"2b83c894",
X"0c515656",
X"fec53f83",
X"c0800852",
X"81daf051",
X"e9b93f81",
X"c80b83c7",
X"d00c7883",
X"32703070",
X"72078025",
X"70872b83",
X"c8940c51",
X"5683c7e8",
X"085256ff",
X"b6973f83",
X"c0800852",
X"81daf851",
X"e9893f82",
X"980b83c7",
X"d00c810b",
X"83c7d45b",
X"5883c7d0",
X"0883197a",
X"32703070",
X"72078025",
X"70872b83",
X"c8940c51",
X"578e3d70",
X"55ff1b54",
X"5757579a",
X"e03f7970",
X"84055b08",
X"51ffb5cd",
X"3f745483",
X"c0800853",
X"775281db",
X"8051e8bb",
X"3fa81783",
X"c7d00c81",
X"18587785",
X"2e098106",
X"ffaf3883",
X"b80b83c7",
X"d00c7888",
X"32703070",
X"72078025",
X"70872b83",
X"c8940c51",
X"5656f7b9",
X"3f81db90",
X"5583c080",
X"08802e8f",
X"3883c7e4",
X"0851ffb4",
X"f83f83c0",
X"80085574",
X"5281db98",
X"51e7e83f",
X"84880b83",
X"c7d00c78",
X"89327030",
X"70720780",
X"2570872b",
X"83c8940c",
X"515781db",
X"a45255e7",
X"c63f868d",
X"a051f8b3",
X"3f805291",
X"3d705255",
X"9ea33f83",
X"5274519e",
X"9c3f6355",
X"74839c38",
X"61195978",
X"80258538",
X"74599039",
X"89792585",
X"38885987",
X"39788926",
X"82fb3878",
X"822b5581",
X"d5c41508",
X"04f5d43f",
X"83c08008",
X"61575575",
X"812e0981",
X"06893883",
X"c0800810",
X"55903975",
X"ff2e0981",
X"06883883",
X"c0800881",
X"2c559075",
X"25853890",
X"55883974",
X"80248338",
X"81557451",
X"f5ae3f82",
X"b03999e5",
X"3f83c080",
X"08610555",
X"74802585",
X"38805588",
X"39877525",
X"83388755",
X"74518dc8",
X"3f828e39",
X"f59e3f83",
X"c0800861",
X"05557480",
X"25853880",
X"55883986",
X"75258338",
X"86557451",
X"f5973f81",
X"ec396087",
X"3862802e",
X"81e33883",
X"c39c0883",
X"c3980cad",
X"e50b83c3",
X"a00c83c7",
X"e80851d6",
X"da3ffa8f",
X"3f81c639",
X"60568076",
X"259838ad",
X"840b83c3",
X"a00c83c7",
X"c4157008",
X"5255d6bb",
X"3f740852",
X"92397580",
X"25923883",
X"c7c41508",
X"51ffb2bf",
X"3f8052fc",
X"1951b839",
X"62802e81",
X"8c3883c7",
X"c4157008",
X"83c7d408",
X"720c83c7",
X"d40cfc1a",
X"70535155",
X"8c953f83",
X"c0800856",
X"80518c8b",
X"3f83c080",
X"08527451",
X"88a43f75",
X"52805188",
X"9d3f80d5",
X"39605580",
X"7525b638",
X"83c3a408",
X"83c3980c",
X"ade50b83",
X"c3a00c83",
X"c7e40851",
X"d5c53f83",
X"c7e40851",
X"d2e63f83",
X"c0800881",
X"ff067052",
X"55f3f73f",
X"74802e9d",
X"388155a1",
X"39748025",
X"943883c7",
X"e40851ff",
X"b1b13f80",
X"51f3db3f",
X"84396287",
X"387a802e",
X"f9b73880",
X"557483c0",
X"800c953d",
X"0d04fe3d",
X"0d83c880",
X"5180f4a0",
X"3f83c7f0",
X"5180f498",
X"3ff3f73f",
X"83c08008",
X"802e8638",
X"8051818a",
X"39f3fc3f",
X"83c08008",
X"80fe38f4",
X"9c3f83c0",
X"8008802e",
X"b9388151",
X"f1d93f80",
X"51f3b23f",
X"eecd3f80",
X"0b83c7d0",
X"0cf8cf3f",
X"83c08008",
X"53ff0b83",
X"c7d00cf0",
X"b93f7280",
X"cb3883c7",
X"cc3351f3",
X"8c3f7251",
X"f1a93f80",
X"c039f3c4",
X"3f83c080",
X"08802eb5",
X"388151f1",
X"963f8051",
X"f2ef3fee",
X"8a3fad84",
X"0b83c3a0",
X"0c83c7d4",
X"0851d3e7",
X"3fff0b83",
X"c7d00cef",
X"f53f83c7",
X"d4085280",
X"51868b3f",
X"8151f4b6",
X"3f843d0d",
X"04fb3d0d",
X"805283c8",
X"805180e3",
X"a73f8152",
X"83c7f051",
X"80e39d3f",
X"800b83c7",
X"cc349080",
X"80528684",
X"808051ff",
X"b3c63f83",
X"c0800881",
X"973889dc",
X"3f81dfe4",
X"51ffb885",
X"3f83c080",
X"08559c80",
X"0a5480c0",
X"805381db",
X"ac5283c0",
X"800851f6",
X"883f83c7",
X"e8085381",
X"dbbc5274",
X"51ffb2ce",
X"3f83c080",
X"088438f6",
X"963f83c7",
X"ec085381",
X"dbc85274",
X"51ffb2b6",
X"3f83c080",
X"08b63887",
X"3dfc0554",
X"84808053",
X"86a88080",
X"5283c7ec",
X"0851ffb0",
X"c13f83c0",
X"80089338",
X"75848080",
X"2e098106",
X"8938810b",
X"83c7cc34",
X"8739800b",
X"83c7cc34",
X"83c7cc33",
X"51f1823f",
X"8151f2ee",
X"3f938d3f",
X"8151f2e6",
X"3f8151fc",
X"fd3ffa39",
X"83c08c08",
X"0283c08c",
X"0cfb3d0d",
X"0281dbd4",
X"0b83c39c",
X"0c81dbd8",
X"0b83c394",
X"0c81dbdc",
X"0b83c3a4",
X"0c83c08c",
X"08fc050c",
X"800b83c7",
X"d40b83c0",
X"8c08f805",
X"0c83c08c",
X"08f4050c",
X"ffb0d13f",
X"83c08008",
X"8605fc06",
X"83c08c08",
X"f0050c02",
X"83c08c08",
X"f0050831",
X"0d833d70",
X"83c08c08",
X"f8050870",
X"840583c0",
X"8c08f805",
X"0c0c51ff",
X"ad993f83",
X"c08c08f4",
X"05088105",
X"83c08c08",
X"f4050c83",
X"c08c08f4",
X"0508872e",
X"098106ff",
X"ab388694",
X"808051ea",
X"af3fff0b",
X"83c7d00c",
X"800b83c8",
X"940c84d8",
X"c00b83c8",
X"900c8151",
X"edd93f81",
X"51edfe3f",
X"8051edf9",
X"3f8151ee",
X"9f3f8251",
X"eec73f80",
X"51eeef3f",
X"8051ef99",
X"3f80d0af",
X"528051df",
X"933ffccd",
X"3f83c08c",
X"08fc0508",
X"0d800b83",
X"c0800c87",
X"3d0d83c0",
X"8c0c0480",
X"3d0d81ff",
X"51800b83",
X"c8a41234",
X"ff115170",
X"f438823d",
X"0d04ff3d",
X"0d737033",
X"53518111",
X"33713471",
X"81123483",
X"3d0d04fb",
X"3d0d7779",
X"56568070",
X"71555552",
X"717525ac",
X"38721670",
X"33701470",
X"81ff0655",
X"51515171",
X"74278938",
X"81127081",
X"ff065351",
X"71811470",
X"83ffff06",
X"55525474",
X"7324d638",
X"7183c080",
X"0c873d0d",
X"04fb3d0d",
X"7756d6dd",
X"3f83c080",
X"08802ef6",
X"3883cac0",
X"08860570",
X"81ff0652",
X"53d4df3f",
X"810b9088",
X"d4349088",
X"d4337081",
X"ff065153",
X"728b38f9",
X"dd3f8351",
X"eecd3fea",
X"39805574",
X"1675822b",
X"54549088",
X"c0133374",
X"34811555",
X"74852e09",
X"8106e838",
X"810b9088",
X"d4347533",
X"83c8a434",
X"81163383",
X"c8a53482",
X"163383c8",
X"a6348316",
X"3383c8a7",
X"34845283",
X"c8a451fe",
X"ba3f83c0",
X"800881ff",
X"06841733",
X"57537276",
X"2e098106",
X"8c38d586",
X"3f83c080",
X"08802e9c",
X"3883cac0",
X"08a82e09",
X"81068b38",
X"83cad808",
X"83cac00c",
X"8739a80b",
X"83cac00c",
X"80e451ed",
X"c63f873d",
X"0d04f43d",
X"0d7e6059",
X"55805d80",
X"75822b71",
X"83cac412",
X"0c83cadc",
X"175b5b57",
X"76793477",
X"772e83b7",
X"38765277",
X"51ffabe2",
X"3f8e3dfc",
X"05549053",
X"83caac52",
X"7751ffab",
X"9d3f7c56",
X"75902e09",
X"81068393",
X"3883caac",
X"51fd933f",
X"83caae51",
X"fd8c3f83",
X"cab051fd",
X"853f7683",
X"cabc0c77",
X"51ffa8e9",
X"3f81d9d4",
X"5283c080",
X"0851cb82",
X"3f83c080",
X"08812e09",
X"810680d4",
X"387683ca",
X"d40c820b",
X"83caac34",
X"ff960b83",
X"caad3477",
X"51ffabaf",
X"3f83c080",
X"085583c0",
X"80087725",
X"883883c0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83caae34",
X"7483caaf",
X"347683ca",
X"b034ff80",
X"0b83cab1",
X"34819039",
X"83caac33",
X"83caad33",
X"71882b07",
X"565b7483",
X"ffff2e09",
X"810680e8",
X"38fe800b",
X"83cad40c",
X"810b83ca",
X"bc0cff0b",
X"83caac34",
X"ff0b83ca",
X"ad347751",
X"ffaabc3f",
X"83c08008",
X"83cae00c",
X"83c08008",
X"5583c080",
X"08802588",
X"3883c080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"caae3474",
X"83caaf34",
X"7683cab0",
X"34ff800b",
X"83cab134",
X"810b83ca",
X"bb34a539",
X"7485962e",
X"09810680",
X"fe387583",
X"cad40c77",
X"51ffa9f0",
X"3f83cabb",
X"3383c080",
X"08075574",
X"83cabb34",
X"83cabb33",
X"81065574",
X"802e8338",
X"845783ca",
X"b03383ca",
X"b1337188",
X"2b07565c",
X"7481802e",
X"098106a1",
X"3883caae",
X"3383caaf",
X"3371882b",
X"07565bad",
X"80752787",
X"38768207",
X"579c3976",
X"81075796",
X"39748280",
X"2e098106",
X"87387683",
X"07578739",
X"7481ff26",
X"8a387783",
X"cac41b0c",
X"7679348e",
X"3d0d0480",
X"3d0d7284",
X"2983cac4",
X"05700883",
X"c0800c51",
X"823d0d04",
X"803d0d72",
X"7083c89c",
X"0c708429",
X"81df9805",
X"700883ca",
X"d80c5151",
X"823d0d04",
X"fe3d0d81",
X"51de3f80",
X"0b83caa8",
X"0c800b83",
X"caa40cff",
X"0b83c8a0",
X"0ca80b83",
X"cac00cae",
X"51cf873f",
X"800b83ca",
X"c4545280",
X"73708405",
X"550c8112",
X"5271842e",
X"098106ef",
X"38843d0d",
X"04fe3d0d",
X"74028405",
X"96052253",
X"5371802e",
X"96387270",
X"81055433",
X"51cf923f",
X"ff127083",
X"ffff0651",
X"52e73984",
X"3d0d04fe",
X"3d0d0292",
X"05225382",
X"ac51e8bb",
X"3f80c351",
X"ceef3f81",
X"9651e8af",
X"3f725283",
X"c8a451ff",
X"b43f7252",
X"83c8a451",
X"f8d13f83",
X"c0800881",
X"ff0651ce",
X"cc3f843d",
X"0d04ffb1",
X"3d0d80d1",
X"3df80551",
X"f8fb3f83",
X"caa80881",
X"0583caa8",
X"0c80cf3d",
X"33cf1170",
X"81ff0651",
X"56567483",
X"2688e638",
X"758f06ff",
X"05567583",
X"c8a0082e",
X"9b387583",
X"26963875",
X"83c8a00c",
X"75842983",
X"cac40570",
X"08535575",
X"51f9fb3f",
X"80762488",
X"c2387584",
X"2983cac4",
X"05557408",
X"802e88b3",
X"3883c8a0",
X"08842983",
X"cac40570",
X"08028805",
X"82b90533",
X"525b5574",
X"80d22e84",
X"b0387480",
X"d2249038",
X"74bf2e9c",
X"387480d0",
X"2e81d538",
X"87f23974",
X"80d32e80",
X"d3387480",
X"d72e81c4",
X"3887e139",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"055656cd",
X"c83f80c1",
X"51cd823f",
X"f6cd3f83",
X"cadb3383",
X"c8a43481",
X"5283c8a4",
X"51cea33f",
X"8151fde7",
X"3f748b38",
X"83cad808",
X"83cac00c",
X"8739a80b",
X"83cac00c",
X"cd933f80",
X"c151cccd",
X"3ff6983f",
X"900b83ca",
X"bb338106",
X"56567480",
X"2e833898",
X"5683cab0",
X"3383cab1",
X"3371882b",
X"07565974",
X"81802e09",
X"81069c38",
X"83caae33",
X"83caaf33",
X"71882b07",
X"5657ad80",
X"75278c38",
X"75818007",
X"56853975",
X"a0075675",
X"83c8a434",
X"ff0b83c8",
X"a534e00b",
X"83c8a634",
X"800b83c8",
X"a7348452",
X"83c8a451",
X"cd983f84",
X"51869b39",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"055659cc",
X"883f7951",
X"ffa49d3f",
X"83c08008",
X"802e8a38",
X"80ce51cb",
X"b43f85f1",
X"3980c151",
X"cbab3fcc",
X"a03fcad5",
X"3f83cad4",
X"08588375",
X"259b3883",
X"cab03383",
X"cab13371",
X"882b07fc",
X"1771297a",
X"05838005",
X"5a51578d",
X"39748180",
X"2918ff80",
X"05588180",
X"57805676",
X"762e9238",
X"cb873f83",
X"c0800883",
X"c8a41734",
X"811656eb",
X"39caf63f",
X"83c08008",
X"81ff0677",
X"5383c8a4",
X"5256f4c3",
X"3f83c080",
X"0881ff06",
X"5575752e",
X"09810681",
X"95389451",
X"e3f93fca",
X"f03f80c1",
X"51caaa3f",
X"cb9f3f77",
X"527951ff",
X"a2b03f80",
X"5e80d13d",
X"fdf40554",
X"765383c8",
X"a4527951",
X"ffa0bd3f",
X"0282b905",
X"33558159",
X"7480d72e",
X"09810680",
X"c5387752",
X"7951ffa2",
X"813f80d1",
X"3dfdf005",
X"5476538f",
X"3d70537a",
X"5258ffa1",
X"b93f8056",
X"76762ea2",
X"38751883",
X"c8a41733",
X"71337072",
X"32703070",
X"80257030",
X"7f06811d",
X"5d5f5151",
X"51525b55",
X"db3982ac",
X"51e2f43f",
X"78802e86",
X"3880c351",
X"843980ce",
X"51c99e3f",
X"ca933fc8",
X"c83f83d8",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055955",
X"80705d59",
X"80e451e2",
X"be3fc9b5",
X"3f80c151",
X"c8ef3f83",
X"cabc0879",
X"2e82d638",
X"83cae008",
X"80fc0555",
X"80fd5274",
X"5185c13f",
X"83c08008",
X"5b778224",
X"b238ff18",
X"70872b83",
X"ffff8006",
X"81dde405",
X"83c8a459",
X"57558180",
X"55757081",
X"05573377",
X"70810559",
X"34ff1570",
X"81ff0651",
X"5574ea38",
X"82853977",
X"82e82e81",
X"a3387782",
X"e92e0981",
X"0681aa38",
X"78587787",
X"32703070",
X"72078025",
X"7a8a3270",
X"30707207",
X"80257307",
X"53545a51",
X"57557580",
X"2e973878",
X"78269238",
X"a00b83c8",
X"a41a3481",
X"197081ff",
X"065a55eb",
X"39811870",
X"81ff0659",
X"558a7827",
X"ffbc388f",
X"5883c89f",
X"183383c8",
X"a41934ff",
X"187081ff",
X"06595577",
X"8426ea38",
X"9058800b",
X"83c8a419",
X"34811870",
X"81ff0670",
X"982b5259",
X"55748025",
X"e93880c6",
X"557a858f",
X"24843880",
X"c2557483",
X"c8a43480",
X"f10b83c8",
X"a734810b",
X"83c8a834",
X"7a83c8a5",
X"347a882c",
X"557483c8",
X"a63480cb",
X"3982f078",
X"2580c438",
X"7780fd29",
X"fd97d305",
X"527951ff",
X"9edc3f80",
X"d13dfdec",
X"055480fd",
X"5383c8a4",
X"527951ff",
X"9e943f7b",
X"81195956",
X"7580fc24",
X"83387858",
X"77882c55",
X"7483c9a1",
X"347783c9",
X"a2347583",
X"c9a33481",
X"805980cc",
X"3983cad4",
X"08578378",
X"259b3883",
X"cab03383",
X"cab13371",
X"882b07fc",
X"1a712979",
X"05838005",
X"5951598d",
X"39778180",
X"2917ff80",
X"05578180",
X"59765279",
X"51ff9dea",
X"3f80d13d",
X"fdec0554",
X"785383c8",
X"a4527951",
X"ff9da33f",
X"7851f6bf",
X"3fc6b63f",
X"c4eb3f8b",
X"3983caa4",
X"08810583",
X"caa40c80",
X"d13d0d04",
X"f6e03ffc",
X"39fc3d0d",
X"76787184",
X"2983cac4",
X"05700851",
X"53535370",
X"9e3880ce",
X"723480cf",
X"0b811334",
X"80ce0b82",
X"133480c5",
X"0b831334",
X"70841334",
X"80e73983",
X"cadc1333",
X"5480d272",
X"3473822a",
X"70810651",
X"5180cf53",
X"70843880",
X"d7537281",
X"1334a00b",
X"82133473",
X"83065170",
X"812e9e38",
X"70812488",
X"3870802e",
X"8f389f39",
X"70822e92",
X"3870832e",
X"92389339",
X"80d8558e",
X"3980d355",
X"893980cd",
X"55843980",
X"c4557483",
X"133480c4",
X"0b841334",
X"800b8513",
X"34863d0d",
X"0483c89c",
X"0883c080",
X"0c04803d",
X"0d83c89c",
X"08842981",
X"dfb80570",
X"0883c080",
X"0c51823d",
X"0d04fc3d",
X"0d767853",
X"54815380",
X"55873971",
X"10731054",
X"52737226",
X"5172802e",
X"a7387080",
X"2e863871",
X"8025e838",
X"72802e98",
X"38717426",
X"89387372",
X"31757407",
X"56547281",
X"2a72812a",
X"5353e539",
X"73517883",
X"38745170",
X"83c0800c",
X"863d0d04",
X"fe3d0d80",
X"53755274",
X"51ffa33f",
X"843d0d04",
X"fe3d0d81",
X"53755274",
X"51ff933f",
X"843d0d04",
X"fb3d0d77",
X"79555580",
X"56747625",
X"86387430",
X"55815673",
X"80258838",
X"73307681",
X"32575480",
X"53735274",
X"51fee73f",
X"83c08008",
X"5475802e",
X"873883c0",
X"80083054",
X"7383c080",
X"0c873d0d",
X"04fa3d0d",
X"787a5755",
X"80577477",
X"25863874",
X"30558157",
X"759f2c54",
X"81537574",
X"32743152",
X"7451feaa",
X"3f83c080",
X"08547680",
X"2e873883",
X"c0800830",
X"547383c0",
X"800c883d",
X"0d04fc3d",
X"0d765580",
X"750c800b",
X"84160c80",
X"0b88160c",
X"800b8c16",
X"0c83c880",
X"5180dad4",
X"3f83c7f0",
X"5180dacc",
X"3f87a680",
X"337081ff",
X"065152da",
X"f53f7181",
X"2a813272",
X"81327181",
X"06718106",
X"3184180c",
X"54547183",
X"2a813272",
X"822a8132",
X"71810671",
X"81063177",
X"0c535387",
X"a0903370",
X"09810688",
X"170c5283",
X"c0800880",
X"2e80c238",
X"83c08008",
X"812a7081",
X"0683c080",
X"08810631",
X"84170c52",
X"83c08008",
X"832a83c0",
X"8008822a",
X"71810671",
X"81063177",
X"0c535383",
X"c0800884",
X"2a810688",
X"160c83c0",
X"8008852a",
X"81068c16",
X"0c863d0d",
X"04fe3d0d",
X"74765452",
X"7151febe",
X"3f72812e",
X"a2388173",
X"268d3872",
X"822ea838",
X"72832e9c",
X"38e63971",
X"08e23884",
X"1208dd38",
X"881208d8",
X"38a53988",
X"1208812e",
X"9e389139",
X"88120881",
X"2e953871",
X"08913884",
X"12088c38",
X"8c120881",
X"2e098106",
X"ffb23884",
X"3d0d04fb",
X"3d0d7802",
X"84059f05",
X"33555680",
X"0b81d7d8",
X"56538173",
X"2b740652",
X"71802e83",
X"38815274",
X"70820556",
X"22707390",
X"2b079080",
X"9c0c5181",
X"13537288",
X"2e098106",
X"d9388053",
X"83cae813",
X"33517081",
X"ff2eb238",
X"701081d5",
X"f8057022",
X"55518073",
X"17703370",
X"1081d5f8",
X"05702251",
X"51515252",
X"73712e91",
X"38811252",
X"71862e09",
X"8106f138",
X"7390809c",
X"0c811353",
X"72862e09",
X"8106ffb8",
X"38805372",
X"16703351",
X"517081ff",
X"2e943870",
X"1081d5f8",
X"05702270",
X"84808007",
X"90809c0c",
X"51518113",
X"5372862e",
X"098106d7",
X"38805372",
X"16517033",
X"83cae814",
X"34811353",
X"72862e09",
X"8106ec38",
X"873d0d04",
X"04ff3d0d",
X"74028405",
X"8f053352",
X"52708838",
X"71908094",
X"0c8e3970",
X"812e0981",
X"06863871",
X"9080980c",
X"833d0d04",
X"fb3d0d02",
X"9f053379",
X"982b7098",
X"2c7c982b",
X"70982c83",
X"cb841570",
X"3370982b",
X"70982c51",
X"585c5a51",
X"55515454",
X"70732e09",
X"81069438",
X"83cae414",
X"3370982b",
X"70982c51",
X"52567072",
X"2eb13872",
X"75347183",
X"cae41534",
X"83cae533",
X"83cb8533",
X"71982b71",
X"902b0783",
X"cae43370",
X"882b7207",
X"83cb8433",
X"71079080",
X"b80c5259",
X"53545287",
X"3d0d04fe",
X"3d0d7481",
X"11337133",
X"71882b07",
X"83c0800c",
X"5351843d",
X"0d0483ca",
X"f03383c0",
X"800c04f5",
X"3d0d02bb",
X"05330284",
X"05bf0533",
X"02880580",
X"c3053302",
X"8c0580c6",
X"0522665c",
X"5a5e5c56",
X"7a557b54",
X"8953a152",
X"7d5180d0",
X"c03f83c0",
X"800881ff",
X"0683c080",
X"0c8d3d0d",
X"0483c08c",
X"080283c0",
X"8c0cf53d",
X"0d83c08c",
X"08880508",
X"83c08c08",
X"8f053383",
X"c08c0892",
X"0522028c",
X"05739005",
X"83c08c08",
X"e8050c83",
X"c08c08f8",
X"050c83c0",
X"8c08f005",
X"0c83c08c",
X"08ec050c",
X"83c08c08",
X"f4050c80",
X"0b83c08c",
X"08f00508",
X"83c08c08",
X"e0050c83",
X"c08c08fc",
X"050c83c0",
X"8c08f005",
X"0889278a",
X"38890b83",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08860587",
X"fffc0683",
X"c08c08e0",
X"050c0283",
X"c08c08e0",
X"0508310d",
X"853d7055",
X"83c08c08",
X"ec050854",
X"83c08c08",
X"f0050853",
X"83c08c08",
X"f4050852",
X"83c08c08",
X"e4050c80",
X"d9f23f83",
X"c0800881",
X"ff0683c0",
X"8c08e405",
X"0883c08c",
X"08ec050c",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508802e",
X"8c3883c0",
X"8c08f805",
X"080d89c8",
X"3983c08c",
X"08f00508",
X"802e89a6",
X"3883c08c",
X"08ec0508",
X"81053383",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08842ea9",
X"38840b83",
X"c08c08e0",
X"05082588",
X"c73883c0",
X"8c08e005",
X"08852e85",
X"9b3883c0",
X"8c08e005",
X"08a12e87",
X"ad3888ac",
X"39800b83",
X"c08c08ec",
X"05088505",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"fc050c83",
X"c08c08e0",
X"0508832e",
X"09810688",
X"833883c0",
X"8c08e805",
X"08810533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"05088126",
X"87e63881",
X"0b83c08c",
X"08e00508",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08fc05",
X"0c83c08c",
X"08ec0508",
X"82053383",
X"c08c08e0",
X"05088705",
X"3483c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c800b83",
X"c08c08e0",
X"05088b05",
X"3483c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08f405",
X"0c800b83",
X"c08c08e0",
X"05088c05",
X"3483c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c800b83",
X"c08c08e0",
X"05088d05",
X"3483c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08f405",
X"0c800b83",
X"c08c08e0",
X"05088e05",
X"2383c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c800b83",
X"c08c08e0",
X"05088a05",
X"3483c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080570",
X"940508fc",
X"ffff0671",
X"94050c83",
X"c08c08e0",
X"050c83c0",
X"8c08ec05",
X"08860533",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c83c0",
X"8c08e005",
X"0883c08c",
X"08fc0508",
X"2e098106",
X"b63883c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c83c0",
X"8c08fc05",
X"0883c08c",
X"08e00508",
X"8b053483",
X"c08c08ec",
X"05088705",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e0050881",
X"2e8f3883",
X"c08c08e0",
X"0508822e",
X"b738848c",
X"3983c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08f405",
X"0c820b83",
X"c08c08e0",
X"05088a05",
X"3483d939",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"83c08c08",
X"fc050883",
X"c08c08e0",
X"05088a05",
X"3483a139",
X"83c08c08",
X"fc050880",
X"2e839538",
X"83c08c08",
X"ec050883",
X"05338306",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508832e",
X"09810682",
X"f33883c0",
X"8c08ec05",
X"08820533",
X"70982b83",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08e00508",
X"802582cc",
X"3883c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08f405",
X"0c83c08c",
X"08ec0508",
X"86053383",
X"c08c08e0",
X"050880d6",
X"053483c0",
X"8c08e005",
X"08840583",
X"c08c08ec",
X"05088205",
X"338f0683",
X"c08c08e4",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08e40508",
X"83c08c08",
X"e0050834",
X"83c08c08",
X"ec050884",
X"053383c0",
X"8c08e005",
X"08810534",
X"800b83c0",
X"8c08e005",
X"08820534",
X"83c08c08",
X"e0050808",
X"ff83ff06",
X"82800783",
X"c08c08e0",
X"05080c83",
X"c08c08e8",
X"05088105",
X"33810583",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"0883c08c",
X"08e80508",
X"81053481",
X"833983c0",
X"8c08fc05",
X"08802e80",
X"f73883c0",
X"8c08ec05",
X"08860533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508a22e",
X"09810680",
X"d73883c0",
X"8c08ec05",
X"08880533",
X"83c08c08",
X"ec050887",
X"05337182",
X"80290583",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"5283c08c",
X"08e4050c",
X"83c08c08",
X"f4050c83",
X"c08c08e4",
X"050883c0",
X"8c08e005",
X"08880523",
X"83c08c08",
X"ec050833",
X"83c08c08",
X"f0050871",
X"317083ff",
X"ff0683c0",
X"8c08f005",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"ec050805",
X"83c08c08",
X"ec050cf6",
X"d03983c0",
X"8c08f805",
X"080d83c0",
X"8c08f005",
X"0883c08c",
X"08e0050c",
X"83c08c08",
X"f805080d",
X"83c08c08",
X"e0050883",
X"c0800c8d",
X"3d0d83c0",
X"8c0c0483",
X"c08c0802",
X"83c08c0c",
X"e63d0d83",
X"c08c0888",
X"05080284",
X"0583c08c",
X"08e8050c",
X"83c08c08",
X"d4050c80",
X"0b83cb8c",
X"3483c08c",
X"08d40508",
X"900583c0",
X"8c08c005",
X"0c800b83",
X"c08c08c0",
X"05083480",
X"0b83c08c",
X"08c00508",
X"81053480",
X"0b83c08c",
X"08c4050c",
X"83c08c08",
X"c4050880",
X"d82983c0",
X"8c08c005",
X"080583c0",
X"8c08ffb4",
X"050c800b",
X"83c08c08",
X"ffb40508",
X"80d8050c",
X"83c08c08",
X"ffb40508",
X"840583c0",
X"8c08ffb4",
X"050c83c0",
X"8c08c405",
X"0883c08c",
X"08ffb405",
X"0834880b",
X"83c08c08",
X"ffb40508",
X"81053480",
X"0b83c08c",
X"08ffb405",
X"08820534",
X"83c08c08",
X"ffb40508",
X"08ffa1ff",
X"06a08007",
X"83c08c08",
X"ffb40508",
X"0c83c08c",
X"08c40508",
X"81057081",
X"ff0683c0",
X"8c08c405",
X"0c83c08c",
X"08ffb405",
X"0c810b83",
X"c08c08c4",
X"050827fe",
X"db3883c0",
X"8c08ec05",
X"705483c0",
X"8c08c805",
X"0c925283",
X"c08c08d4",
X"05085180",
X"cd993f83",
X"c0800881",
X"ff067083",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b805088d",
X"ea3883c0",
X"8c08f405",
X"51f18c3f",
X"83c08008",
X"83ffff06",
X"83c08c08",
X"f6055283",
X"c08c08e4",
X"050cf0f3",
X"3f83c080",
X"0883ffff",
X"0683c08c",
X"08fd0533",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"c4050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08e0",
X"050c83c0",
X"8c08c405",
X"0883c08c",
X"08ffbc05",
X"082780fe",
X"3883c08c",
X"08c80508",
X"5483c08c",
X"08c40508",
X"53895283",
X"c08c08d4",
X"05085180",
X"cc9e3f83",
X"c0800881",
X"ff0683c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"050880f2",
X"3883c08c",
X"08ee0551",
X"eff13f83",
X"c0800883",
X"ffff0653",
X"83c08c08",
X"c4050852",
X"83c08c08",
X"d4050851",
X"f0b33f83",
X"c08c08c4",
X"05088105",
X"7081ff06",
X"83c08c08",
X"c4050c83",
X"c08c08ff",
X"b4050cfe",
X"f13983c0",
X"8c08c005",
X"08810533",
X"83c08c08",
X"ffb4050c",
X"81db0b83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"b4050880",
X"2e8be038",
X"943983c0",
X"8c08ffb8",
X"050883c0",
X"8c08ffbc",
X"050c8bcb",
X"3983c08c",
X"08f10533",
X"5283c08c",
X"08d40508",
X"5180cb9c",
X"3f800b83",
X"c08c08c0",
X"05088105",
X"3383c08c",
X"08ffb405",
X"0c83c08c",
X"08c4050c",
X"83c08c08",
X"c4050883",
X"c08c08ff",
X"b4050827",
X"89e63883",
X"c08c08c4",
X"050880d8",
X"297083c0",
X"8c08c005",
X"08057088",
X"05708305",
X"3383c08c",
X"08cc050c",
X"83c08c08",
X"c8050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08d8",
X"050c83c0",
X"8c08cc05",
X"0887a638",
X"83c08c08",
X"c8050822",
X"02840571",
X"860587ff",
X"fc0683c0",
X"8c08ffb4",
X"050c83c0",
X"8c08dc05",
X"0c83c08c",
X"08ffb805",
X"0c0283c0",
X"8c08ffb4",
X"0508310d",
X"893d7059",
X"83c08c08",
X"ffb80508",
X"5883c08c",
X"08ffbc05",
X"08870533",
X"5783c08c",
X"08ffb405",
X"0ca25583",
X"c08c08cc",
X"05085486",
X"53818152",
X"83c08c08",
X"d4050851",
X"be933f83",
X"c0800881",
X"ff0683c0",
X"8c08d005",
X"0c83c08c",
X"08d00508",
X"81c13883",
X"c08c08ff",
X"bc050896",
X"055383c0",
X"8c08ffb8",
X"05085283",
X"c08c08ff",
X"b4050851",
X"a1c63f83",
X"c0800881",
X"ff0683c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb4",
X"0508802e",
X"81853883",
X"c08c08ff",
X"bc050894",
X"0583c08c",
X"08ffbc05",
X"08960533",
X"70862a83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08cc",
X"050c83c0",
X"8c08ffb4",
X"0508832e",
X"09810680",
X"c63883c0",
X"8c08ffb4",
X"050883c0",
X"8c08c805",
X"08820534",
X"83caf033",
X"70810583",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b4050883",
X"caf03483",
X"c08c08ff",
X"b8050883",
X"c08c08cc",
X"05083483",
X"c08c08dc",
X"05080d83",
X"c08c08d0",
X"050881ff",
X"0683c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"08fbff38",
X"83c08c08",
X"d8050883",
X"c08c08c0",
X"05080588",
X"05708205",
X"335183c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb4",
X"0508832e",
X"09810680",
X"e33883c0",
X"8c08ffb8",
X"050883c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb4",
X"05088105",
X"7081ff06",
X"5183c08c",
X"08ffb405",
X"0c810b83",
X"c08c08ff",
X"b4050827",
X"dd38800b",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb40508",
X"81057081",
X"ff065183",
X"c08c08ff",
X"b4050c97",
X"0b83c08c",
X"08ffb405",
X"0827dd38",
X"83c08c08",
X"e4050880",
X"f9327030",
X"70802551",
X"5183c08c",
X"08ffb405",
X"0c83c08c",
X"08e00508",
X"912e0981",
X"0680f938",
X"83c08c08",
X"ffb40508",
X"802e80ec",
X"3883c08c",
X"08c40508",
X"80e23885",
X"0b83c08c",
X"08c00508",
X"a60534a0",
X"0b83c08c",
X"08c00508",
X"a7053485",
X"0b83c08c",
X"08c00508",
X"a8053480",
X"c00b83c0",
X"8c08c005",
X"08a90534",
X"860b83c0",
X"8c08c005",
X"08aa0534",
X"900b83c0",
X"8c08c005",
X"08ab0534",
X"860b83c0",
X"8c08c005",
X"08ac0534",
X"a00b83c0",
X"8c08c005",
X"08ad0534",
X"83c08c08",
X"e4050889",
X"d8327030",
X"70802551",
X"5183c08c",
X"08ffb405",
X"0c83c08c",
X"08e00508",
X"83edec2e",
X"09810680",
X"f6388170",
X"83c08c08",
X"ffb40508",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb405",
X"08802e80",
X"ce3883c0",
X"8c08c405",
X"0880c438",
X"840b83c0",
X"8c08c005",
X"08aa0534",
X"80c00b83",
X"c08c08c0",
X"0508ab05",
X"34840b83",
X"c08c08c0",
X"0508ac05",
X"34900b83",
X"c08c08c0",
X"0508ad05",
X"3483c08c",
X"08ffb805",
X"0883c08c",
X"08c00508",
X"8c053483",
X"c08c08e4",
X"050880f9",
X"32703070",
X"80255151",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"e0050886",
X"2e098106",
X"80c33881",
X"7083c08c",
X"08ffb405",
X"080683c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb4",
X"0508802e",
X"9c3883c0",
X"8c08c405",
X"08933883",
X"c08c08ff",
X"b8050883",
X"c08c08c0",
X"05088d05",
X"3483c08c",
X"08c40508",
X"80d82983",
X"c08c08c0",
X"05080570",
X"84057083",
X"053383c0",
X"8c08ffb4",
X"050c83c0",
X"8c08c805",
X"0c83c08c",
X"08ffbc05",
X"0c805880",
X"5783c08c",
X"08ffb405",
X"08568055",
X"80548a53",
X"a15283c0",
X"8c08d405",
X"0851b78d",
X"3f83c080",
X"0881ff06",
X"7030709f",
X"2a5183c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"0508a02e",
X"8c3883c0",
X"8c08ffb4",
X"0508f6c2",
X"3883c08c",
X"08ffbc05",
X"088b0533",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb40508",
X"802eb338",
X"83c08c08",
X"c8050883",
X"053383c0",
X"8c08ffb4",
X"050c8058",
X"805783c0",
X"8c08ffb4",
X"05085680",
X"5580548b",
X"53a15283",
X"c08c08d4",
X"050851b6",
X"883f83c0",
X"8c08c405",
X"08810570",
X"81ff0683",
X"c08c08c0",
X"05088105",
X"335283c0",
X"8c08c405",
X"0c83c08c",
X"08ffb405",
X"0cf68939",
X"800b83c0",
X"8c08c405",
X"0c83c08c",
X"08c40508",
X"80d82983",
X"c08c08d4",
X"05080570",
X"9a053383",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b4050882",
X"2e098106",
X"a93883cb",
X"8c568155",
X"805483c0",
X"8c08ffb4",
X"05085383",
X"c08c08ff",
X"b8050897",
X"05335283",
X"c08c08d4",
X"050851e4",
X"8a3f83c0",
X"8c08c405",
X"08810570",
X"81ff0683",
X"c08c08c4",
X"050c83c0",
X"8c08ffb4",
X"050c810b",
X"83c08c08",
X"c4050827",
X"fefb3881",
X"0b83c08c",
X"08c00508",
X"34800b83",
X"c08c08ff",
X"bc050c83",
X"c08c08e8",
X"05080d83",
X"c08c08ff",
X"bc050883",
X"c0800c9c",
X"3d0d83c0",
X"8c0c04f5",
X"3d0d901e",
X"57800b81",
X"18335459",
X"78732781",
X"9d387880",
X"d829178a",
X"11335454",
X"72832e09",
X"810680f8",
X"38941433",
X"5ba98c3f",
X"83c08008",
X"5a805675",
X"81c4291a",
X"87113354",
X"5472802e",
X"80c03873",
X"0881d5ec",
X"2e098106",
X"b5388074",
X"59557480",
X"d829189a",
X"11335454",
X"72832e09",
X"81069238",
X"a4147033",
X"54547a73",
X"278738ff",
X"13537274",
X"34811570",
X"81ff0656",
X"53817527",
X"d1388116",
X"7081ff06",
X"57538f76",
X"27ffa438",
X"83caf033",
X"ff055372",
X"83caf034",
X"81197081",
X"ff068119",
X"335e5a53",
X"7b7926fe",
X"e538800b",
X"83c0800c",
X"8d3d0d04",
X"83c08c08",
X"0283c08c",
X"0ce63d0d",
X"83c08c08",
X"88050802",
X"84057190",
X"05703370",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"c8050c83",
X"c08c08dc",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08ffa405",
X"08802e94",
X"b538800b",
X"83c08c08",
X"c8050881",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08d405",
X"0c83c08c",
X"08d40508",
X"83c08c08",
X"ffa40508",
X"2593fd38",
X"83c08c08",
X"d4050880",
X"d82983c0",
X"8c08c805",
X"08058405",
X"70860533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffa40508",
X"802e9389",
X"38a6b23f",
X"83c08c08",
X"ffb80508",
X"80d40508",
X"83c08008",
X"2692f238",
X"0283c08c",
X"08ffb805",
X"08810533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"d8050c83",
X"c08c08ff",
X"a4050883",
X"c08c08fc",
X"052383c0",
X"8c08ffa4",
X"05088605",
X"83fc0683",
X"c08c08ff",
X"a4050c02",
X"83c08c08",
X"ffa40508",
X"310d853d",
X"705583c0",
X"8c08fc05",
X"5483c08c",
X"08ffb805",
X"085383c0",
X"8c08e005",
X"085283c0",
X"8c08c005",
X"0cae8a3f",
X"83c08008",
X"81ff0683",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050891",
X"bb3883c0",
X"8c08ffb8",
X"05088705",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e80",
X"d53883c0",
X"8c08ffb8",
X"05088605",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08822e09",
X"8106b338",
X"83c08c08",
X"fc052283",
X"c08c08ff",
X"a4050c87",
X"0b83c08c",
X"08ffa405",
X"08279738",
X"83c08c08",
X"c0050882",
X"055283c0",
X"8c08c005",
X"083351db",
X"a63f83c0",
X"8c08ffb8",
X"05088605",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08832e09",
X"810690a4",
X"3883c08c",
X"08ffb805",
X"08920570",
X"82053383",
X"c08c08fc",
X"052283c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08c405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffa805",
X"08268fe4",
X"38800b83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffb00508",
X"1083c08c",
X"0805f805",
X"83c08c08",
X"ffb00508",
X"842983c0",
X"8c08ffb0",
X"05081005",
X"83c08c08",
X"c4050805",
X"70840570",
X"3383c08c",
X"08c00508",
X"05703383",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"b4050883",
X"c08c08ff",
X"bc050823",
X"83c08c08",
X"ffa80508",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050890",
X"2e098106",
X"be3883c0",
X"8c08ffa8",
X"05083383",
X"c08c08c0",
X"05080581",
X"05703370",
X"82802983",
X"c08c08ff",
X"b4050805",
X"515183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffbc",
X"05082383",
X"c08c08ff",
X"ac050886",
X"052283c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa8",
X"0508a238",
X"83c08c08",
X"ffac0508",
X"88052283",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050881",
X"ff2e80e5",
X"3883c08c",
X"08ffbc05",
X"08227083",
X"c08c08ff",
X"a8050831",
X"70828029",
X"713183c0",
X"8c08ffac",
X"05088805",
X"227083c0",
X"8c08ffa8",
X"05083170",
X"73355383",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"ac050c51",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffbc0508",
X"2383c08c",
X"08ffb005",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a4050c81",
X"0b83c08c",
X"08ffb005",
X"0827fce0",
X"3883c08c",
X"08f80522",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"bf269138",
X"83c08c08",
X"e4050882",
X"0783c08c",
X"08e4050c",
X"81c00b83",
X"c08c08ff",
X"a4050827",
X"913883c0",
X"8c08e405",
X"08810783",
X"c08c08e4",
X"050c83c0",
X"8c08fa05",
X"2283c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08bf2691",
X"3883c08c",
X"08e40508",
X"880783c0",
X"8c08e405",
X"0c81c00b",
X"83c08c08",
X"ffa40508",
X"27913883",
X"c08c08e4",
X"05088407",
X"83c08c08",
X"e4050c80",
X"0b83c08c",
X"08ffb005",
X"0c83c08c",
X"08ffb005",
X"081083c0",
X"8c08c405",
X"08057090",
X"05703383",
X"c08c08c0",
X"05080570",
X"33728105",
X"33707206",
X"51535183",
X"c08c08ff",
X"a8050c51",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9b38",
X"900b83c0",
X"8c08ffb0",
X"05082b83",
X"c08c08e4",
X"05080783",
X"c08c08e4",
X"050c83c0",
X"8c08ffb0",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa4050c",
X"970b83c0",
X"8c08ffb0",
X"050827fe",
X"f43883c0",
X"8c08ffb8",
X"05089005",
X"3383c08c",
X"08e40508",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"c4050c83",
X"c08c08ff",
X"b4050883",
X"c08c08ff",
X"b805088c",
X"05082e83",
X"ff3883c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffb8",
X"05088c05",
X"0c83c08c",
X"08ffb805",
X"08890533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e83b9",
X"3883c08c",
X"08e40583",
X"c08c08ff",
X"b405088f",
X"0683c08c",
X"08e4050c",
X"83c08c08",
X"cc050c80",
X"0b83c08c",
X"08f0050c",
X"800b83c0",
X"8c08f405",
X"23800b81",
X"d7e83383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"bc05082e",
X"82d33883",
X"c08c08f0",
X"0581d7e8",
X"0b83c08c",
X"08ffac05",
X"0c83c08c",
X"08d0050c",
X"83c08c08",
X"ffac0508",
X"3383c08c",
X"08ffac05",
X"08810533",
X"81722b81",
X"722b0770",
X"83c08c08",
X"ffb40508",
X"065283c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffa8",
X"05082e09",
X"810681be",
X"3883c08c",
X"08ffbc05",
X"08852680",
X"f63883c0",
X"8c08ffac",
X"05088205",
X"337081ff",
X"0683c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa405",
X"08802e80",
X"ca3883c0",
X"8c08ffbc",
X"050883c0",
X"8c08ffbc",
X"05088105",
X"7081ff06",
X"83c08c08",
X"d0050873",
X"055383c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb0",
X"050883c0",
X"8c08ffa4",
X"05083483",
X"c08c08ff",
X"ac050883",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"9d38810b",
X"83c08c08",
X"ffa40508",
X"2b83c08c",
X"08cc0508",
X"080783c0",
X"8c08cc05",
X"080c83c0",
X"8c08ffac",
X"05088405",
X"703383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa4",
X"0508fdc8",
X"3883c08c",
X"08f00552",
X"8051d0c3",
X"3f83c08c",
X"08e40508",
X"5283c08c",
X"08c40508",
X"51d1fe3f",
X"83c08c08",
X"fb053370",
X"81800a29",
X"810a0570",
X"982c5583",
X"c08c08ff",
X"a4050c83",
X"c08c08f9",
X"05337081",
X"800a2981",
X"0a057098",
X"2c5583c0",
X"8c08ffa4",
X"050c83c0",
X"8c08c405",
X"085383c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa8",
X"050cd1d4",
X"3f83c08c",
X"08ffb805",
X"08880533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e84e0",
X"3883c08c",
X"08ffb805",
X"08900533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"812684c0",
X"38807081",
X"d89c0b81",
X"d89c0b81",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffb4",
X"05082e81",
X"ae3883c0",
X"8c08ffac",
X"05088429",
X"83c08c08",
X"ffa80508",
X"05703383",
X"c08c08c0",
X"05080570",
X"33728105",
X"33707206",
X"51535183",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2eaa3881",
X"0b83c08c",
X"08ffac05",
X"082b83c0",
X"8c08ffb4",
X"05080770",
X"83ffff06",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffac0508",
X"81057081",
X"ff0681d8",
X"9c718429",
X"71057081",
X"05335153",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"fed43883",
X"c08c08ff",
X"b805088a",
X"052283c0",
X"8c08c005",
X"0c83c08c",
X"08ffb405",
X"0883c08c",
X"08c00508",
X"2e82ad38",
X"800b83c0",
X"8c08e805",
X"0c800b83",
X"c08c08ec",
X"05238070",
X"83c08c08",
X"e80583c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffb0",
X"050c81af",
X"3983c08c",
X"08ffb405",
X"0883c08c",
X"08ffac05",
X"082c7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"80e73883",
X"c08c08ff",
X"b0050883",
X"c08c08ff",
X"b0050881",
X"057081ff",
X"0683c08c",
X"08ffbc05",
X"08730583",
X"c08c08ff",
X"b8050890",
X"053383c0",
X"8c08ffac",
X"05088429",
X"05535383",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a8050881",
X"d89e0533",
X"83c08c08",
X"ffa40508",
X"3483c08c",
X"08ffac05",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a4050c8f",
X"0b83c08c",
X"08ffac05",
X"082783c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb0",
X"05088526",
X"8c3883c0",
X"8c08ffa4",
X"0508fea9",
X"3883c08c",
X"08e80552",
X"8051caf3",
X"3f83c08c",
X"08ffb405",
X"0883c08c",
X"08ffb805",
X"088a0523",
X"83c08c08",
X"ffb80508",
X"80d20533",
X"83c08c08",
X"ffb80508",
X"80d40508",
X"0583c08c",
X"08ffb805",
X"0880d405",
X"0c83c08c",
X"08d80508",
X"0d83c08c",
X"08d40508",
X"81800a29",
X"81800a05",
X"70982c83",
X"c08c08c8",
X"05088105",
X"3383c08c",
X"08ffa805",
X"0c5183c0",
X"8c08d405",
X"0c83c08c",
X"08ffa805",
X"0883c08c",
X"08d40508",
X"24ec8538",
X"800b83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08dc05",
X"080d83c0",
X"8c08ffa8",
X"050883c0",
X"800c9c3d",
X"0d83c08c",
X"0c04f33d",
X"0d02bf05",
X"33028405",
X"80c30533",
X"83cb8c33",
X"5a5b5979",
X"802e8d38",
X"78780657",
X"76802e8e",
X"38818939",
X"78780657",
X"76802e80",
X"ff3883cb",
X"8c33707a",
X"07585879",
X"88387809",
X"70790651",
X"577683cb",
X"8c349297",
X"3f83c080",
X"085e805c",
X"8f5d7d1c",
X"87113358",
X"5876802e",
X"80c13877",
X"0881d5ec",
X"2e098106",
X"b638805b",
X"815a7d1c",
X"701c9a11",
X"33595959",
X"76822e09",
X"81069438",
X"83cb8c56",
X"81558054",
X"76539718",
X"33527851",
X"cbc53fff",
X"1a80d81c",
X"5c5a7980",
X"25d038ff",
X"1d81c41d",
X"5d5d7c80",
X"25ffa738",
X"8f3d0d04",
X"e93d0d69",
X"6c028805",
X"80ea0522",
X"5c5a5b80",
X"7071415e",
X"58ff7879",
X"7a7b7c7d",
X"464c4a45",
X"405d4362",
X"993d3462",
X"02840580",
X"dd053477",
X"792280ff",
X"ff065445",
X"72792379",
X"782e8887",
X"387a7081",
X"055c3370",
X"842a718c",
X"0670822a",
X"5a565683",
X"06ff1b70",
X"83ffff06",
X"5c545680",
X"5475742e",
X"91387a70",
X"81055c33",
X"ff1b7083",
X"ffff065c",
X"54548176",
X"279b3873",
X"81ff067b",
X"7081055d",
X"33557482",
X"802905ff",
X"1b7083ff",
X"ff065c54",
X"54827627",
X"aa387383",
X"ffff067b",
X"7081055d",
X"3370902b",
X"72077d70",
X"81055f33",
X"70982b72",
X"07fe1f70",
X"83ffff06",
X"40525252",
X"5254547e",
X"802e80c4",
X"387686f7",
X"38748a2e",
X"09810694",
X"38811f70",
X"81ff0681",
X"1e7081ff",
X"065f5240",
X"5386dc39",
X"748c2e09",
X"810686d3",
X"38ff1f70",
X"81ff06ff",
X"1e7081ff",
X"065f5240",
X"537b6325",
X"86bd38ff",
X"4386b839",
X"76812e83",
X"bb387681",
X"24893876",
X"802e8d38",
X"86a53976",
X"822e84a6",
X"38869c39",
X"f8155372",
X"84268495",
X"38728429",
X"81d8dc05",
X"53720804",
X"64802e80",
X"cd387822",
X"83808006",
X"53728380",
X"802e0981",
X"06bc3880",
X"56756427",
X"a438751e",
X"7083ffff",
X"0677101b",
X"90117283",
X"2a585157",
X"51537375",
X"34728706",
X"81712b51",
X"53728116",
X"34811670",
X"81ff0657",
X"53977627",
X"cc387f84",
X"0740800b",
X"993d4356",
X"61167033",
X"70982b70",
X"982c5151",
X"51538073",
X"2480fb38",
X"6073291e",
X"7083ffff",
X"067a2283",
X"80800652",
X"58537283",
X"80802e09",
X"810680de",
X"38608832",
X"70307072",
X"07802563",
X"90327030",
X"70720780",
X"25730753",
X"54585155",
X"5373802e",
X"bd387687",
X"065372b6",
X"38758429",
X"76100579",
X"11841179",
X"832a5757",
X"51537375",
X"34608116",
X"34658614",
X"23668814",
X"23758738",
X"7f810740",
X"8d397581",
X"2e098106",
X"85387f82",
X"07408116",
X"7081ff06",
X"57538176",
X"27fee538",
X"6361291e",
X"7083ffff",
X"065f5380",
X"704642ff",
X"02840580",
X"dd0534ff",
X"0b993d34",
X"83f53981",
X"1c7081ff",
X"065d5380",
X"4273812e",
X"0981068e",
X"38778180",
X"0a298180",
X"0a055880",
X"d3397380",
X"2e893873",
X"822e0981",
X"068d387c",
X"81800a29",
X"81800a05",
X"5da43981",
X"5f83b839",
X"ff1c7081",
X"ff065d53",
X"7b632583",
X"38ff437c",
X"802e9238",
X"7c81800a",
X"2981ff0a",
X"055d7c98",
X"2c5d8393",
X"3977802e",
X"92387781",
X"800a2981",
X"ff0a0558",
X"77982c58",
X"82fd3977",
X"53839e39",
X"74892680",
X"f4387484",
X"2981d8f0",
X"05537208",
X"0473872e",
X"82e13873",
X"852e82db",
X"3873882e",
X"82d53873",
X"8c2e82cf",
X"3873892e",
X"09810686",
X"38814582",
X"c2397381",
X"2e098106",
X"82b93862",
X"802582b3",
X"387b982b",
X"70982c51",
X"4382a839",
X"7383ffff",
X"0646829f",
X"397383ff",
X"ff064782",
X"96397381",
X"ff064182",
X"8e397381",
X"1a348287",
X"397381ff",
X"064481ff",
X"397e5382",
X"a0397481",
X"2e81e338",
X"74812489",
X"3874802e",
X"8d3881e7",
X"3974822e",
X"81d83881",
X"de397456",
X"7b833881",
X"56745373",
X"862e0981",
X"06973875",
X"81065372",
X"802e8e38",
X"782282ff",
X"ff06fe80",
X"800753b6",
X"397b8338",
X"81537382",
X"2e098106",
X"97387281",
X"06537280",
X"2e8e3878",
X"2281ffff",
X"06818080",
X"07539339",
X"7b9638fc",
X"14537281",
X"268e3878",
X"22ff8080",
X"07537279",
X"2380e539",
X"80557381",
X"2e098106",
X"83387355",
X"77537780",
X"2e893874",
X"81065372",
X"80ca3872",
X"d0155455",
X"72812683",
X"38815577",
X"802eb938",
X"74810653",
X"72802eb0",
X"38782283",
X"80800653",
X"72838080",
X"2e098106",
X"9f3873b0",
X"2e098106",
X"87386199",
X"3d349139",
X"73b12e09",
X"81068938",
X"61028405",
X"80dd0534",
X"61810553",
X"8c396174",
X"31810553",
X"84396114",
X"537283ff",
X"ff064279",
X"f7fb387d",
X"832a5372",
X"821a3478",
X"22838080",
X"06537283",
X"80802e09",
X"81068838",
X"81537f87",
X"2e833880",
X"537283c0",
X"800c993d",
X"0d04fd3d",
X"0d758311",
X"33821233",
X"71982b71",
X"902b0781",
X"14337088",
X"2b720775",
X"33710783",
X"c0800c52",
X"53545654",
X"52853d0d",
X"04f63d0d",
X"02b70533",
X"028405bb",
X"05330288",
X"05bf0533",
X"5b5b5b80",
X"58805778",
X"882b7a07",
X"5680557a",
X"548153a3",
X"527c5192",
X"cc3f83c0",
X"800881ff",
X"0683c080",
X"0c8c3d0d",
X"04f63d0d",
X"02b70533",
X"028405bb",
X"05330288",
X"05bf0533",
X"5b5b5b80",
X"58805778",
X"882b7a07",
X"5680557a",
X"548353a3",
X"527c5192",
X"903f83c0",
X"800881ff",
X"0683c080",
X"0c8c3d0d",
X"04f73d0d",
X"02b30533",
X"028405b6",
X"0522605a",
X"58568055",
X"80548053",
X"81a3527b",
X"5191e23f",
X"83c08008",
X"81ff0683",
X"c0800c8b",
X"3d0d04ee",
X"3d0d6490",
X"115c5c80",
X"7b34800b",
X"841c0c80",
X"0b881c34",
X"810b891c",
X"34880b8a",
X"1c34800b",
X"8b1c3488",
X"1b08c106",
X"8107881c",
X"0c8f3d70",
X"545d8852",
X"7b519beb",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"81a93890",
X"3d335e81",
X"db5a7d89",
X"2e098106",
X"8199387c",
X"5392527b",
X"519bc43f",
X"83c08008",
X"81ff0670",
X"5b597881",
X"82387c58",
X"88577856",
X"a9557854",
X"865381a0",
X"527b5190",
X"d03f83c0",
X"800881ff",
X"06705b59",
X"7880e038",
X"02ba0533",
X"7b347c54",
X"78537d52",
X"7b519bac",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"80c13802",
X"bd053352",
X"7b519bc4",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"aa38817b",
X"335a5a79",
X"79269938",
X"80547953",
X"88527b51",
X"fdbb3f81",
X"1a7081ff",
X"067c3352",
X"5b59e439",
X"810b881c",
X"34805a79",
X"83c0800c",
X"943d0d04",
X"800b83c0",
X"800c04f9",
X"3d0d7902",
X"8405ab05",
X"338e3d70",
X"54585858",
X"ffbeb03f",
X"8a3d8a05",
X"51ffbea7",
X"3f7551fc",
X"8d3f83c0",
X"80088486",
X"812ebe38",
X"83c08008",
X"84868126",
X"993883c0",
X"80088482",
X"802e80e6",
X"3883c080",
X"08848281",
X"2e9f3881",
X"b43983c0",
X"800880c0",
X"82832e80",
X"f43883c0",
X"800880c0",
X"86832e80",
X"e8388199",
X"3983c09c",
X"33558056",
X"74762e09",
X"8106818b",
X"38745476",
X"53915277",
X"51fbd63f",
X"74547653",
X"90527751",
X"fbcb3f74",
X"54765384",
X"527751fb",
X"fc3f810b",
X"83c09c34",
X"81b15680",
X"de398054",
X"76539152",
X"7751fba9",
X"3f805476",
X"53905277",
X"51fb9e3f",
X"800b83c0",
X"9c347652",
X"87183351",
X"97963fb5",
X"39805476",
X"53945277",
X"51fb823f",
X"80547653",
X"90527751",
X"faf73f75",
X"51ffbcdb",
X"3f83c080",
X"08892a81",
X"06537652",
X"87183351",
X"90cd3f80",
X"0b83c09c",
X"34805675",
X"83c0800c",
X"893d0d04",
X"f23d0d60",
X"90115a58",
X"800b881a",
X"33715956",
X"5674762e",
X"82a53882",
X"ac3f8419",
X"0883c080",
X"08268295",
X"3878335a",
X"810b8e3d",
X"23903df8",
X"1155f405",
X"53991852",
X"77518ae5",
X"3f83c080",
X"0881ff06",
X"70575574",
X"772e0981",
X"0681d938",
X"86397456",
X"81d23981",
X"5682578e",
X"3d337706",
X"5574802e",
X"bb38800b",
X"8d3d3490",
X"3df00554",
X"84537552",
X"7751facd",
X"3f83c080",
X"0881ff06",
X"55749d38",
X"7b537552",
X"7751fce7",
X"3f83c080",
X"0881ff06",
X"557481b1",
X"2e818b38",
X"74ffb338",
X"761081fc",
X"06811770",
X"81ff0658",
X"56578776",
X"27ffa838",
X"8156757a",
X"2680eb38",
X"800b8d3d",
X"348c3d70",
X"55578453",
X"75527751",
X"f9f73f83",
X"c0800881",
X"ff065574",
X"80c13876",
X"51ffbad7",
X"3f83c080",
X"08828706",
X"55748281",
X"2e098106",
X"aa3802ae",
X"05338107",
X"55740284",
X"05ae0534",
X"7b537552",
X"7751fbeb",
X"3f83c080",
X"0881ff06",
X"557481b1",
X"2e903874",
X"feb83881",
X"167081ff",
X"065755ff",
X"91398056",
X"7581ff06",
X"56973f83",
X"c080088f",
X"d005841a",
X"0c755776",
X"83c0800c",
X"903d0d04",
X"049080a0",
X"0883c080",
X"0c04ff3d",
X"0d7387e8",
X"2951ff90",
X"9e3f833d",
X"0d040483",
X"cb900b83",
X"c0800c04",
X"fd3d0d75",
X"77545480",
X"0b83caf0",
X"34728a38",
X"9090800b",
X"84150c90",
X"3972812e",
X"09810688",
X"38909880",
X"0b84150c",
X"84140883",
X"cb880c80",
X"0b88150c",
X"800b8c15",
X"0c83cb88",
X"0853820b",
X"87801434",
X"8151ff9e",
X"3f83cb88",
X"0853800b",
X"88143483",
X"cb880853",
X"810b8780",
X"143483cb",
X"88085380",
X"0b8c1434",
X"83cb8808",
X"53800ba4",
X"14349174",
X"34800b83",
X"c0a03480",
X"0b83c0a4",
X"34800b83",
X"c0a83480",
X"547381c4",
X"2983cb94",
X"0553800b",
X"83143481",
X"147081ff",
X"0655538f",
X"7427e638",
X"853d0d04",
X"fe3d0d74",
X"76821133",
X"70bf0681",
X"712bff05",
X"56515152",
X"53907127",
X"8338ff52",
X"76517171",
X"2383cb88",
X"08518713",
X"33901234",
X"800b83c0",
X"a434800b",
X"83c0a834",
X"8813338a",
X"14335252",
X"71802eaa",
X"387081ff",
X"06518452",
X"70833870",
X"527183c0",
X"a4348a13",
X"33703070",
X"8025842b",
X"70880751",
X"51525370",
X"83c0a834",
X"90397081",
X"ff065170",
X"83389852",
X"7183c0a8",
X"34800b83",
X"c0800c84",
X"3d0d04f1",
X"3d0d6165",
X"68028c05",
X"80cb0533",
X"02900580",
X"ce052202",
X"940580d6",
X"05224240",
X"415a4040",
X"fd8b3f83",
X"c08008a7",
X"88055b80",
X"70715b5b",
X"52839439",
X"83cb8808",
X"517d9412",
X"3483c0a4",
X"33810755",
X"80705456",
X"7f862680",
X"ea387f84",
X"2981d9a4",
X"0583cb88",
X"08535170",
X"0804800b",
X"841334a1",
X"39773370",
X"30708025",
X"83713151",
X"51525370",
X"8413348d",
X"39810b84",
X"1334b839",
X"830b8413",
X"34817054",
X"56ad3981",
X"0b841334",
X"a2397733",
X"70307080",
X"25837131",
X"51515253",
X"70841334",
X"80783352",
X"52708338",
X"81527178",
X"34815374",
X"88075583",
X"c0a83383",
X"cb880852",
X"57810b81",
X"d0123483",
X"cb880851",
X"810b8190",
X"12347e80",
X"2eae3872",
X"802ea938",
X"7eff1e52",
X"547083ff",
X"ff065372",
X"83ffff2e",
X"97387370",
X"81055533",
X"83cb8808",
X"53517081",
X"c01334ff",
X"1351de39",
X"83cb8808",
X"a8113353",
X"51768812",
X"3483cb88",
X"08517471",
X"3481ff52",
X"913983cb",
X"8808a011",
X"33708106",
X"51525370",
X"8f38fafd",
X"3f7a83c0",
X"800826e6",
X"38818839",
X"810ba014",
X"3483cb88",
X"08a81133",
X"80ff0670",
X"78075253",
X"5170802e",
X"80ed3871",
X"862a7081",
X"06515170",
X"802e9138",
X"80783352",
X"53708338",
X"81537278",
X"3480e039",
X"71842a70",
X"81065151",
X"70802e9b",
X"38811970",
X"83ffff06",
X"7d30709f",
X"2a51525a",
X"51787c2e",
X"098106af",
X"38a43971",
X"832a7081",
X"06515170",
X"802e9338",
X"811a7081",
X"ff065b51",
X"79832e09",
X"81069038",
X"8a3971a3",
X"06517080",
X"2e853871",
X"519239f9",
X"e43f7a83",
X"c0800826",
X"fce23871",
X"81bf0651",
X"7083c080",
X"0c913d0d",
X"04f63d0d",
X"02b30533",
X"028405b7",
X"05330288",
X"05ba0522",
X"59595980",
X"0b8c3d34",
X"8c3dfc05",
X"56805580",
X"54765377",
X"527851fb",
X"f23f83c0",
X"800881ff",
X"0683c080",
X"0c8c3d0d",
X"04f33d0d",
X"7f626402",
X"8c0580c2",
X"05227222",
X"81153342",
X"5f415e59",
X"59807823",
X"7d537833",
X"528151ff",
X"a03f83c0",
X"800881ff",
X"06567580",
X"2e863875",
X"5481ad39",
X"83cb8808",
X"a8113382",
X"1b337086",
X"2a708106",
X"73982b53",
X"51575c56",
X"57798025",
X"83388156",
X"73762e87",
X"3881f054",
X"81823981",
X"8c173370",
X"81ff0679",
X"227d7131",
X"902b7090",
X"2c700970",
X"9f2c7206",
X"70525253",
X"51535757",
X"54757424",
X"83387555",
X"74848080",
X"29fc8080",
X"0570902c",
X"515574ff",
X"2e943883",
X"cb880881",
X"80113351",
X"54737c70",
X"81055e34",
X"db397722",
X"76055473",
X"78237909",
X"709f2a70",
X"8106821c",
X"3381bf06",
X"71862b07",
X"51515154",
X"73821a34",
X"7c76268a",
X"38772254",
X"7a7426fe",
X"bb388054",
X"7383c080",
X"0c8f3d0d",
X"04f93d0d",
X"7a57800b",
X"893d2389",
X"3dfc0553",
X"76527951",
X"f8da3f83",
X"c0800881",
X"ff067057",
X"55749638",
X"7c547b53",
X"883d2252",
X"7651fde5",
X"3f83c080",
X"0881ff06",
X"567583c0",
X"800c893d",
X"0d04f03d",
X"0d626602",
X"880580ce",
X"0522415d",
X"5e800284",
X"0580d205",
X"227f8105",
X"33ff115a",
X"5d5a5d81",
X"da5876bf",
X"2680e938",
X"78802e80",
X"e1387a58",
X"787b2783",
X"38785882",
X"1e337087",
X"2a585a76",
X"923d3492",
X"3dfc0556",
X"77557b54",
X"7e537d33",
X"528251f8",
X"de3f83c0",
X"800881ff",
X"065d800b",
X"923d3358",
X"5a76802e",
X"8338815a",
X"821e3380",
X"ff067a87",
X"2b075776",
X"821f347c",
X"91387878",
X"317083ff",
X"ff06791e",
X"5e5a57ff",
X"9b397c58",
X"7783c080",
X"0c923d0d",
X"04f83d0d",
X"7b028405",
X"b2052258",
X"58800b8a",
X"3d238a3d",
X"fc055377",
X"527a51f6",
X"f73f83c0",
X"800881ff",
X"06705755",
X"7496387d",
X"54765389",
X"3d225277",
X"51feaf3f",
X"83c08008",
X"81ff0656",
X"7583c080",
X"0c8a3d0d",
X"04ec3d0d",
X"666e0288",
X"0580df05",
X"33028c05",
X"80e30533",
X"02900580",
X"e7053302",
X"940580eb",
X"05330298",
X"0580ee05",
X"22414341",
X"5f5c4057",
X"0280f205",
X"22963d23",
X"963df005",
X"53841770",
X"53775259",
X"f6863f83",
X"c0800881",
X"ff065877",
X"81e53877",
X"7a818006",
X"58408077",
X"25833881",
X"4079943d",
X"347b0284",
X"0580c905",
X"347c0284",
X"0580ca05",
X"347d0284",
X"0580cb05",
X"347a953d",
X"347a882a",
X"57760284",
X"0580cd05",
X"34953d22",
X"57760284",
X"0580ce05",
X"3476882a",
X"57760284",
X"0580cf05",
X"3477923d",
X"34963dec",
X"11575788",
X"55f41754",
X"923d2253",
X"77527751",
X"f6953f83",
X"c0800881",
X"ff065877",
X"80ed387e",
X"802e80cb",
X"38923d22",
X"79085858",
X"7f802e9c",
X"38768180",
X"8007790c",
X"7e54963d",
X"fc055377",
X"83ffff06",
X"527851f9",
X"fc3f9939",
X"76828080",
X"07790c7e",
X"54953d22",
X"537783ff",
X"ff065278",
X"51fc8f3f",
X"83c08008",
X"81ff0658",
X"779d3892",
X"3d225380",
X"527f3070",
X"80258471",
X"31535157",
X"f9873f83",
X"c0800881",
X"ff065877",
X"83c0800c",
X"963d0d04",
X"f63d0d7c",
X"028405b7",
X"05335b5b",
X"80588057",
X"80568055",
X"79548553",
X"80527a51",
X"fda33f83",
X"c0800881",
X"ff065978",
X"85387987",
X"1c347883",
X"c0800c8c",
X"3d0d04f9",
X"3d0d02a7",
X"05330284",
X"05ab0533",
X"028805af",
X"05335859",
X"57800b83",
X"cb973354",
X"5472742e",
X"9f388114",
X"7081ff06",
X"5553738f",
X"2681b638",
X"7381c429",
X"83cb9405",
X"83113351",
X"5372e338",
X"7381c429",
X"83cb9005",
X"55800b87",
X"16347688",
X"1634758a",
X"16347789",
X"16348075",
X"0c83cb88",
X"088c160c",
X"800b8416",
X"34880b85",
X"1634800b",
X"86163484",
X"1508ffa1",
X"ff06a080",
X"0784160c",
X"81147081",
X"ff065353",
X"7451febc",
X"3f83c080",
X"0881ff06",
X"70555372",
X"80cd388a",
X"39730875",
X"0c725480",
X"c2397281",
X"dfd85556",
X"81dfd808",
X"802eb238",
X"75842914",
X"70087653",
X"70085154",
X"54722d83",
X"c0800881",
X"ff065372",
X"802ece38",
X"81167081",
X"ff0681df",
X"d8718429",
X"11535657",
X"537208d0",
X"38805473",
X"83c0800c",
X"893d0d04",
X"f93d0d79",
X"57800b84",
X"180883cb",
X"880c58f0",
X"883f8817",
X"0883c080",
X"082783ed",
X"38effa3f",
X"83c08008",
X"81058818",
X"0c83cb88",
X"08b81133",
X"7081ff06",
X"51515473",
X"812ea438",
X"73812488",
X"3873782e",
X"8a38b839",
X"73822e95",
X"38b13976",
X"3381f006",
X"5473902e",
X"a6389177",
X"34a13973",
X"58763381",
X"f0065473",
X"902e0981",
X"069138ef",
X"a83f83c0",
X"800881c8",
X"058c180c",
X"a0773480",
X"567581c4",
X"2983cb97",
X"11335555",
X"73802eaa",
X"3883cb90",
X"15700856",
X"5474802e",
X"9d388815",
X"08802e96",
X"388c1408",
X"83cb8808",
X"2e098106",
X"89387351",
X"88150854",
X"732d8116",
X"7081ff06",
X"57548f76",
X"27ffba38",
X"76335473",
X"b02e8199",
X"3873b024",
X"8f387391",
X"2eab3873",
X"a02e80f5",
X"3882a639",
X"7380d02e",
X"81e43873",
X"80d0248b",
X"387380c0",
X"2e819938",
X"828f3973",
X"81802e81",
X"fb388285",
X"39805675",
X"81c42983",
X"cb941183",
X"11335659",
X"5573802e",
X"a83883cb",
X"90157008",
X"56547480",
X"2e9b388c",
X"140883cb",
X"88082e09",
X"81068e38",
X"73518415",
X"0854732d",
X"800b8319",
X"34811670",
X"81ff0657",
X"548f7627",
X"ffb93892",
X"773481b5",
X"39edc23f",
X"8c170883",
X"c0800827",
X"81a738b0",
X"773481a1",
X"3983cb88",
X"0854800b",
X"8c153483",
X"cb880854",
X"840b8815",
X"3480c077",
X"34ed963f",
X"83c08008",
X"b2058c18",
X"0c80fa39",
X"ed873f8c",
X"170883c0",
X"80082780",
X"ec3883cb",
X"88085481",
X"0b8c1534",
X"83cb8808",
X"54800b88",
X"153483cb",
X"88085488",
X"0ba01534",
X"ecdb3f83",
X"c0800894",
X"058c180c",
X"80d07734",
X"bc3983cb",
X"8808a011",
X"3370832a",
X"70810651",
X"51555573",
X"802ea638",
X"880ba016",
X"34ecae3f",
X"8c170883",
X"c0800827",
X"9438ff80",
X"77348e39",
X"77538052",
X"8051fa8b",
X"3fff9077",
X"3483cb88",
X"08a01133",
X"70832a70",
X"81065151",
X"55557380",
X"2e863888",
X"0ba01634",
X"893d0d04",
X"f63d0d02",
X"b3053302",
X"8405b705",
X"335b5b80",
X"0b83cb94",
X"70841272",
X"745d5957",
X"5b585683",
X"15335372",
X"802e80f3",
X"38733353",
X"7a732e09",
X"810680e7",
X"38811433",
X"5379732e",
X"09810680",
X"da388055",
X"7481c429",
X"83cb9805",
X"7033831b",
X"33585553",
X"73762e09",
X"81068a38",
X"81133352",
X"7351ff9c",
X"3f811570",
X"81ff0656",
X"538f7527",
X"d338800b",
X"83cb9019",
X"70085654",
X"5573752e",
X"91387251",
X"84140853",
X"722d83c0",
X"800881ff",
X"0655800b",
X"83183474",
X"53a03981",
X"1681c419",
X"81c41781",
X"c41781c4",
X"1d81c41c",
X"5c5d5757",
X"59568f76",
X"25fee838",
X"80537283",
X"c0800c8c",
X"3d0d04f8",
X"3d0d02ae",
X"05227d59",
X"57805681",
X"55805486",
X"53818052",
X"7a51f595",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8a3d0d04",
X"f73d0d02",
X"b2052202",
X"8405b705",
X"33605a5b",
X"57805682",
X"55795486",
X"53818052",
X"7b51f4e5",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8b3d0d04",
X"f83d0d02",
X"af053359",
X"80588057",
X"80568055",
X"78548953",
X"80527a51",
X"f4bb3f83",
X"c0800881",
X"ff0683c0",
X"800c8a3d",
X"0d040000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002b19",
X"00002b5a",
X"00002b7c",
X"00002b9e",
X"00002bc4",
X"00002bc4",
X"00002bc4",
X"00002bc4",
X"00002c35",
X"00002c86",
X"000041fb",
X"00004a3f",
X"00004af8",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3f00",
X"0c0c4000",
X"0a0a4100",
X"0b0b4100",
X"07074100",
X"0a0b4300",
X"080b4200",
X"04044500",
X"05054400",
X"06060004",
X"08080004",
X"09090004",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"00005784",
X"00005a8b",
X"00005897",
X"00005a8b",
X"000058d4",
X"00005925",
X"00005964",
X"0000596d",
X"00005a8b",
X"00005a8b",
X"00005a8b",
X"00005a8b",
X"00005976",
X"0000597e",
X"00005985",
X"00005b8b",
X"00005c84",
X"00005d98",
X"0000608e",
X"000060a9",
X"00006095",
X"000060a9",
X"000060b0",
X"000060bb",
X"000060c2",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"43505520",
X"54757262",
X"6f3a2564",
X"78000000",
X"44726976",
X"65205475",
X"72626f3a",
X"25730000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"66726565",
X"7a65722e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"5374616e",
X"64617264",
X"00000000",
X"46617374",
X"28362900",
X"46617374",
X"28352900",
X"46617374",
X"28342900",
X"46617374",
X"28332900",
X"46617374",
X"28322900",
X"46617374",
X"28312900",
X"46617374",
X"28302900",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00006d00",
X"00006d04",
X"00006d0c",
X"00006d18",
X"00006d24",
X"00006d30",
X"00006d3c",
X"00006d40",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00000028",
X"00000006",
X"00000005",
X"00000004",
X"00000003",
X"00000002",
X"00000001",
X"00000000",
X"00006de0",
X"00006dec",
X"00006df4",
X"00006dfc",
X"00006e04",
X"00006e0c",
X"00006e14",
X"00006e1c",
X"00006c98",
X"00006aec",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"69383030",
X"00000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
