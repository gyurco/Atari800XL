
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f2",
X"c0738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80f5",
X"f40c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f0",
X"802d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580efbf",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80dad004",
X"fd3d0d75",
X"705254ae",
X"a53f83e0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83e0",
X"8008732e",
X"a13883e0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183e0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83e2c008",
X"248a38b4",
X"f63fff0b",
X"83e2c00c",
X"800b83e0",
X"800c04ff",
X"3d0d7352",
X"83e09c08",
X"722e8d38",
X"d93f7151",
X"96993f71",
X"83e09c0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"558154bc",
X"15088191",
X"387451cf",
X"3f795880",
X"7a2580f7",
X"3883e2f0",
X"0870892a",
X"5783ff06",
X"78848072",
X"31565657",
X"73782583",
X"38735575",
X"83e2c008",
X"2e8438ff",
X"893f83e2",
X"c0088025",
X"a6387589",
X"2b5198dc",
X"3f83e2f0",
X"088f3dfc",
X"11555c54",
X"8152f81b",
X"5196c63f",
X"761483e2",
X"f00c7583",
X"e2c00c74",
X"53765278",
X"51b3a73f",
X"83e08008",
X"83e2f008",
X"1683e2f0",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8b3861",
X"7a710c54",
X"75547580",
X"2e833881",
X"547383e0",
X"800c8e3d",
X"0d04fc3d",
X"0dfe9b3f",
X"7651feaf",
X"3f863dfc",
X"05537852",
X"775195e9",
X"3f797571",
X"0c5483e0",
X"80085483",
X"e0800880",
X"2e833881",
X"547383e0",
X"800c863d",
X"0d04fe3d",
X"0d7583e2",
X"c0085353",
X"80722489",
X"3871732e",
X"8438fdd6",
X"3f7451fd",
X"ea3f7251",
X"97ae3f83",
X"e0800852",
X"83e08008",
X"802e8338",
X"81527183",
X"e0800c84",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"e0800c51",
X"823d0d04",
X"80c40b83",
X"e0800c04",
X"fd3d0d75",
X"77715470",
X"535553a9",
X"fd3f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfceb3f",
X"735193ab",
X"3f7383e0",
X"9c0c83e0",
X"80085383",
X"e0800880",
X"2e833881",
X"537283e0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcbf3f",
X"72802ea5",
X"38bc1308",
X"527351a9",
X"873f83e0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"e0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83e0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83e2c0",
X"0c7483e0",
X"a00c7583",
X"e2bc0caf",
X"db3f83e0",
X"800881ff",
X"06528153",
X"71993883",
X"e2d8518e",
X"943f83e0",
X"80085283",
X"e0800880",
X"2e833872",
X"52715372",
X"83e0800c",
X"843d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"51a6f83f",
X"83e08008",
X"557483e0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"e0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283e2bc",
X"085180de",
X"c23f83e0",
X"800857f9",
X"e13f7952",
X"83e2c451",
X"95b73f83",
X"e0800854",
X"805383e0",
X"8008732e",
X"09810682",
X"833883e0",
X"a0080b0b",
X"80f3f453",
X"705256a6",
X"b53f0b0b",
X"80f3f452",
X"80c01651",
X"a6a83f75",
X"bc170c73",
X"82c0170c",
X"810b82c4",
X"170c810b",
X"82c8170c",
X"7382cc17",
X"0cff1782",
X"d0175557",
X"81913983",
X"e0ac3370",
X"822a7081",
X"06515455",
X"72818038",
X"74812a81",
X"06587780",
X"f6387484",
X"2a810682",
X"c4150c83",
X"e0ac3381",
X"0682c815",
X"0c795273",
X"51a5cf3f",
X"7351a5e6",
X"3f83e080",
X"081453af",
X"73708105",
X"553472bc",
X"150c83e0",
X"ad527251",
X"a5b03f83",
X"e0a40882",
X"c0150c83",
X"e0ba5280",
X"c01451a5",
X"9d3f7880",
X"2e8d3873",
X"51782d83",
X"e0800880",
X"2e993877",
X"82cc150c",
X"75802e86",
X"387382cc",
X"170c7382",
X"d015ff19",
X"59555676",
X"802e9b38",
X"83e0a452",
X"83e2c451",
X"94ad3f83",
X"e080088a",
X"3883e0ad",
X"335372fe",
X"d2387880",
X"2e893883",
X"e0a00851",
X"fcb83f83",
X"e0a00853",
X"7283e080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb53f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f690",
X"3f83e080",
X"08745387",
X"3d705355",
X"55f6b03f",
X"f7903f73",
X"51d33f63",
X"53745283",
X"e0800851",
X"fab83f92",
X"3d0d0471",
X"83e0800c",
X"0480c012",
X"83e0800c",
X"04803d0d",
X"7282c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"e0800c51",
X"823d0d04",
X"f93d0d79",
X"83e09008",
X"57578177",
X"27819638",
X"76881708",
X"27818e38",
X"75335574",
X"822e8938",
X"74832eb3",
X"3880fe39",
X"74547610",
X"83fe0653",
X"76882a8c",
X"17080552",
X"893dfc05",
X"51aa893f",
X"83e08008",
X"80df3802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d13984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"51a9d93f",
X"83e08008",
X"b038029f",
X"05330284",
X"059e0533",
X"71982b71",
X"902b0702",
X"8c059d05",
X"3370882b",
X"72078d3d",
X"337180ff",
X"fffe8006",
X"07515253",
X"57585683",
X"39815574",
X"83e0800c",
X"893d0d04",
X"fb3d0d83",
X"e09008fe",
X"19881208",
X"fe055556",
X"54805674",
X"73278d38",
X"82143375",
X"71299416",
X"08055753",
X"7583e080",
X"0c873d0d",
X"04fc3d0d",
X"7652800b",
X"83e09008",
X"70335152",
X"5370832e",
X"09810691",
X"38951233",
X"94133371",
X"982b7190",
X"2b075555",
X"519b1233",
X"9a133371",
X"882b0774",
X"0783e080",
X"0c55863d",
X"0d04fc3d",
X"0d7683e0",
X"90085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"fed63f83",
X"e0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183e080",
X"0c863d0d",
X"04fa3d0d",
X"7883e090",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fcb13f",
X"81527183",
X"e0800827",
X"a8388352",
X"83e08008",
X"88170827",
X"9c3883e0",
X"80088c16",
X"0c83e080",
X"0851fdbc",
X"3f83e080",
X"0890160c",
X"73752380",
X"527183e0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585e5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"9f269138",
X"7a51fdd2",
X"3f83e080",
X"0856807d",
X"34838139",
X"933d841c",
X"08705859",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"3880705a",
X"5c887f08",
X"5f5a7b81",
X"1d7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535e57",
X"557480e7",
X"3876ae2e",
X"09810683",
X"38815578",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675bb",
X"3888598b",
X"5affab39",
X"76982b55",
X"74802587",
X"3880f1d0",
X"173357ff",
X"9f175574",
X"99268938",
X"e0177081",
X"ff065855",
X"78811a70",
X"81ff0672",
X"1b535b57",
X"55767534",
X"fef8397b",
X"1e7f0c80",
X"5576a026",
X"83388155",
X"748b1934",
X"7a51fc82",
X"3f83e080",
X"0880f538",
X"a0547a22",
X"70852b83",
X"e0065455",
X"901b0852",
X"7c51a494",
X"3f83e080",
X"085783e0",
X"80088181",
X"387c3355",
X"74802e80",
X"f4388b1d",
X"3370832a",
X"70810651",
X"565674b4",
X"388b7d84",
X"1d0883e0",
X"8008595b",
X"5b58ff18",
X"5877ff2e",
X"9a387970",
X"81055b33",
X"79708105",
X"5b337171",
X"31525656",
X"75802ee2",
X"38863975",
X"802e9638",
X"7a51fbe5",
X"3fff8639",
X"83e08008",
X"5683e080",
X"08b63883",
X"39765684",
X"1b088b11",
X"33515574",
X"a7388b1d",
X"3370842a",
X"70810651",
X"56567489",
X"38835694",
X"39815690",
X"397c51fa",
X"943f83e0",
X"8008881c",
X"0cfd8139",
X"7583e080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"51a2d93f",
X"835683e0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"51a2ad3f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"7651a284",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583e080",
X"0c8a3d0d",
X"04eb3d0d",
X"675a800b",
X"83e0900c",
X"a1a63f83",
X"e0800881",
X"06558256",
X"7483ef38",
X"7475538f",
X"3d705357",
X"59feca3f",
X"83e08008",
X"81ff0657",
X"76812e09",
X"810680d4",
X"38905483",
X"be537452",
X"7551a198",
X"3f83e080",
X"0880c938",
X"8f3d3355",
X"74802e80",
X"c93802bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"33710770",
X"587b575e",
X"525e5759",
X"57fdee3f",
X"83e08008",
X"81ff0657",
X"76832e09",
X"81068638",
X"815682f2",
X"3976802e",
X"86388656",
X"82e839a4",
X"548d5378",
X"527551a0",
X"af3f8156",
X"83e08008",
X"82d43802",
X"be053302",
X"8405bd05",
X"3371882b",
X"07595d77",
X"ab380280",
X"ce053302",
X"840580cd",
X"05337198",
X"2b71902b",
X"07973d33",
X"70882b72",
X"07029405",
X"80cb0533",
X"71075452",
X"5e575956",
X"02b70533",
X"78712902",
X"8805b605",
X"33028c05",
X"b5053371",
X"882b0770",
X"1d707f8c",
X"050c5f59",
X"57595d8e",
X"3d33821b",
X"3402b905",
X"33903d33",
X"71882b07",
X"5a5c7884",
X"1b2302bb",
X"05330284",
X"05ba0533",
X"71882b07",
X"565c74ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"07515253",
X"575e5c74",
X"76317831",
X"79842a90",
X"3d335471",
X"71315356",
X"5680cfa7",
X"3f83e080",
X"08820570",
X"881c0c83",
X"e08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83e0900c",
X"80567583",
X"e0800c97",
X"3d0d04e9",
X"3d0d83e0",
X"90085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e53f83e0",
X"80085483",
X"e0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f489",
X"3f83e080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383e080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83e09008",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0e93f",
X"83e08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"833f83e0",
X"80085583",
X"e0800880",
X"2eff8938",
X"83e08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"519ad53f",
X"83e08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83e0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83e09008",
X"55568555",
X"73802e81",
X"e3388114",
X"33810653",
X"84557280",
X"2e81d538",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b9388214",
X"3370892b",
X"56537680",
X"2eb73874",
X"52ff1651",
X"80caa83f",
X"83e08008",
X"ff187654",
X"70535853",
X"80ca983f",
X"83e08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed63f83",
X"e0800853",
X"810b83e0",
X"8008278b",
X"38881408",
X"83e08008",
X"26883880",
X"0b811534",
X"b03983e0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc53f",
X"83e08008",
X"8c3883e0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683e0",
X"800805a8",
X"150c8055",
X"7483e080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83e09008",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1cf3f",
X"83e08008",
X"5583e080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef5",
X"3f83e080",
X"0888170c",
X"7551efa6",
X"3f83e080",
X"08557483",
X"e0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683e0",
X"9008802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f53f83e0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"96de3f83",
X"e0800841",
X"83e08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"eddf3f83",
X"e0800841",
X"83e08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"8e843f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f03f83e0",
X"80088332",
X"70307072",
X"079f2c83",
X"e0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"8c903f75",
X"83e0800c",
X"9e3d0d04",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"7751e0d2",
X"3f83e080",
X"0880d738",
X"78902e09",
X"810680ce",
X"3802ab05",
X"3380f5fc",
X"0b80f5fc",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ad388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"56848880",
X"80527751",
X"e0803f83",
X"e0800886",
X"3878752e",
X"85388056",
X"85398117",
X"33567583",
X"e0800c8e",
X"3d0d04fc",
X"3d0d7670",
X"52558b96",
X"3f83e080",
X"0815ff05",
X"5473752e",
X"8e387333",
X"5372ae2e",
X"8638ff14",
X"54ef3977",
X"52811451",
X"8aae3f83",
X"e0800830",
X"7083e080",
X"08078025",
X"83e0800c",
X"53863d0d",
X"04fc3d0d",
X"76705255",
X"e6ed3f83",
X"e0800854",
X"815383e0",
X"800880c1",
X"387451e6",
X"b03f83e0",
X"800880f4",
X"845383e0",
X"80085253",
X"ff913f83",
X"e08008a1",
X"3880f488",
X"527251ff",
X"823f83e0",
X"80089238",
X"80f48c52",
X"7251fef3",
X"3f83e080",
X"08802e83",
X"38815473",
X"537283e0",
X"800c863d",
X"0d04fd3d",
X"0d757052",
X"54e68c3f",
X"815383e0",
X"80089838",
X"7351e5d5",
X"3f83e388",
X"085283e0",
X"800851fe",
X"ba3f83e0",
X"80085372",
X"83e0800c",
X"853d0d04",
X"df3d0da4",
X"3d087052",
X"5edbfa3f",
X"83e08008",
X"33953d56",
X"54739638",
X"80f8f852",
X"7451898e",
X"3f9a397d",
X"527851de",
X"fb3f84cd",
X"397d51db",
X"e03f83e0",
X"80085274",
X"51db903f",
X"80438042",
X"80418040",
X"83e39008",
X"52943d70",
X"525de1e3",
X"3f83e080",
X"0859800b",
X"83e08008",
X"555b83e0",
X"80087b2e",
X"9438811b",
X"74525be4",
X"e53f83e0",
X"80085483",
X"e08008ee",
X"38805aff",
X"5f790970",
X"9f2c7b06",
X"5b547a7a",
X"248438ff",
X"1b5af61a",
X"7009709f",
X"2c72067b",
X"ff125a5a",
X"52555580",
X"75259538",
X"7651e4aa",
X"3f83e080",
X"0876ff18",
X"58555773",
X"8024ed38",
X"747f2e86",
X"38a0a83f",
X"745f78ff",
X"1b70585d",
X"58807a25",
X"95387751",
X"e4803f83",
X"e0800876",
X"ff185855",
X"58738024",
X"ed38800b",
X"83e7c00c",
X"800b83e7",
X"e40c80f4",
X"90518d8d",
X"3f81800b",
X"83e7e40c",
X"80f49851",
X"8cff3fa8",
X"0b83e7c0",
X"0c76802e",
X"80e43883",
X"e7c00877",
X"79327030",
X"70720780",
X"2570872b",
X"83e7e40c",
X"51567853",
X"5656e3b7",
X"3f83e080",
X"08802e88",
X"3880f4a0",
X"518cc63f",
X"7651e2f9",
X"3f83e080",
X"085280f5",
X"ac518cb5",
X"3f7651e3",
X"813f83e0",
X"800883e7",
X"c0085557",
X"75742586",
X"38a81656",
X"f7397583",
X"e7c00c86",
X"f07624ff",
X"98388798",
X"0b83e7c0",
X"0c77802e",
X"b1387751",
X"e2b73f83",
X"e0800878",
X"5255e2d7",
X"3f80f4a8",
X"5483e080",
X"088d3887",
X"39807634",
X"81ce3980",
X"f4a45474",
X"53735280",
X"f3f8518b",
X"d43f8054",
X"80f48051",
X"8bcb3f81",
X"145473a8",
X"2e098106",
X"ef38868d",
X"a0519cad",
X"3f805290",
X"3d705257",
X"bffa3f83",
X"527651bf",
X"f33f6281",
X"8f386180",
X"2e80fb38",
X"7b5473ff",
X"2e963878",
X"802e8189",
X"387851e1",
X"dd3f83e0",
X"8008ff15",
X"5559e739",
X"78802e80",
X"f4387851",
X"e1d93f83",
X"e0800880",
X"2efc9038",
X"7851e1a1",
X"3f83e080",
X"085280f3",
X"f45183e3",
X"3f83e080",
X"08a3387c",
X"51859b3f",
X"83e08008",
X"5574ff16",
X"56548074",
X"25ae3874",
X"1d703355",
X"5673af2e",
X"fecf38e9",
X"397851e0",
X"e23f83e0",
X"8008527c",
X"5184d33f",
X"8f397f88",
X"29601005",
X"7a056105",
X"5afc9239",
X"62802efb",
X"d3388052",
X"7651bed4",
X"3fa33d0d",
X"04803d0d",
X"9088b833",
X"7081ff06",
X"70842a81",
X"32708106",
X"51515151",
X"70802e8d",
X"38a80b90",
X"88b834b8",
X"0b9088b8",
X"347083e0",
X"800c823d",
X"0d04803d",
X"0d9088b8",
X"337081ff",
X"0670852a",
X"81327081",
X"06515151",
X"5170802e",
X"8d38980b",
X"9088b834",
X"b80b9088",
X"b8347083",
X"e0800c82",
X"3d0d0493",
X"0b9088bc",
X"34ff0b90",
X"88a83404",
X"ff3d0d02",
X"8f053352",
X"800b9088",
X"bc348a51",
X"99f73fdf",
X"3f80f80b",
X"9088a034",
X"800b9088",
X"8834fa12",
X"52719088",
X"8034800b",
X"90889834",
X"71908890",
X"349088b8",
X"52807234",
X"b8723483",
X"3d0d0480",
X"3d0d028b",
X"05335170",
X"9088b434",
X"febf3f83",
X"e0800880",
X"2ef63882",
X"3d0d0480",
X"3d0d8439",
X"a3ce3ffe",
X"d93f83e0",
X"8008802e",
X"f3389088",
X"b4337081",
X"ff0683e0",
X"800c5182",
X"3d0d0480",
X"3d0da30b",
X"9088bc34",
X"ff0b9088",
X"a8349088",
X"b851a871",
X"34b87134",
X"823d0d04",
X"803d0d90",
X"88bc3370",
X"81c00670",
X"30708025",
X"83e0800c",
X"51515182",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067083",
X"2a813270",
X"81065151",
X"51517080",
X"2ee838b0",
X"0b9088b8",
X"34b80b90",
X"88b83482",
X"3d0d0480",
X"3d0d9080",
X"ac088106",
X"83e0800c",
X"823d0d04",
X"fd3d0d75",
X"77545480",
X"73259438",
X"73708105",
X"55335280",
X"f4ac5187",
X"843fff13",
X"53e93985",
X"3d0d04fd",
X"3d0d7577",
X"53547333",
X"51708938",
X"71335170",
X"802ea138",
X"73337233",
X"52537271",
X"278538ff",
X"51943970",
X"73278538",
X"81518b39",
X"81148113",
X"5354d339",
X"80517083",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"54547233",
X"7081ff06",
X"52527080",
X"2ea33871",
X"81ff0681",
X"14ffbf12",
X"53545270",
X"99268938",
X"a0127081",
X"ff065351",
X"71747081",
X"055634d2",
X"39807434",
X"853d0d04",
X"ffbd3d0d",
X"80c63d08",
X"52a53d70",
X"5254ffb3",
X"3f80c73d",
X"0852853d",
X"705253ff",
X"a63f7252",
X"7351fedf",
X"3f80c53d",
X"0d04fe3d",
X"0d747653",
X"53717081",
X"05533351",
X"70737081",
X"05553470",
X"f038843d",
X"0d04fe3d",
X"0d745280",
X"72335253",
X"70732e8d",
X"38811281",
X"14713353",
X"545270f5",
X"387283e0",
X"800c843d",
X"0d04f63d",
X"0d7c7e60",
X"625a5d5b",
X"56805981",
X"55853974",
X"7a295574",
X"527551b6",
X"fe3f83e0",
X"80087a27",
X"ee387480",
X"2e80dd38",
X"74527551",
X"b6e93f83",
X"e0800875",
X"53765254",
X"b6ed3f83",
X"e080087a",
X"53755256",
X"b6d13f83",
X"e0800879",
X"30707b07",
X"9f2a7077",
X"80240751",
X"51545572",
X"873883e0",
X"8008c538",
X"768118b0",
X"16555858",
X"8974258b",
X"38b71453",
X"7a853880",
X"d7145372",
X"78348119",
X"59ff9f39",
X"8077348c",
X"3d0d04f7",
X"3d0d7b7d",
X"7f620290",
X"05bb0533",
X"5759565a",
X"5ab05872",
X"8338a058",
X"75707081",
X"05523371",
X"59545590",
X"39807425",
X"8e38ff14",
X"77708105",
X"59335454",
X"72ef3873",
X"ff155553",
X"80732589",
X"38775279",
X"51782def",
X"39753375",
X"57537280",
X"2e903872",
X"52795178",
X"2d757081",
X"05573353",
X"ed398b3d",
X"0d04ee3d",
X"0d646669",
X"69707081",
X"0552335b",
X"4a5c5e5e",
X"76802e82",
X"f93876a5",
X"2e098106",
X"82e03880",
X"70416770",
X"70810552",
X"33714a59",
X"575f76b0",
X"2e098106",
X"8c387570",
X"81055733",
X"76485781",
X"5fd01756",
X"75892680",
X"da387667",
X"5c59805c",
X"9339778a",
X"2480c338",
X"7b8a2918",
X"7b708105",
X"5d335a5c",
X"d0197081",
X"ff065858",
X"897727a4",
X"38ff9f19",
X"7081ff06",
X"ffa91b5a",
X"51568576",
X"279238ff",
X"bf197081",
X"ff065156",
X"7585268a",
X"38c91958",
X"778025ff",
X"b9387a47",
X"7b407881",
X"ff065776",
X"80e42e80",
X"e5387680",
X"e424a738",
X"7680d82e",
X"81863876",
X"80d82490",
X"3876802e",
X"81cc3876",
X"a52e81b6",
X"3881b939",
X"7680e32e",
X"818c3881",
X"af397680",
X"f52e9b38",
X"7680f524",
X"8b387680",
X"f32e8181",
X"38819939",
X"7680f82e",
X"80ca3881",
X"8f39913d",
X"70555780",
X"538a5279",
X"841b7108",
X"535b56fc",
X"813f7655",
X"ab397984",
X"1b710894",
X"3d705b5b",
X"525b5675",
X"80258c38",
X"753056ad",
X"78340280",
X"c1055776",
X"5480538a",
X"527551fb",
X"d53f7755",
X"7e54b839",
X"913d7055",
X"7780d832",
X"70307080",
X"25565158",
X"56905279",
X"841b7108",
X"535b57fb",
X"b13f7555",
X"db397984",
X"1b831233",
X"545b5698",
X"3979841b",
X"7108575b",
X"5680547f",
X"537c527d",
X"51fc9c3f",
X"87397652",
X"7d517c2d",
X"66703358",
X"810547fd",
X"8339943d",
X"0d047283",
X"e0940c71",
X"83e0980c",
X"04fb3d0d",
X"883d7070",
X"84055208",
X"57547553",
X"83e09408",
X"5283e098",
X"0851fcc6",
X"3f873d0d",
X"04ff3d0d",
X"73700853",
X"51029305",
X"33723470",
X"08810571",
X"0c833d0d",
X"04fc3d0d",
X"873d8811",
X"557854bd",
X"b95351fc",
X"993f8052",
X"873d51d1",
X"3f863d0d",
X"04fc3d0d",
X"76557483",
X"e398082e",
X"af388053",
X"745187c1",
X"3f83e080",
X"0881ff06",
X"ff147081",
X"ff067230",
X"709f2a51",
X"52555354",
X"72802e84",
X"3871dd38",
X"73fe3874",
X"83e3980c",
X"863d0d04",
X"ff3d0dff",
X"0b83e398",
X"0c84a53f",
X"81518785",
X"3f83e080",
X"0881ff06",
X"5271ee38",
X"81d33f71",
X"83e0800c",
X"833d0d04",
X"fc3d0d76",
X"028405a2",
X"05220288",
X"05a60522",
X"7a545555",
X"55ff823f",
X"72802ea0",
X"3883e3ac",
X"14337570",
X"81055734",
X"81147083",
X"ffff06ff",
X"157083ff",
X"ff065652",
X"5552dd39",
X"800b83e0",
X"800c863d",
X"0d04fc3d",
X"0d76787a",
X"11565355",
X"80537174",
X"2e933872",
X"15517033",
X"83e3ac13",
X"34811281",
X"145452ea",
X"39800b83",
X"e0800c86",
X"3d0d04fd",
X"3d0d9054",
X"83e39808",
X"5186f43f",
X"83e08008",
X"81ff06ff",
X"15713071",
X"30707307",
X"9f2a729f",
X"2a065255",
X"52555372",
X"db38853d",
X"0d04803d",
X"0d83e3a4",
X"081083e3",
X"9c080790",
X"80a80c82",
X"3d0d0480",
X"0b83e3a4",
X"0ce43f04",
X"810b83e3",
X"a40cdb3f",
X"04ed3f04",
X"7183e3a0",
X"0c04803d",
X"0d8051f4",
X"3f810b83",
X"e3a40c81",
X"0b83e39c",
X"0cffbb3f",
X"823d0d04",
X"803d0d72",
X"30707407",
X"802583e3",
X"9c0c51ff",
X"a53f823d",
X"0d04803d",
X"0d028b05",
X"339080a4",
X"0c9080a8",
X"08708106",
X"515170f5",
X"389080a4",
X"087081ff",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d81ff51",
X"d13f83e0",
X"800881ff",
X"0683e080",
X"0c823d0d",
X"04803d0d",
X"73902b73",
X"079080b4",
X"0c823d0d",
X"0404fb3d",
X"0d780284",
X"059f0533",
X"70982b55",
X"57557280",
X"259b3875",
X"80ff0656",
X"805280f7",
X"51e03f83",
X"e0800881",
X"ff065473",
X"812680ff",
X"388051fe",
X"e73fffa2",
X"3f8151fe",
X"df3fff9a",
X"3f7551fe",
X"ed3f7498",
X"2a51fee6",
X"3f74902a",
X"7081ff06",
X"5253feda",
X"3f74882a",
X"7081ff06",
X"5253fece",
X"3f7481ff",
X"0651fec6",
X"3f815575",
X"80c02e09",
X"81068638",
X"8195558d",
X"397580c8",
X"2e098106",
X"84388187",
X"557451fe",
X"a53f8a55",
X"fec83f83",
X"e0800881",
X"ff067098",
X"2b545472",
X"80258c38",
X"ff157081",
X"ff065653",
X"74e23873",
X"83e0800c",
X"873d0d04",
X"fa3d0dfd",
X"c53f8051",
X"fdda3f8a",
X"54fe933f",
X"ff147081",
X"ff065553",
X"73f33873",
X"74535580",
X"c051fea6",
X"3f83e080",
X"0881ff06",
X"5473812e",
X"09810682",
X"9f3883aa",
X"5280c851",
X"fe8c3f83",
X"e0800881",
X"ff065372",
X"812e0981",
X"0681a838",
X"7454873d",
X"74115456",
X"fdc83f83",
X"e0800873",
X"34811470",
X"81ff0655",
X"53837427",
X"e538029a",
X"05335372",
X"812e0981",
X"0681d938",
X"029b0533",
X"5380ce90",
X"547281aa",
X"2e8d3881",
X"c73980e4",
X"518a9e3f",
X"ff145473",
X"802e81b8",
X"38820a52",
X"81e951fd",
X"a53f83e0",
X"800881ff",
X"065372de",
X"38725280",
X"fa51fd92",
X"3f83e080",
X"0881ff06",
X"53728190",
X"38725473",
X"1653fcd6",
X"3f83e080",
X"08733481",
X"147081ff",
X"06555383",
X"7427e838",
X"873d3370",
X"862a7081",
X"06515454",
X"8c557280",
X"e3388455",
X"80de3974",
X"5281e951",
X"fccc3f83",
X"e0800881",
X"ff065382",
X"5581e956",
X"81732786",
X"38735580",
X"c15680ce",
X"90548a39",
X"80e45189",
X"903fff14",
X"5473802e",
X"a9388052",
X"7551fc9a",
X"3f83e080",
X"0881ff06",
X"5372e138",
X"84805280",
X"d051fc86",
X"3f83e080",
X"0881ff06",
X"5372802e",
X"83388055",
X"7483e3a8",
X"348051fb",
X"873ffbc2",
X"3f883d0d",
X"04fb3d0d",
X"7754800b",
X"83e3a833",
X"70832a70",
X"81065155",
X"57557275",
X"2e098106",
X"85387389",
X"2b547352",
X"80d151fb",
X"bd3f83e0",
X"800881ff",
X"065372bd",
X"3882b8c0",
X"54fb833f",
X"83e08008",
X"81ff0653",
X"7281ff2e",
X"09810689",
X"38ff1454",
X"73e7389f",
X"397281fe",
X"2e098106",
X"963883e7",
X"ac5283e3",
X"ac51faed",
X"3ffad33f",
X"fad03f83",
X"39815580",
X"51fa893f",
X"fac43f74",
X"81ff0683",
X"e0800c87",
X"3d0d04fb",
X"3d0d7783",
X"e3ac5654",
X"8151f9ec",
X"3f83e3a8",
X"3370832a",
X"70810651",
X"54567285",
X"3873892b",
X"54735280",
X"d851fab6",
X"3f83e080",
X"0881ff06",
X"537280e4",
X"3881ff51",
X"f9d43f81",
X"fe51f9ce",
X"3f848053",
X"74708105",
X"563351f9",
X"c13fff13",
X"7083ffff",
X"06515372",
X"eb387251",
X"f9b03f72",
X"51f9ab3f",
X"f9d03f83",
X"e080089f",
X"0653a788",
X"5472852e",
X"8c389939",
X"80e45186",
X"c83fff14",
X"54f9b33f",
X"83e08008",
X"81ff2e84",
X"3873e938",
X"8051f8e4",
X"3ff99f3f",
X"800b83e0",
X"800c873d",
X"0d047183",
X"e7b00c88",
X"80800b83",
X"e7ac0c84",
X"80800b83",
X"e7b40c04",
X"fd3d0d77",
X"70175577",
X"05ff1a53",
X"5371ff2e",
X"94387370",
X"81055533",
X"51707370",
X"81055534",
X"ff1252e9",
X"39853d0d",
X"04fc3d0d",
X"87a68155",
X"743383e7",
X"b834a054",
X"83a08053",
X"83e7b008",
X"5283e7ac",
X"0851ffb8",
X"3fa05483",
X"a4805383",
X"e7b00852",
X"83e7ac08",
X"51ffa53f",
X"905483a8",
X"805383e7",
X"b0085283",
X"e7ac0851",
X"ff923fa0",
X"53805283",
X"e7b40883",
X"a0800551",
X"85a03fa0",
X"53805283",
X"e7b40883",
X"a4800551",
X"85903f90",
X"53805283",
X"e7b40883",
X"a8800551",
X"85803fff",
X"753483a0",
X"80548053",
X"83e7b008",
X"5283e7b4",
X"0851fecc",
X"3f80d080",
X"5483b080",
X"5383e7b0",
X"085283e7",
X"b40851fe",
X"b73f86b3",
X"3fa25480",
X"5383e7b4",
X"088c8005",
X"5280f6f0",
X"51fea13f",
X"860b87a8",
X"8334800b",
X"87a88234",
X"800b87a0",
X"9a34af0b",
X"87a09634",
X"bf0b87a0",
X"9734800b",
X"87a09834",
X"9f0b87a0",
X"9934800b",
X"87a09b34",
X"e00b87a8",
X"8934a20b",
X"87a88034",
X"830b87a4",
X"8f34820b",
X"87a88134",
X"863d0d04",
X"fd3d0d83",
X"a0805480",
X"5383e7b4",
X"085283e7",
X"b00851fd",
X"bf3f80d0",
X"805483b0",
X"805383e7",
X"b4085283",
X"e7b00851",
X"fdaa3fa0",
X"5483a080",
X"5383e7b4",
X"085283e7",
X"b00851fd",
X"973fa054",
X"83a48053",
X"83e7b408",
X"5283e7b0",
X"0851fd84",
X"3f905483",
X"a8805383",
X"e7b40852",
X"83e7b008",
X"51fcf13f",
X"83e7b833",
X"87a68134",
X"853d0d04",
X"803d0d90",
X"80900881",
X"0683e080",
X"0c823d0d",
X"04ff3d0d",
X"90809070",
X"0870fe06",
X"7607720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870812c",
X"810683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fd067610",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70822cbf",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"83067682",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870882c",
X"870683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"f1ff0676",
X"882b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087091",
X"2cbf0683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fc87ff",
X"ff067691",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870992c",
X"810683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"ffbf0a06",
X"76992b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80800870",
X"882c8106",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"70892c81",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708a2c",
X"810683e0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708b",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8c2cbf06",
X"83e0800c",
X"51823d0d",
X"04fe3d0d",
X"7481e629",
X"872a9080",
X"a00c843d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"81055434",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727084",
X"05540cff",
X"1151f039",
X"843d0d04",
X"fe3d0d84",
X"80805380",
X"5288800a",
X"51ffb33f",
X"81808053",
X"80528280",
X"0a51c63f",
X"843d0d04",
X"803d0d81",
X"51fcaa3f",
X"72802e90",
X"388051fd",
X"fe3fcd3f",
X"83e7bc33",
X"51fdf43f",
X"8151fcbb",
X"3f8051fc",
X"b63f8051",
X"fc873f82",
X"3d0d04fd",
X"3d0d7552",
X"805480ff",
X"72258838",
X"810bff80",
X"135354ff",
X"bf125170",
X"99268638",
X"e012529e",
X"39ff9f12",
X"51997127",
X"9538d012",
X"e0137054",
X"54518971",
X"2788388f",
X"73278338",
X"80527380",
X"2e853881",
X"80125271",
X"81ff0683",
X"e0800c85",
X"3d0d0480",
X"3d0d84d8",
X"c0518071",
X"70810553",
X"347084e0",
X"c02e0981",
X"06f03882",
X"3d0d04fe",
X"3d0d0297",
X"053351ff",
X"863f83e0",
X"800881ff",
X"0683e7c0",
X"08545280",
X"73249b38",
X"83e7e008",
X"137283e7",
X"e4080753",
X"53717334",
X"83e7c008",
X"810583e7",
X"c00c843d",
X"0d04fa3d",
X"0d82800a",
X"1b558057",
X"883dfc05",
X"54795374",
X"527851ff",
X"bbb83f88",
X"3d0d04fe",
X"3d0d83e7",
X"d8085274",
X"51c29c3f",
X"83e08008",
X"8c387653",
X"755283e7",
X"d80851c6",
X"3f843d0d",
X"04fe3d0d",
X"83e7d808",
X"53755274",
X"51ffbcda",
X"3f83e080",
X"088d3877",
X"53765283",
X"e7d80851",
X"ffa03f84",
X"3d0d04fe",
X"3d0d83e7",
X"d80851ff",
X"bbcd3f83",
X"e0800881",
X"80802e09",
X"81068738",
X"8f808053",
X"9b3983e7",
X"d80851ff",
X"bbb13f83",
X"e0800880",
X"d0802e09",
X"81069238",
X"8fb08053",
X"83e08008",
X"5283e7d8",
X"0851fed6",
X"3f843d0d",
X"04803d0d",
X"fa903f83",
X"e0800884",
X"2980f794",
X"05700883",
X"e0800c51",
X"823d0d04",
X"ed3d0d80",
X"44804380",
X"42804180",
X"705a5bfd",
X"ce3f800b",
X"83e7c00c",
X"800b83e7",
X"e40c80f4",
X"f851ead5",
X"3f81800b",
X"83e7e40c",
X"80f4fc51",
X"eac73f80",
X"d00b83e7",
X"c00c7830",
X"707a0780",
X"2570872b",
X"83e7e40c",
X"5155f981",
X"3f83e080",
X"085280f5",
X"8451eaa1",
X"3f80f80b",
X"83e7c00c",
X"78813270",
X"30707207",
X"80257087",
X"2b83e7e4",
X"0c515656",
X"feef3f83",
X"e0800852",
X"80f59051",
X"e9f73f81",
X"a00b83e7",
X"c00c7882",
X"32703070",
X"72078025",
X"70872b83",
X"e7e40c51",
X"5683e7d8",
X"085256ff",
X"b6d73f83",
X"e0800852",
X"80f59851",
X"e9c73f81",
X"f00b83e7",
X"c00c810b",
X"83e7c45b",
X"5883e7c0",
X"0882197a",
X"32703070",
X"72078025",
X"70872b83",
X"e7e40c51",
X"578e3d70",
X"55ff1b54",
X"57575799",
X"ac3f7970",
X"84055b08",
X"51ffb68d",
X"3f745483",
X"e0800853",
X"775280f5",
X"a051e8f9",
X"3fa81783",
X"e7c00c81",
X"18587785",
X"2e098106",
X"ffaf3883",
X"900b83e7",
X"c00c7887",
X"32703070",
X"72078025",
X"70872b83",
X"e7e40c51",
X"5656f7f7",
X"3f80f5b0",
X"5583e080",
X"08802e8f",
X"3883e7d4",
X"0851ffb5",
X"b83f83e0",
X"80085574",
X"5280f5b8",
X"51e8a63f",
X"83e00b83",
X"e7c00c78",
X"88327030",
X"70720780",
X"2570872b",
X"83e7e40c",
X"515780f5",
X"c45255e8",
X"843f868d",
X"a051f8f1",
X"3f805291",
X"3d705255",
X"9cbe3f83",
X"5274519c",
X"b73f6355",
X"7482fa38",
X"61195978",
X"80258538",
X"74599039",
X"88792585",
X"38885987",
X"39788826",
X"82d93878",
X"822b5580",
X"f3d01508",
X"04f6923f",
X"83e08008",
X"61575575",
X"812e0981",
X"06893883",
X"e0800810",
X"55903975",
X"ff2e0981",
X"06883883",
X"e0800881",
X"2c559075",
X"25853890",
X"55883974",
X"80248338",
X"81557451",
X"f5ec3f82",
X"8e39f5fe",
X"3f83e080",
X"08610555",
X"74802585",
X"38805588",
X"39837525",
X"83388355",
X"7451f5f7",
X"3f81ec39",
X"60873862",
X"802e81e3",
X"3883e38c",
X"0883e388",
X"0cade60b",
X"83e3900c",
X"83e7d808",
X"51d7bd3f",
X"fadd3f81",
X"c6396056",
X"80762598",
X"38ad850b",
X"83e3900c",
X"83e7b815",
X"70085255",
X"d79e3f74",
X"08529239",
X"75802592",
X"3883e7b8",
X"150851ff",
X"b3a13f80",
X"52fd1951",
X"b8396280",
X"2e818c38",
X"83e7b815",
X"700883e7",
X"c408720c",
X"83e7c40c",
X"fd1a7053",
X"51558ba7",
X"3f83e080",
X"08568051",
X"8b9d3f83",
X"e0800852",
X"745187b4",
X"3f755280",
X"5187ad3f",
X"80d53960",
X"55807525",
X"b63883e3",
X"940883e3",
X"880cade6",
X"0b83e390",
X"0c83e7d4",
X"0851d6a8",
X"3f83e7d4",
X"0851d3c8",
X"3f83e080",
X"0881ff06",
X"705255f4",
X"d73f7480",
X"2e9d3881",
X"55a13974",
X"80259438",
X"83e7d408",
X"51ffb293",
X"3f8051f4",
X"bb3f8439",
X"6287387a",
X"802efa83",
X"38805574",
X"83e0800c",
X"953d0d04",
X"fe3d0df4",
X"e73f83e0",
X"8008802e",
X"86388051",
X"818a39f4",
X"ec3f83e0",
X"800880fe",
X"38f58c3f",
X"83e08008",
X"802eb938",
X"8151f2c9",
X"3f8051f4",
X"a23fefbd",
X"3f800b83",
X"e7c00cf9",
X"ab3f83e0",
X"800853ff",
X"0b83e7c0",
X"0cf1a93f",
X"7280cb38",
X"83e7bc33",
X"51f3fc3f",
X"7251f299",
X"3f80c039",
X"f4b43f83",
X"e0800880",
X"2eb53881",
X"51f2863f",
X"8051f3df",
X"3feefa3f",
X"ad850b83",
X"e3900c83",
X"e7c40851",
X"d4da3fff",
X"0b83e7c0",
X"0cf0e53f",
X"83e7c408",
X"52805185",
X"ab3f8151",
X"f5a63f84",
X"3d0d04fc",
X"3d0d800b",
X"83e7bc34",
X"84808052",
X"848a8080",
X"51ffb4cc",
X"3f83e080",
X"0880cd38",
X"88f63f80",
X"f8e851ff",
X"b98b3f83",
X"e0800855",
X"8e808054",
X"80c08053",
X"80f5cc52",
X"83e08008",
X"51f6fa3f",
X"83e7d808",
X"5380f5dc",
X"527451ff",
X"b3d43f83",
X"e0800884",
X"38f7883f",
X"83e7bc33",
X"51f2d03f",
X"8151f4bc",
X"3f92e93f",
X"8151f4b4",
X"3f8151fd",
X"eb3ffa39",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"0280f5e8",
X"0b83e38c",
X"0c80f5ec",
X"0b83e384",
X"0c80f5f0",
X"0b83e394",
X"0c83e08c",
X"08fc050c",
X"800b83e7",
X"c40b83e0",
X"8c08f805",
X"0c83e08c",
X"08f4050c",
X"ffb2a13f",
X"83e08008",
X"8605fc06",
X"83e08c08",
X"f0050c02",
X"83e08c08",
X"f0050831",
X"0d833d70",
X"83e08c08",
X"f8050870",
X"840583e0",
X"8c08f805",
X"0c0c51ff",
X"aee93f83",
X"e08c08f4",
X"05088105",
X"83e08c08",
X"f4050c83",
X"e08c08f4",
X"0508872e",
X"098106ff",
X"ab388484",
X"808051eb",
X"fd3fff0b",
X"83e7c00c",
X"800b83e7",
X"e40c84d8",
X"c00b83e7",
X"e00c8151",
X"efa73f81",
X"51efcc3f",
X"8051efc7",
X"3f8151ef",
X"ed3f8251",
X"f0953f80",
X"51f0bd3f",
X"8051f0e7",
X"3f80d09b",
X"528051e0",
X"e13ffdab",
X"3f83e08c",
X"08fc0508",
X"0d800b83",
X"e0800c87",
X"3d0d83e0",
X"8c0c0480",
X"3d0d81ff",
X"51800b83",
X"e7f01234",
X"ff115170",
X"f438823d",
X"0d04ff3d",
X"0d737033",
X"53518111",
X"33713471",
X"81123483",
X"3d0d04fb",
X"3d0d7779",
X"56568070",
X"71555552",
X"717525ac",
X"38721670",
X"33701470",
X"81ff0655",
X"51515171",
X"74278938",
X"81127081",
X"ff065351",
X"71811470",
X"83ffff06",
X"55525474",
X"7324d638",
X"7183e080",
X"0c873d0d",
X"04fb3d0d",
X"7756d8ab",
X"3f83e080",
X"08802ef6",
X"3883ea8c",
X"08860570",
X"81ff0652",
X"53d6ad3f",
X"810b9088",
X"d4349088",
X"d4337081",
X"ff065153",
X"728b38fa",
X"cb3f8351",
X"f09b3fea",
X"39805574",
X"1675822b",
X"54549088",
X"c0133374",
X"34811555",
X"74852e09",
X"8106e838",
X"810b9088",
X"d4347533",
X"83e7f034",
X"81163383",
X"e7f13482",
X"163383e7",
X"f2348316",
X"3383e7f3",
X"34845283",
X"e7f051fe",
X"ba3f83e0",
X"800881ff",
X"06841733",
X"57537276",
X"2e098106",
X"8c38d6d4",
X"3f83e080",
X"08802e9a",
X"3883ea8c",
X"08a82e09",
X"81068938",
X"860b83ea",
X"8c0c8739",
X"a80b83ea",
X"8c0c80e4",
X"51ef963f",
X"873d0d04",
X"f43d0d7e",
X"60595580",
X"5d807582",
X"2b7183ea",
X"90120c83",
X"eaa4175b",
X"5b577679",
X"3477772e",
X"83b93876",
X"527751ff",
X"adb43f8e",
X"3dfc0554",
X"905383e9",
X"f8527751",
X"ffacef3f",
X"7c567590",
X"2e098106",
X"83953883",
X"e9f851fd",
X"953f83e9",
X"fa51fd8e",
X"3f83e9fc",
X"51fd873f",
X"7683ea88",
X"0c7751ff",
X"aabb3f0b",
X"0b80f488",
X"5283e080",
X"0851ccd3",
X"3f83e080",
X"08812e09",
X"810680d4",
X"387683ea",
X"a00c820b",
X"83e9f834",
X"ff960b83",
X"e9f93477",
X"51ffacff",
X"3f83e080",
X"085583e0",
X"80087725",
X"883883e0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83e9fa34",
X"7483e9fb",
X"347683e9",
X"fc34ff80",
X"0b83e9fd",
X"34819039",
X"83e9f833",
X"83e9f933",
X"71882b07",
X"565b7483",
X"ffff2e09",
X"810680e8",
X"38fe800b",
X"83eaa00c",
X"810b83ea",
X"880cff0b",
X"83e9f834",
X"ff0b83e9",
X"f9347751",
X"ffac8c3f",
X"83e08008",
X"83eaa80c",
X"83e08008",
X"5583e080",
X"08802588",
X"3883e080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"e9fa3474",
X"83e9fb34",
X"7683e9fc",
X"34ff800b",
X"83e9fd34",
X"810b83ea",
X"8734a539",
X"7485962e",
X"09810680",
X"fe387583",
X"eaa00c77",
X"51ffabc0",
X"3f83ea87",
X"3383e080",
X"08075574",
X"83ea8734",
X"83ea8733",
X"81065574",
X"802e8338",
X"845783e9",
X"fc3383e9",
X"fd337188",
X"2b07565c",
X"7481802e",
X"098106a1",
X"3883e9fa",
X"3383e9fb",
X"3371882b",
X"07565bad",
X"80752787",
X"38768207",
X"579c3976",
X"81075796",
X"39748280",
X"2e098106",
X"87387683",
X"07578739",
X"7481ff26",
X"8a387783",
X"ea901b0c",
X"7679348e",
X"3d0d0480",
X"3d0d7284",
X"2983ea90",
X"05700883",
X"e0800c51",
X"823d0d04",
X"fe3d0d80",
X"0b83e9f4",
X"0c800b83",
X"e9f00cff",
X"0b83e7ec",
X"0ca80b83",
X"ea8c0cae",
X"51d0f53f",
X"800b83ea",
X"90545280",
X"73708405",
X"550c8112",
X"5271842e",
X"098106ef",
X"38843d0d",
X"04fe3d0d",
X"74028405",
X"96052253",
X"5371802e",
X"96387270",
X"81055433",
X"51d1803f",
X"ff127083",
X"ffff0651",
X"52e73984",
X"3d0d04fe",
X"3d0d0292",
X"05225382",
X"ac51eaa9",
X"3f80c351",
X"d0dd3f81",
X"9651ea9d",
X"3f725283",
X"e7f051ff",
X"b43f7252",
X"83e7f051",
X"f8f13f83",
X"e0800881",
X"ff0651d0",
X"ba3f843d",
X"0d04ffb1",
X"3d0d80d1",
X"3df80551",
X"f99b3f83",
X"e9f40881",
X"0583e9f4",
X"0c80cf3d",
X"33cf1170",
X"81ff0651",
X"56567483",
X"2688e238",
X"758f06ff",
X"05567583",
X"e7ec082e",
X"9b387583",
X"26963875",
X"83e7ec0c",
X"75842983",
X"ea900570",
X"08535575",
X"51fa993f",
X"80762488",
X"be387584",
X"2983ea90",
X"05557408",
X"802e88af",
X"3883e7ec",
X"08842983",
X"ea900570",
X"08028805",
X"82b90533",
X"525b5574",
X"80d22e84",
X"ac387480",
X"d2249038",
X"74bf2e9c",
X"387480d0",
X"2e81d138",
X"87ee3974",
X"80d32e80",
X"cf387480",
X"d72e81c0",
X"3887dd39",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"055656cf",
X"b63f80c1",
X"51cef03f",
X"f6ed3f86",
X"0b83e7f0",
X"34815283",
X"e7f051d0",
X"933f8151",
X"fde93f74",
X"8938860b",
X"83ea8c0c",
X"8739a80b",
X"83ea8c0c",
X"cf853f80",
X"c151cebf",
X"3ff6bc3f",
X"900b83ea",
X"87338106",
X"56567480",
X"2e833898",
X"5683e9fc",
X"3383e9fd",
X"3371882b",
X"07565974",
X"81802e09",
X"81069c38",
X"83e9fa33",
X"83e9fb33",
X"71882b07",
X"5657ad80",
X"75278c38",
X"75818007",
X"56853975",
X"a0075675",
X"83e7f034",
X"ff0b83e7",
X"f134e00b",
X"83e7f234",
X"800b83e7",
X"f3348452",
X"83e7f051",
X"cf8a3f84",
X"51869b39",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"055659cd",
X"fa3f7951",
X"ffa6913f",
X"83e08008",
X"802e8a38",
X"80ce51cd",
X"a63f85f1",
X"3980c151",
X"cd9d3fce",
X"923fccc7",
X"3f83eaa0",
X"08588375",
X"259b3883",
X"e9fc3383",
X"e9fd3371",
X"882b07fc",
X"1771297a",
X"05838005",
X"5a51578d",
X"39748180",
X"2918ff80",
X"05588180",
X"57805676",
X"762e9238",
X"ccf93f83",
X"e0800883",
X"e7f01734",
X"811656eb",
X"39cce83f",
X"83e08008",
X"81ff0677",
X"5383e7f0",
X"5256f4e7",
X"3f83e080",
X"0881ff06",
X"5575752e",
X"09810681",
X"95389451",
X"e5eb3fcc",
X"e23f80c1",
X"51cc9c3f",
X"cd913f77",
X"527951ff",
X"a4a43f80",
X"5e80d13d",
X"fdf40554",
X"765383e7",
X"f0527951",
X"ffa2b13f",
X"0282b905",
X"33558159",
X"7480d72e",
X"09810680",
X"c5387752",
X"7951ffa3",
X"f53f80d1",
X"3dfdf005",
X"5476538f",
X"3d70537a",
X"5258ffa3",
X"ad3f8056",
X"76762ea2",
X"38751883",
X"e7f01733",
X"71337072",
X"32703070",
X"80257030",
X"7f06811d",
X"5d5f5151",
X"51525b55",
X"db3982ac",
X"51e4e63f",
X"78802e86",
X"3880c351",
X"843980ce",
X"51cb903f",
X"cc853fca",
X"ba3f83d8",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055955",
X"80705d59",
X"80e451e4",
X"b03fcba7",
X"3f80c151",
X"cae13f83",
X"ea880879",
X"2e82d638",
X"83eaa808",
X"80fc0555",
X"80fd5274",
X"5185a03f",
X"83e08008",
X"5b778224",
X"b238ff18",
X"70872b83",
X"ffff8006",
X"80f7b405",
X"83e7f059",
X"57558180",
X"55757081",
X"05573377",
X"70810559",
X"34ff1570",
X"81ff0651",
X"5574ea38",
X"82853977",
X"82e82e81",
X"a3387782",
X"e92e0981",
X"0681aa38",
X"78587787",
X"32703070",
X"72078025",
X"7a8a3270",
X"30707207",
X"80257307",
X"53545a51",
X"57557580",
X"2e973878",
X"78269238",
X"a00b83e7",
X"f01a3481",
X"197081ff",
X"065a55eb",
X"39811870",
X"81ff0659",
X"558a7827",
X"ffbc388f",
X"5883e7eb",
X"183383e7",
X"f01934ff",
X"187081ff",
X"06595577",
X"8426ea38",
X"9058800b",
X"83e7f019",
X"34811870",
X"81ff0670",
X"982b5259",
X"55748025",
X"e93880c6",
X"557a858f",
X"24843880",
X"c2557483",
X"e7f03480",
X"f10b83e7",
X"f334810b",
X"83e7f434",
X"7a83e7f1",
X"347a882c",
X"557483e7",
X"f23480cb",
X"3982f078",
X"2580c438",
X"7780fd29",
X"fd97d305",
X"527951ff",
X"a0d03f80",
X"d13dfdec",
X"055480fd",
X"5383e7f0",
X"527951ff",
X"a0883f7b",
X"81195956",
X"7580fc24",
X"83387858",
X"77882c55",
X"7483e8ed",
X"347783e8",
X"ee347583",
X"e8ef3481",
X"805980cc",
X"3983eaa0",
X"08578378",
X"259b3883",
X"e9fc3383",
X"e9fd3371",
X"882b07fc",
X"1a712979",
X"05838005",
X"5951598d",
X"39778180",
X"2917ff80",
X"05578180",
X"59765279",
X"51ff9fde",
X"3f80d13d",
X"fdec0554",
X"785383e7",
X"f0527951",
X"ff9f973f",
X"7851f6c3",
X"3fc8a83f",
X"c6dd3f8b",
X"3983e9f0",
X"08810583",
X"e9f00c80",
X"d13d0d04",
X"f6e43ffc",
X"39fc3d0d",
X"76787184",
X"2983ea90",
X"05700851",
X"53535370",
X"9e3880ce",
X"723480cf",
X"0b811334",
X"80ce0b82",
X"133480c5",
X"0b831334",
X"70841334",
X"80e73983",
X"eaa41333",
X"5480d272",
X"3473822a",
X"70810651",
X"5180cf53",
X"70843880",
X"d7537281",
X"1334a00b",
X"82133473",
X"83065170",
X"812e9e38",
X"70812488",
X"3870802e",
X"8f389f39",
X"70822e92",
X"3870832e",
X"92389339",
X"80d8558e",
X"3980d355",
X"893980cd",
X"55843980",
X"c4557483",
X"133480c4",
X"0b841334",
X"800b8513",
X"34863d0d",
X"04fc3d0d",
X"76785354",
X"81538055",
X"87397110",
X"73105452",
X"73722651",
X"72802ea7",
X"3870802e",
X"86387180",
X"25e83872",
X"802e9838",
X"71742689",
X"38737231",
X"75740756",
X"5472812a",
X"72812a53",
X"53e53973",
X"51788338",
X"74517083",
X"e0800c86",
X"3d0d04fe",
X"3d0d8053",
X"75527451",
X"ffa33f84",
X"3d0d04fe",
X"3d0d8153",
X"75527451",
X"ff933f84",
X"3d0d04fb",
X"3d0d7779",
X"55558056",
X"74762586",
X"38743055",
X"81567380",
X"25883873",
X"30768132",
X"57548053",
X"73527451",
X"fee73f83",
X"e0800854",
X"75802e87",
X"3883e080",
X"08305473",
X"83e0800c",
X"873d0d04",
X"fa3d0d78",
X"7a575580",
X"57747725",
X"86387430",
X"55815775",
X"9f2c5481",
X"53757432",
X"74315274",
X"51feaa3f",
X"83e08008",
X"5476802e",
X"873883e0",
X"80083054",
X"7383e080",
X"0c883d0d",
X"04fd3d0d",
X"75548074",
X"0c800b84",
X"150c800b",
X"88150c80",
X"0b8c150c",
X"87a68033",
X"7081ff06",
X"5151dd98",
X"3f70812a",
X"81327181",
X"32718106",
X"71810631",
X"84170c53",
X"5370832a",
X"81327182",
X"2a813271",
X"81067181",
X"0631760c",
X"525287a0",
X"90337009",
X"81068816",
X"0c5183e0",
X"8008802e",
X"80c23883",
X"e0800881",
X"2a708106",
X"83e08008",
X"81063184",
X"160c5183",
X"e0800883",
X"2a83e080",
X"08822a71",
X"81067181",
X"0631760c",
X"525283e0",
X"8008842a",
X"81068815",
X"0c83e080",
X"08852a81",
X"068c150c",
X"853d0d04",
X"fe3d0d74",
X"76545271",
X"51fece3f",
X"72812ea2",
X"38817326",
X"8d387282",
X"2ea83872",
X"832e9c38",
X"e6397108",
X"e2388412",
X"08dd3888",
X"1208d838",
X"a5398812",
X"08812e9e",
X"38913988",
X"1208812e",
X"95387108",
X"91388412",
X"088c388c",
X"1208812e",
X"098106ff",
X"b238843d",
X"0d040000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002ad9",
X"00002b1a",
X"00002b3c",
X"00002b62",
X"00002b62",
X"00002b62",
X"00002b62",
X"00002bd3",
X"00002c24",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00003a34",
X"00003a38",
X"00003a40",
X"00003a4c",
X"00003a58",
X"00003a64",
X"00003a70",
X"00003a74",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
