
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f8",
X"e4738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80fb",
X"bc0c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f3",
X"912d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580f1a5",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"96ea0480",
X"3d0d80fd",
X"80087008",
X"810683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d80fd",
X"80087008",
X"70fe0676",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80fd8008",
X"70087081",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80fd8008",
X"700870fd",
X"06761007",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"fd800870",
X"0870822c",
X"bf0683e0",
X"800c5151",
X"823d0d04",
X"ff3d0d80",
X"fd800870",
X"0870fe83",
X"0676822b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80fd8008",
X"70087088",
X"2c870683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80fd8008",
X"700870f1",
X"ff067688",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d80fd80",
X"08700870",
X"8b2cbf06",
X"83e0800c",
X"5151823d",
X"0d04ff3d",
X"0d80fd80",
X"08700870",
X"f88fff06",
X"768b2b07",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"fd900870",
X"0870882c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fd900870",
X"0870892c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fd900870",
X"08708a2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fd900870",
X"08708b2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"fd3d0d75",
X"81e62987",
X"2a80fcf0",
X"0854730c",
X"853d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d848080",
X"53805288",
X"800a51ff",
X"b33f8180",
X"80538052",
X"82800a51",
X"c63f843d",
X"0d04803d",
X"0d8151fc",
X"ce3f7280",
X"2e8338d2",
X"3f8151fc",
X"f03f8051",
X"fceb3f80",
X"51fcb83f",
X"823d0d04",
X"fd3d0d75",
X"52805480",
X"ff722588",
X"38810bff",
X"80135354",
X"ffbf1251",
X"70992686",
X"38e01252",
X"9e39ff9f",
X"12519971",
X"279538d0",
X"12e01370",
X"54545189",
X"71278838",
X"8f732783",
X"38805273",
X"802e8538",
X"81801252",
X"7181ff06",
X"83e0800c",
X"853d0d04",
X"803d0d86",
X"b8c05180",
X"71708105",
X"53347086",
X"c0c02e09",
X"8106f038",
X"823d0d04",
X"fe3d0d02",
X"97053351",
X"ff863f83",
X"e0800881",
X"ff0683e0",
X"9c085452",
X"8073249b",
X"3883e0b8",
X"08137283",
X"e0bc0807",
X"53537173",
X"3483e09c",
X"08810583",
X"e09c0c84",
X"3d0d04fa",
X"3d0d8280",
X"0a1b5580",
X"57883dfc",
X"05547953",
X"74527851",
X"b5963f88",
X"3d0d04fe",
X"3d0d83e0",
X"b0085274",
X"51bbf83f",
X"83e08008",
X"8c387653",
X"755283e0",
X"b00851c7",
X"3f843d0d",
X"04fe3d0d",
X"83e0b008",
X"53755274",
X"51b6b83f",
X"83e08008",
X"8d387753",
X"765283e0",
X"b00851ff",
X"a23f843d",
X"0d04fe3d",
X"0d83e0b4",
X"0851b5ac",
X"3f83e080",
X"08818080",
X"2e098106",
X"883883c1",
X"8080539b",
X"3983e0b4",
X"0851b590",
X"3f83e080",
X"0880d080",
X"2e098106",
X"933883c1",
X"b0805383",
X"e0800852",
X"83e0b408",
X"51fed83f",
X"843d0d04",
X"803d0dfa",
X"cc3f83e0",
X"80088429",
X"80fbc405",
X"700883e0",
X"800c5182",
X"3d0d04ee",
X"3d0d8043",
X"80428041",
X"80705a5b",
X"fdd23f80",
X"0b83e09c",
X"0c800b83",
X"e0bc0c0b",
X"0b80fa80",
X"51affa3f",
X"81800b83",
X"e0bc0c0b",
X"0b80fa84",
X"51afea3f",
X"80d00b83",
X"e09c0c78",
X"30707a07",
X"80257087",
X"2b83e0bc",
X"0c5155f9",
X"b73f83e0",
X"8008520b",
X"0b80fa8c",
X"51afc23f",
X"80f80b83",
X"e09c0c78",
X"81327030",
X"70720780",
X"2570872b",
X"83e0bc0c",
X"515656fe",
X"eb3f83e0",
X"8008520b",
X"0b80fa98",
X"51af963f",
X"81a00b83",
X"e09c0c78",
X"82327030",
X"70720780",
X"2570872b",
X"83e0bc0c",
X"515683e0",
X"b4085256",
X"b0b13f83",
X"e0800852",
X"0b0b80fa",
X"a051aee5",
X"3f81f00b",
X"83e09c0c",
X"810b83e0",
X"a05b5883",
X"e09c0882",
X"197a3270",
X"30707207",
X"80257087",
X"2b83e0bc",
X"0c51578e",
X"3d7055ff",
X"1b545757",
X"57a4c33f",
X"79708405",
X"5b0851af",
X"e63f7454",
X"83e08008",
X"5377520b",
X"0b80faa8",
X"51ae963f",
X"a81783e0",
X"9c0c8118",
X"5877852e",
X"098106ff",
X"ae388390",
X"0b83e09c",
X"0c788732",
X"70307072",
X"07802570",
X"872b83e0",
X"bc0c5156",
X"0b0b80fa",
X"b85256ad",
X"e03f83e0",
X"0b83e09c",
X"0c788832",
X"70307072",
X"07802570",
X"872b83e0",
X"bc0c5156",
X"0b0b80fa",
X"cc5256ad",
X"bc3f868d",
X"a051f990",
X"3f805291",
X"3d705255",
X"8ba53f83",
X"5274518b",
X"9e3f6119",
X"59788025",
X"85388059",
X"90398879",
X"25853888",
X"59873978",
X"882682ae",
X"3878822b",
X"5580f8f4",
X"150804f6",
X"e33f83e0",
X"80086157",
X"5575812e",
X"09810689",
X"3883e080",
X"08105590",
X"3975ff2e",
X"09810688",
X"3883e080",
X"08812c55",
X"90752585",
X"38905588",
X"39748024",
X"83388155",
X"7451f6c0",
X"3f81e339",
X"f6d33f83",
X"e0800861",
X"05557480",
X"25853880",
X"55883987",
X"75258338",
X"87557451",
X"f6cf3f81",
X"c1396087",
X"3862802e",
X"81b838a0",
X"990b83e0",
X"d00c83e0",
X"b408518c",
X"a93ffafe",
X"3f81a339",
X"60568076",
X"2598389f",
X"b80b83e0",
X"d00c83e0",
X"94157008",
X"52558c8a",
X"3f740852",
X"91397580",
X"25913883",
X"e0941508",
X"51ada23f",
X"8052fd19",
X"51b83962",
X"802e80ea",
X"3883e094",
X"15700883",
X"e0a00872",
X"0c83e0a0",
X"0cfd1a70",
X"53515596",
X"f93f83e0",
X"80085680",
X"5196ef3f",
X"83e08008",
X"52745193",
X"8e3f7552",
X"80519387",
X"3fb43962",
X"802eaf38",
X"a0990b83",
X"e0d00c83",
X"e0b00851",
X"8ba03f83",
X"e0b00851",
X"acb13f9c",
X"800a5380",
X"c0805283",
X"e0800851",
X"f9993f81",
X"558c3962",
X"87387a80",
X"2efac538",
X"80557483",
X"e0800c94",
X"3d0d04fe",
X"3d0df5c0",
X"3f83e080",
X"08802e86",
X"38805180",
X"f639f5c8",
X"3f83e080",
X"0880ea38",
X"f5ee3f83",
X"e0800880",
X"2eaa3881",
X"51f3c03f",
X"839b3f80",
X"0b83e09c",
X"0cf9f43f",
X"83e08008",
X"53ff0b83",
X"e09c0c85",
X"ee3f72bd",
X"387251f3",
X"9e3fbb39",
X"f5a23f83",
X"e0800880",
X"2eb03881",
X"51f38c3f",
X"82e73f9f",
X"b80b83e0",
X"d00c83e0",
X"a0085189",
X"fd3fff0b",
X"83e09c0c",
X"85b93f83",
X"e0a00852",
X"805191bb",
X"3f8151f6",
X"8d3f843d",
X"0d0483e0",
X"8c080283",
X"e08c0cfa",
X"3d0d800b",
X"83e0a00b",
X"83e08c08",
X"fc050c83",
X"e08c08f8",
X"050caded",
X"3f83e080",
X"088605fc",
X"0683e08c",
X"08f4050c",
X"0283e08c",
X"08f40508",
X"310d853d",
X"7083e08c",
X"08fc0508",
X"70840583",
X"e08c08fc",
X"050c0c51",
X"aab73f83",
X"e08c08f8",
X"05088105",
X"83e08c08",
X"f8050c83",
X"e08c08f8",
X"0508862e",
X"098106ff",
X"ad388688",
X"80805181",
X"aa3fff0b",
X"83e09c0c",
X"800b83e0",
X"bc0c86b8",
X"c00b83e0",
X"b80c8151",
X"f1c93f81",
X"51f1f23f",
X"8051f1ed",
X"3f8151f2",
X"973f8151",
X"f2f43f82",
X"51f2be3f",
X"8e845280",
X"51a7fb3f",
X"84808052",
X"86848080",
X"51add63f",
X"83e08008",
X"80d33893",
X"d23f80fe",
X"c851b295",
X"3f83e080",
X"0883e0b4",
X"08540b0b",
X"80fad453",
X"83e08008",
X"5283e08c",
X"08f4050c",
X"ace93f83",
X"e0800884",
X"38f6bf3f",
X"9c800a54",
X"80c08053",
X"0b0b80fa",
X"e05283e0",
X"8c08f405",
X"0851f681",
X"3f8151f3",
X"f13f9daa",
X"3f8151f3",
X"e93ffccf",
X"3ffc3971",
X"83e0c40c",
X"8880800b",
X"83e0c00c",
X"8480800b",
X"83e0c80c",
X"04f03d0d",
X"80fbf808",
X"54733383",
X"e0cc3483",
X"a0805683",
X"e0c40816",
X"83e0c008",
X"17565474",
X"33743483",
X"e0c80816",
X"54807434",
X"81165675",
X"83a0a02e",
X"098106db",
X"3883a480",
X"5683e0c4",
X"081683e0",
X"c0081756",
X"54743374",
X"3483e0c8",
X"08165480",
X"74348116",
X"567583a4",
X"a02e0981",
X"06db3883",
X"a8805683",
X"e0c40816",
X"83e0c008",
X"17565474",
X"33743483",
X"e0c80816",
X"54807434",
X"81165675",
X"83a8902e",
X"098106db",
X"3880fbf8",
X"0854ff74",
X"34805683",
X"e0c40816",
X"83e0c808",
X"17555573",
X"33753481",
X"16567583",
X"a0802e09",
X"8106e438",
X"83b08056",
X"83e0c408",
X"1683e0c8",
X"08175555",
X"73337534",
X"81165675",
X"8480802e",
X"098106e4",
X"38f2ed3f",
X"893d58a2",
X"5380f998",
X"52775180",
X"dcbc3f80",
X"578c8056",
X"83e0c808",
X"16771955",
X"55733375",
X"34811681",
X"18585676",
X"a22e0981",
X"06e63880",
X"fc9c0854",
X"86743480",
X"fca00854",
X"80743480",
X"fc980854",
X"80743480",
X"fc880854",
X"af743480",
X"fc940854",
X"bf743480",
X"fc900854",
X"80743480",
X"fc8c0854",
X"9f743480",
X"fc840854",
X"80743480",
X"fbf00854",
X"e0743480",
X"fbe80854",
X"76743480",
X"fbe40854",
X"83743480",
X"fbec0854",
X"82743492",
X"3d0d04fe",
X"3d0d8053",
X"83e0c808",
X"1383e0c4",
X"08145252",
X"70337234",
X"81135372",
X"83a0802e",
X"098106e4",
X"3883b080",
X"5383e0c8",
X"081383e0",
X"c4081452",
X"52703372",
X"34811353",
X"72848080",
X"2e098106",
X"e43883a0",
X"805383e0",
X"c8081383",
X"e0c40814",
X"52527033",
X"72348113",
X"537283a0",
X"a02e0981",
X"06e43883",
X"a4805383",
X"e0c80813",
X"83e0c408",
X"14525270",
X"33723481",
X"13537283",
X"a4a02e09",
X"8106e438",
X"83a88053",
X"83e0c808",
X"1383e0c4",
X"08145252",
X"70337234",
X"81135372",
X"83a8902e",
X"098106e4",
X"3880fbf8",
X"085183e0",
X"cc337134",
X"843d0d04",
X"fd3d0d75",
X"5480740c",
X"800b8415",
X"0c800b88",
X"150c80fb",
X"fc087033",
X"7081ff06",
X"70812a81",
X"32718132",
X"71810671",
X"81063184",
X"1a0c5656",
X"70832a81",
X"3271822a",
X"81327181",
X"06718106",
X"31790c52",
X"55515151",
X"80fbf408",
X"70337009",
X"81068817",
X"0c515185",
X"3d0d04fe",
X"3d0d7476",
X"54527151",
X"ff9a3f72",
X"812ea238",
X"8173268d",
X"3872822e",
X"ab387283",
X"2e9f38e6",
X"397108e2",
X"38841208",
X"dd388812",
X"08d838a0",
X"39881208",
X"812e0981",
X"06cc3894",
X"39881208",
X"812e8d38",
X"71088938",
X"84120880",
X"2effb738",
X"843d0d04",
X"fc3d0d76",
X"70525580",
X"c7933f83",
X"e0800815",
X"ff055473",
X"752e8e38",
X"73335372",
X"ae2e8638",
X"ff1454ef",
X"39775281",
X"145180c6",
X"aa3f83e0",
X"80083070",
X"83e08008",
X"07802583",
X"e0800c53",
X"863d0d04",
X"fc3d0d76",
X"705255ab",
X"fe3f83e0",
X"80085481",
X"5383e080",
X"0880c138",
X"7451abc1",
X"3f83e080",
X"0880fb80",
X"5383e080",
X"085253ff",
X"8f3f83e0",
X"8008a138",
X"80fb8452",
X"7251ff80",
X"3f83e080",
X"08923880",
X"fb885272",
X"51fef13f",
X"83e08008",
X"802e8338",
X"81547353",
X"7283e080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"ab9d3f81",
X"5383e080",
X"08973873",
X"51aae63f",
X"80fb8c52",
X"83e08008",
X"51feb93f",
X"83e08008",
X"537283e0",
X"800c853d",
X"0d04e03d",
X"0da33d08",
X"70525ea1",
X"8e3f83e0",
X"80083394",
X"3d565473",
X"943880fe",
X"e0527451",
X"84d0397d",
X"527851a4",
X"903f84db",
X"397d51a0",
X"f63f83e0",
X"80085274",
X"51a0a63f",
X"83e0d008",
X"52933d70",
X"525ba780",
X"3f83e080",
X"0859800b",
X"83e08008",
X"555c83e0",
X"80087c2e",
X"9438811c",
X"74525caa",
X"813f83e0",
X"80085483",
X"e08008ee",
X"38805aff",
X"7a437a42",
X"7a415f79",
X"09709f2c",
X"7b065b54",
X"7b7a2484",
X"38ff1c5a",
X"f61a7009",
X"709f2c72",
X"067bff12",
X"5a5a5255",
X"55807525",
X"95387651",
X"a9c03f83",
X"e0800876",
X"ff185855",
X"57738024",
X"ed38747f",
X"2e8638eb",
X"e33f745f",
X"78ff1b70",
X"585e5880",
X"7a259538",
X"7751a996",
X"3f83e080",
X"0876ff18",
X"58555873",
X"8024ed38",
X"800b83e0",
X"9c0c800b",
X"83e0bc0c",
X"80fb9051",
X"9deb3f81",
X"800b83e0",
X"bc0c80fb",
X"98519ddd",
X"3fa80b83",
X"e09c0c76",
X"802e80e4",
X"3883e09c",
X"08777932",
X"70307072",
X"07802570",
X"872b83e0",
X"bc0c5156",
X"78535656",
X"a8cd3f83",
X"e0800880",
X"2e883880",
X"fba0519d",
X"a43f7651",
X"a88f3f83",
X"e0800852",
X"80fab451",
X"9d933f76",
X"51a8973f",
X"83e08008",
X"83e09c08",
X"55577574",
X"258638a8",
X"1656f739",
X"7583e09c",
X"0c86f076",
X"24ff9838",
X"87980b83",
X"e09c0c77",
X"802eb138",
X"7751a7cd",
X"3f83e080",
X"08785255",
X"a7ed3f80",
X"fba85483",
X"e080088d",
X"38873980",
X"7634fda0",
X"3980fba4",
X"54745373",
X"5280faf0",
X"519cb23f",
X"805480fb",
X"b0519ca9",
X"3f811454",
X"73a82e09",
X"8106ef38",
X"868da051",
X"e7f23f80",
X"52903d70",
X"5254fa87",
X"3f835273",
X"51fa803f",
X"61802e81",
X"9c387c54",
X"73ff2e96",
X"3878802e",
X"819d3878",
X"51a6f73f",
X"83e08008",
X"ff155559",
X"e7397880",
X"2e818838",
X"7851a6f3",
X"3f83e080",
X"08802efc",
X"96387851",
X"a6bb3f83",
X"e0800883",
X"e0800853",
X"80faf852",
X"54bfe33f",
X"83e08008",
X"a5387a51",
X"80c19a3f",
X"83e08008",
X"5574ff16",
X"56548074",
X"25fbfd38",
X"741b7033",
X"555673af",
X"2efecc38",
X"e8397a51",
X"80c0f63f",
X"825380fa",
X"fc5283e0",
X"80081b51",
X"80d29b3f",
X"7a5180c0",
X"e03f7352",
X"83e08008",
X"1b5180c0",
X"b83ffbc4",
X"397f8829",
X"6010057a",
X"0561055a",
X"fbf539a2",
X"3d0d0480",
X"3d0d81ff",
X"51800b83",
X"e0dc1234",
X"ff115170",
X"f438823d",
X"0d04ff3d",
X"0d737033",
X"53518111",
X"33713471",
X"81123483",
X"3d0d04fb",
X"3d0d7779",
X"56568070",
X"71555552",
X"717525ac",
X"38721670",
X"33701470",
X"81ff0655",
X"51515171",
X"74278938",
X"81127081",
X"ff065351",
X"71811470",
X"83ffff06",
X"55525474",
X"7324d638",
X"7183e080",
X"0c873d0d",
X"04fd3d0d",
X"7554948f",
X"3f83e080",
X"08802ef6",
X"3883e2f8",
X"08860570",
X"81ff0652",
X"5391e83f",
X"8439eef3",
X"3f93f03f",
X"83e08008",
X"812ef338",
X"92cb3f83",
X"e0800874",
X"3492c23f",
X"83e08008",
X"81153492",
X"b83f83e0",
X"80088215",
X"3492ae3f",
X"83e08008",
X"83153492",
X"a43f83e0",
X"80088415",
X"348439ee",
X"b23f93af",
X"3f83e080",
X"08802ef3",
X"38733383",
X"e0dc3481",
X"143383e0",
X"dd348214",
X"3383e0de",
X"34831433",
X"83e0df34",
X"845283e0",
X"dc51fea7",
X"3f83e080",
X"0881ff06",
X"84153355",
X"5372742e",
X"0981068c",
X"3892a03f",
X"83e08008",
X"802e9a38",
X"83e2f808",
X"a82e0981",
X"06893886",
X"0b83e2f8",
X"0c8739a8",
X"0b83e2f8",
X"0c80e451",
X"e3ea3f85",
X"3d0d04f4",
X"3d0d7e60",
X"5955805d",
X"8075822b",
X"7183e2fc",
X"120c83e3",
X"90175b5b",
X"57767934",
X"77772e83",
X"b1387652",
X"77519be1",
X"3f8e3dfc",
X"05549053",
X"83e2e452",
X"77519b98",
X"3f7c5675",
X"902e0981",
X"06838f38",
X"83e2e451",
X"fd843f83",
X"e2e651fc",
X"fd3f83e2",
X"e851fcf6",
X"3f7683e2",
X"f40c7751",
X"98e53f80",
X"fb845283",
X"e0800851",
X"f5ea3f83",
X"e0800881",
X"2e098106",
X"80d33876",
X"83e38c0c",
X"820b83e2",
X"e434ff96",
X"0b83e2e5",
X"3477519b",
X"ab3f83e0",
X"80085583",
X"e0800877",
X"25883883",
X"e080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583e2e6",
X"347483e2",
X"e7347683",
X"e2e834ff",
X"800b83e2",
X"e934818f",
X"3983e2e4",
X"3383e2e5",
X"3371882b",
X"07565b74",
X"83ffff2e",
X"09810680",
X"e738fe80",
X"0b83e38c",
X"0c810b83",
X"e2f40cff",
X"0b83e2e4",
X"34ff0b83",
X"e2e53477",
X"519ab93f",
X"83e08008",
X"83e3940c",
X"83e08008",
X"5583e080",
X"08802588",
X"3883e080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"e2e63474",
X"83e2e734",
X"7683e2e8",
X"34ff800b",
X"83e2e934",
X"810b83e2",
X"f334a439",
X"7485962e",
X"09810680",
X"fd387583",
X"e38c0c77",
X"5199ee3f",
X"83e2f333",
X"83e08008",
X"07557483",
X"e2f33483",
X"e2f33381",
X"06557480",
X"2e833884",
X"5783e2e8",
X"3383e2e9",
X"3371882b",
X"07565c74",
X"81802e09",
X"8106a138",
X"83e2e633",
X"83e2e733",
X"71882b07",
X"565bad80",
X"75278738",
X"76820757",
X"9c397681",
X"07579639",
X"7482802e",
X"09810687",
X"38768307",
X"57873974",
X"81ff268a",
X"387783e2",
X"fc1b0c76",
X"79348e3d",
X"0d04803d",
X"0d728429",
X"83e2fc05",
X"700883e0",
X"800c5182",
X"3d0d04fe",
X"3d0d800b",
X"83e2e00c",
X"800b83e2",
X"dc0cff0b",
X"83e0d80c",
X"a80b83e2",
X"f80cae51",
X"8ca53f80",
X"0b83e2fc",
X"54528073",
X"70840555",
X"0c811252",
X"71842e09",
X"8106ef38",
X"843d0d04",
X"fe3d0d74",
X"02840596",
X"05225353",
X"71802e96",
X"38727081",
X"05543351",
X"8cc43fff",
X"127083ff",
X"ff065152",
X"e739843d",
X"0d04fe3d",
X"0d029205",
X"225382ac",
X"51df853f",
X"80c3518c",
X"a13f8196",
X"51def93f",
X"725283e0",
X"dc51ffb4",
X"3f725283",
X"e0dc51f8",
X"e63f83e0",
X"800881ff",
X"06518bfe",
X"3f843d0d",
X"04ffb13d",
X"0d80d13d",
X"f80551f9",
X"903f83e2",
X"e0088105",
X"83e2e00c",
X"80cf3d33",
X"cf117081",
X"ff065156",
X"56748326",
X"88cd3875",
X"8f06ff05",
X"567583e0",
X"d8082e9b",
X"38758326",
X"96387583",
X"e0d80c75",
X"842983e2",
X"fc057008",
X"53557551",
X"faa13f80",
X"762488a9",
X"38758429",
X"83e2fc05",
X"55740880",
X"2e889a38",
X"83e0d808",
X"842983e2",
X"fc057008",
X"02880582",
X"b9053352",
X"5b557480",
X"d22e849a",
X"387480d2",
X"24903874",
X"bf2e9c38",
X"7480d02e",
X"81d13887",
X"d9397480",
X"d32e80cf",
X"387480d7",
X"2e81c038",
X"87c83902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"56568b80",
X"3f80c151",
X"8ab43ff6",
X"e23f860b",
X"83e0dc34",
X"815283e0",
X"dc518bef",
X"3f8151fd",
X"e93f7489",
X"38860b83",
X"e2f80c87",
X"39a80b83",
X"e2f80c8a",
X"cf3f80c1",
X"518a833f",
X"f6b13f90",
X"0b83e2f3",
X"33810656",
X"5674802e",
X"83389856",
X"83e2e833",
X"83e2e933",
X"71882b07",
X"56597481",
X"802e0981",
X"069c3883",
X"e2e63383",
X"e2e73371",
X"882b0756",
X"57ad8075",
X"278c3875",
X"81800756",
X"853975a0",
X"07567583",
X"e0dc34ff",
X"0b83e0dd",
X"34e00b83",
X"e0de3480",
X"0b83e0df",
X"34845283",
X"e0dc518a",
X"e63f8451",
X"86863902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"565989c4",
X"3f795194",
X"c03f83e0",
X"8008802e",
X"8a3880ce",
X"5188eb3f",
X"85dd3980",
X"c15188e2",
X"3f89ea3f",
X"87ee3f83",
X"e38c0858",
X"8375259b",
X"3883e2e8",
X"3383e2e9",
X"3371882b",
X"07fc1771",
X"297a0583",
X"80055a51",
X"578d3974",
X"81802918",
X"ff800558",
X"81805780",
X"5676762e",
X"923888c1",
X"3f83e080",
X"0883e0dc",
X"17348116",
X"56eb3988",
X"b03f83e0",
X"800881ff",
X"06775383",
X"e0dc5256",
X"f4dd3f83",
X"e0800881",
X"ff065575",
X"752e0981",
X"06818438",
X"88b23f80",
X"c15187e6",
X"3f88ee3f",
X"77527951",
X"92df3f80",
X"5e80d13d",
X"fdf40554",
X"765383e0",
X"dc527951",
X"90e83f02",
X"82b90533",
X"55815874",
X"80d72e09",
X"8106bc38",
X"80d13dfd",
X"f0055476",
X"538f3d70",
X"537a5259",
X"91ee3f80",
X"5676762e",
X"a2387519",
X"83e0dc17",
X"33713370",
X"72327030",
X"70802570",
X"307e0681",
X"1d5d5e51",
X"5151525b",
X"55db3982",
X"ac51d9d4",
X"3f77802e",
X"863880c3",
X"51843980",
X"ce5186e6",
X"3f87ee3f",
X"85f23f83",
X"d5390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290559",
X"5580705d",
X"5987893f",
X"80c15186",
X"bd3f83e2",
X"f408792e",
X"82db3883",
X"e3940880",
X"fc055580",
X"fd527451",
X"bdc13f83",
X"e080085b",
X"778224b2",
X"38ff1870",
X"872b83ff",
X"ff800680",
X"fd940583",
X"e0dc5957",
X"55818055",
X"75708105",
X"57337770",
X"81055934",
X"ff157081",
X"ff065155",
X"74ea3882",
X"8a397782",
X"e82e81aa",
X"387782e9",
X"2e098106",
X"81b13880",
X"fbac518c",
X"d43f7858",
X"77873270",
X"30707207",
X"80257a8a",
X"32703070",
X"72078025",
X"73075354",
X"5a515755",
X"75802e97",
X"38787826",
X"9238a00b",
X"83e0dc1a",
X"34811970",
X"81ff065a",
X"55eb3981",
X"187081ff",
X"0659558a",
X"7827ffbc",
X"388f5883",
X"e0d71833",
X"83e0dc19",
X"34ff1870",
X"81ff0659",
X"55778426",
X"ea389058",
X"800b83e0",
X"dc193481",
X"187081ff",
X"0670982b",
X"52595574",
X"8025e938",
X"80c6557a",
X"858f2484",
X"3880c255",
X"7483e0dc",
X"3480f10b",
X"83e0df34",
X"810b83e0",
X"e0347a83",
X"e0dd347a",
X"882c5574",
X"83e0de34",
X"80c93982",
X"f0782580",
X"c2387780",
X"fd29fd97",
X"d3055279",
X"518f963f",
X"80d13dfd",
X"ec055480",
X"fd5383e0",
X"dc527951",
X"8eca3f7b",
X"81195956",
X"7580fc24",
X"83387858",
X"77882c55",
X"7483e1d9",
X"347783e1",
X"da347583",
X"e1db3481",
X"805980ca",
X"3983e38c",
X"08578378",
X"259b3883",
X"e2e83383",
X"e2e93371",
X"882b07fc",
X"1a712979",
X"05838005",
X"5951598d",
X"39778180",
X"2917ff80",
X"05578180",
X"59765279",
X"518ea63f",
X"80d13dfd",
X"ec055478",
X"5383e0dc",
X"5279518d",
X"db3f7851",
X"f6d83f84",
X"943f8298",
X"3f8b3983",
X"e2dc0881",
X"0583e2dc",
X"0c80d13d",
X"0d04f6f9",
X"3fdfa83f",
X"f939fc3d",
X"0d767871",
X"842983e2",
X"fc057008",
X"51535353",
X"709e3880",
X"ce723480",
X"cf0b8113",
X"3480ce0b",
X"82133480",
X"c50b8313",
X"34708413",
X"3480e739",
X"83e39013",
X"335480d2",
X"72347382",
X"2a708106",
X"515180cf",
X"53708438",
X"80d75372",
X"811334a0",
X"0b821334",
X"73830651",
X"70812e9e",
X"38708124",
X"88387080",
X"2e8f389f",
X"3970822e",
X"92387083",
X"2e923893",
X"3980d855",
X"8e3980d3",
X"55893980",
X"cd558439",
X"80c45574",
X"83133480",
X"c40b8413",
X"34800b85",
X"1334863d",
X"0d04fe3d",
X"0d80fcac",
X"08703370",
X"81ff0670",
X"842a8132",
X"81065551",
X"52537180",
X"2e8c38a8",
X"733480fc",
X"ac0851b8",
X"71347183",
X"e0800c84",
X"3d0d04fe",
X"3d0d80fc",
X"ac087033",
X"7081ff06",
X"70852a81",
X"32810655",
X"51525371",
X"802e8c38",
X"98733480",
X"fcac0851",
X"b8713471",
X"83e0800c",
X"843d0d04",
X"803d0d80",
X"fca80851",
X"93713480",
X"fcb40851",
X"ff713482",
X"3d0d04fe",
X"3d0d0293",
X"053380fc",
X"a8085353",
X"8072348a",
X"51d3a13f",
X"d33f80fc",
X"b8085280",
X"f8723480",
X"fcd00852",
X"807234fa",
X"1380fcd8",
X"08535372",
X"723480fc",
X"c0085280",
X"723480fc",
X"c8085272",
X"723480fc",
X"ac085280",
X"723480fc",
X"ac0852b8",
X"7234843d",
X"0d04ff3d",
X"0d028f05",
X"3380fcb0",
X"08525271",
X"7134fe9e",
X"3f83e080",
X"08802ef6",
X"38833d0d",
X"04803d0d",
X"8439dc93",
X"3ffeb83f",
X"83e08008",
X"802ef338",
X"80fcb008",
X"70337081",
X"ff0683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fca80851",
X"a3713480",
X"fcb40851",
X"ff713480",
X"fcac0851",
X"a8713480",
X"fcac0851",
X"b8713482",
X"3d0d0480",
X"3d0d80fc",
X"a8087033",
X"7081c006",
X"70307080",
X"2583e080",
X"0c515151",
X"51823d0d",
X"04ff3d0d",
X"80fcac08",
X"70337081",
X"ff067083",
X"2a813270",
X"81065151",
X"51525270",
X"802ee538",
X"b0723480",
X"fcac0851",
X"b8713483",
X"3d0d0480",
X"3d0d80fc",
X"e4087008",
X"810683e0",
X"800c5182",
X"3d0d04fd",
X"3d0d7577",
X"54548073",
X"25943873",
X"70810555",
X"335280fb",
X"b451859d",
X"3fff1353",
X"e939853d",
X"0d04f63d",
X"0d7c7e60",
X"625a5d5b",
X"56805981",
X"55853974",
X"7a295574",
X"527551b5",
X"923f83e0",
X"80087a27",
X"ee387480",
X"2e80dd38",
X"74527551",
X"b4fd3f83",
X"e0800875",
X"53765254",
X"b5a43f83",
X"e080087a",
X"53755256",
X"b4e53f83",
X"e0800879",
X"30707b07",
X"9f2a7077",
X"80240751",
X"51545572",
X"873883e0",
X"8008c538",
X"768118b0",
X"16555858",
X"8974258b",
X"38b71453",
X"7a853880",
X"d7145372",
X"78348119",
X"59ff9f39",
X"8077348c",
X"3d0d04f7",
X"3d0d7b7d",
X"7f620290",
X"05bb0533",
X"5759565a",
X"5ab05872",
X"8338a058",
X"75707081",
X"05523371",
X"59545590",
X"39807425",
X"8e38ff14",
X"77708105",
X"59335454",
X"72ef3873",
X"ff155553",
X"80732589",
X"38775279",
X"51782def",
X"39753375",
X"57537280",
X"2e903872",
X"52795178",
X"2d757081",
X"05573353",
X"ed398b3d",
X"0d04ee3d",
X"0d646669",
X"69707081",
X"0552335b",
X"4a5c5e5e",
X"76802e82",
X"f93876a5",
X"2e098106",
X"82e03880",
X"70416770",
X"70810552",
X"33714a59",
X"575f76b0",
X"2e098106",
X"8c387570",
X"81055733",
X"76485781",
X"5fd01756",
X"75892680",
X"da387667",
X"5c59805c",
X"9339778a",
X"2480c338",
X"7b8a2918",
X"7b708105",
X"5d335a5c",
X"d0197081",
X"ff065858",
X"897727a4",
X"38ff9f19",
X"7081ff06",
X"ffa91b5a",
X"51568576",
X"279238ff",
X"bf197081",
X"ff065156",
X"7585268a",
X"38c91958",
X"778025ff",
X"b9387a47",
X"7b407881",
X"ff065776",
X"80e42e80",
X"e5387680",
X"e424a738",
X"7680d82e",
X"81863876",
X"80d82490",
X"3876802e",
X"81cc3876",
X"a52e81b6",
X"3881b939",
X"7680e32e",
X"818c3881",
X"af397680",
X"f52e9b38",
X"7680f524",
X"8b387680",
X"f32e8181",
X"38819939",
X"7680f82e",
X"80ca3881",
X"8f39913d",
X"70555780",
X"538a5279",
X"841b7108",
X"535b56fc",
X"813f7655",
X"ab397984",
X"1b710894",
X"3d705b5b",
X"525b5675",
X"80258c38",
X"753056ad",
X"78340280",
X"c1055776",
X"5480538a",
X"527551fb",
X"d53f7755",
X"7e54b839",
X"913d7055",
X"7780d832",
X"70307080",
X"25565158",
X"56905279",
X"841b7108",
X"535b57fb",
X"b13f7555",
X"db397984",
X"1b831233",
X"545b5698",
X"3979841b",
X"7108575b",
X"5680547f",
X"537c527d",
X"51fc9c3f",
X"87397652",
X"7d517c2d",
X"66703358",
X"810547fd",
X"8339943d",
X"0d047283",
X"e0900c71",
X"83e0940c",
X"04fb3d0d",
X"883d7070",
X"84055208",
X"57547553",
X"83e09008",
X"5283e094",
X"0851fcc6",
X"3f873d0d",
X"04ff3d0d",
X"73700853",
X"51029305",
X"33723470",
X"08810571",
X"0c833d0d",
X"04fc3d0d",
X"873d8811",
X"55785480",
X"c0c55351",
X"fc983f80",
X"52873d51",
X"d03f863d",
X"0d04fd3d",
X"0d757052",
X"54a58e3f",
X"83e08008",
X"14537274",
X"2e9238ff",
X"13703353",
X"5371af2e",
X"098106ee",
X"38811353",
X"7283e080",
X"0c853d0d",
X"04fd3d0d",
X"75777053",
X"5454c73f",
X"83e08008",
X"732ea138",
X"83e08008",
X"733152ff",
X"125271ff",
X"2e8f3872",
X"70810554",
X"33747081",
X"055634eb",
X"39ff1454",
X"80743485",
X"3d0d0480",
X"3d0d7251",
X"ff903f82",
X"3d0d0471",
X"83e0800c",
X"04803d0d",
X"72518071",
X"34810bbc",
X"120c800b",
X"80c0120c",
X"823d0d04",
X"800b83e5",
X"bc08248a",
X"38a5f83f",
X"ff0b83e5",
X"bc0c800b",
X"83e0800c",
X"04ff3d0d",
X"735283e3",
X"9808722e",
X"8d38d93f",
X"71519785",
X"3f7183e3",
X"980c833d",
X"0d04f43d",
X"0d7e6062",
X"5c5a5581",
X"54bc1508",
X"81913874",
X"51cf3f79",
X"58807a25",
X"80f73883",
X"e5ec0870",
X"892a5783",
X"ff067884",
X"80723156",
X"56577378",
X"25833873",
X"557583e5",
X"bc082e84",
X"38ff893f",
X"83e5bc08",
X"8025a638",
X"75892b51",
X"99f13f83",
X"e5ec088f",
X"3dfc1155",
X"5c548152",
X"f81b5197",
X"d63f7614",
X"83e5ec0c",
X"7583e5bc",
X"0c745376",
X"527851a4",
X"a93f83e0",
X"800883e5",
X"ec081683",
X"e5ec0c78",
X"7631761b",
X"5b595677",
X"8024ff8b",
X"38617a71",
X"0c547554",
X"75802e83",
X"38815473",
X"83e0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"9b3f7651",
X"feaf3f86",
X"3dfc0553",
X"02a20522",
X"52775196",
X"f63f7986",
X"3d22710c",
X"5483e080",
X"085483e0",
X"8008802e",
X"83388154",
X"7383e080",
X"0c863d0d",
X"04fd3d0d",
X"7683e5bc",
X"08535380",
X"72248938",
X"71732e84",
X"38fdd13f",
X"7551fde5",
X"3f725198",
X"be3f7352",
X"73802e83",
X"38815271",
X"83e0800c",
X"853d0d04",
X"803d0d72",
X"80c01108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"72bc1108",
X"83e0800c",
X"51823d0d",
X"0480c40b",
X"83e0800c",
X"04fd3d0d",
X"75777154",
X"70535553",
X"a0e73f82",
X"c81308bc",
X"150c82c0",
X"130880c0",
X"150cfcec",
X"3f735194",
X"983f7383",
X"e3980c83",
X"e0800853",
X"83e08008",
X"802e8338",
X"81537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"5553fcc0",
X"3f72802e",
X"a538bc13",
X"08527351",
X"9ff13f83",
X"e080088f",
X"38775272",
X"51ff9a3f",
X"83e08008",
X"538a3982",
X"cc130853",
X"d8398153",
X"7283e080",
X"0c853d0d",
X"04fe3d0d",
X"ff0b83e5",
X"bc0c7483",
X"e39c0c75",
X"83e5b80c",
X"a0de3f83",
X"e0800881",
X"ff065281",
X"53719938",
X"83e5d451",
X"8f903f83",
X"e0800852",
X"83e08008",
X"802e8338",
X"72527153",
X"7283e080",
X"0c843d0d",
X"04fa3d0d",
X"787a82c4",
X"120882c4",
X"12087072",
X"24595656",
X"57577373",
X"2e098106",
X"913880c0",
X"165280c0",
X"17519de2",
X"3f83e080",
X"08557483",
X"e0800c88",
X"3d0d04f6",
X"3d0d7c5b",
X"807b715c",
X"54577a77",
X"2e8c3881",
X"1a82cc14",
X"08545a72",
X"f6388059",
X"80d9397a",
X"54815780",
X"707b7b31",
X"5a5755ff",
X"18537473",
X"2580c138",
X"82cc1408",
X"527351ff",
X"8c3f800b",
X"83e08008",
X"25a13882",
X"cc140882",
X"cc110882",
X"cc160c74",
X"82cc120c",
X"5375802e",
X"86387282",
X"cc170c72",
X"54805773",
X"82cc1508",
X"81175755",
X"56ffb839",
X"81195980",
X"0bff1b54",
X"54787325",
X"83388154",
X"76813270",
X"75065153",
X"72ff9038",
X"8c3d0d04",
X"f73d0d7b",
X"7d5a5a82",
X"d05283e5",
X"b80851a8",
X"9e3f83e0",
X"800857f9",
X"e33f7952",
X"83e5c051",
X"96c73f83",
X"e0800853",
X"805483e0",
X"8008742e",
X"09810682",
X"833883e3",
X"9c080b0b",
X"80faf853",
X"7052559d",
X"a03f0b0b",
X"80faf852",
X"80c01551",
X"9d933f74",
X"bc160c72",
X"82c0160c",
X"810b82c4",
X"160c810b",
X"82c8160c",
X"ff177357",
X"57819739",
X"83e3a833",
X"70822a70",
X"81065154",
X"54728186",
X"3873812a",
X"81065877",
X"80fc3876",
X"802e8190",
X"3882d015",
X"ff187584",
X"2a810682",
X"c4130c83",
X"e3a83381",
X"0682c813",
X"0c7b5471",
X"5358569c",
X"b43f7551",
X"9ccb3f83",
X"e0800816",
X"53af7370",
X"81055534",
X"72bc170c",
X"83e3a952",
X"72519c95",
X"3f83e3a0",
X"0882c017",
X"0c83e3b6",
X"52839015",
X"519c823f",
X"7782cc17",
X"0c78802e",
X"8d387551",
X"782d83e0",
X"8008802e",
X"8d387480",
X"2e863875",
X"82cc160c",
X"755583e3",
X"a05283e5",
X"c05195e7",
X"3f83e080",
X"088a3883",
X"e3a93353",
X"72fed138",
X"800b82cc",
X"170c7880",
X"2e893883",
X"e39c0851",
X"fcb93f83",
X"e39c0854",
X"7383e080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb63f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f692",
X"3f83e080",
X"08745387",
X"3d705355",
X"55f6b23f",
X"f7923f73",
X"51d33f63",
X"53745283",
X"e0800851",
X"fab93f92",
X"3d0d0471",
X"83e0800c",
X"0480c012",
X"83e0800c",
X"04803d0d",
X"7282c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"e0800c51",
X"823d0d04",
X"f63d0d7c",
X"83e09808",
X"59598179",
X"2782a938",
X"78881908",
X"2782a138",
X"77335675",
X"822e819b",
X"38758224",
X"89387581",
X"2e8d3882",
X"8b397583",
X"2e81b738",
X"82823978",
X"83ffff06",
X"70812a11",
X"7083ffff",
X"067083ff",
X"0671892a",
X"903d5f52",
X"5a515155",
X"7683ff2e",
X"8e388254",
X"76538c18",
X"08155279",
X"51a93975",
X"5476538c",
X"18081552",
X"79519ad8",
X"3f83e080",
X"0881bd38",
X"755483e0",
X"8008538c",
X"18081581",
X"05528c3d",
X"fd05519a",
X"bb3f83e0",
X"800881a0",
X"3802a905",
X"338c3d33",
X"71882b07",
X"7a810671",
X"842a5357",
X"58567486",
X"38769fff",
X"06567555",
X"81803975",
X"54781083",
X"fe065378",
X"882a8c19",
X"0805528c",
X"3dfc0551",
X"99fa3f83",
X"e0800880",
X"df3802a9",
X"05338c3d",
X"3371882b",
X"07565780",
X"d1398454",
X"78822b83",
X"fc065378",
X"872a8c19",
X"0805528c",
X"3dfc0551",
X"99ca3f83",
X"e08008b0",
X"3802ab05",
X"33028405",
X"aa053371",
X"982b7190",
X"2b07028c",
X"05a90533",
X"70882b72",
X"07903d33",
X"7180ffff",
X"fe800607",
X"51525357",
X"58568339",
X"81557483",
X"e0800c8c",
X"3d0d04fb",
X"3d0d83e0",
X"9808fe19",
X"881208fe",
X"05555654",
X"80567473",
X"278d3882",
X"14337571",
X"29941608",
X"05575375",
X"83e0800c",
X"873d0d04",
X"fc3d0d76",
X"83e09808",
X"55558075",
X"23881508",
X"5372812e",
X"88388814",
X"08732685",
X"388152b2",
X"39729038",
X"73335271",
X"832e0981",
X"06853890",
X"14085372",
X"8c160c72",
X"802e8d38",
X"7251ff93",
X"3f83e080",
X"08528539",
X"90140852",
X"7190160c",
X"80527183",
X"e0800c86",
X"3d0d04fa",
X"3d0d7883",
X"e0980871",
X"22810570",
X"83ffff06",
X"57545755",
X"73802e88",
X"38901508",
X"53728638",
X"835280e7",
X"39738f06",
X"527180da",
X"38811390",
X"160c8c15",
X"08537290",
X"38830b84",
X"17225752",
X"73762780",
X"c638bf39",
X"821633ff",
X"0574842a",
X"065271b2",
X"387251fb",
X"db3f8152",
X"7183e080",
X"0827a838",
X"835283e0",
X"80088817",
X"08279c38",
X"83e08008",
X"8c160c83",
X"e0800851",
X"fdf93f83",
X"e0800890",
X"160c7375",
X"23805271",
X"83e0800c",
X"883d0d04",
X"f23d0d60",
X"6264585d",
X"5b753355",
X"74a02e09",
X"81068838",
X"81167044",
X"56ef3962",
X"70335656",
X"74af2e09",
X"81068438",
X"81164380",
X"0b881c0c",
X"62703351",
X"5574a026",
X"91387a51",
X"fdd23f83",
X"e0800856",
X"807c3483",
X"a839933d",
X"841c0870",
X"585a5f8a",
X"55a07670",
X"81055834",
X"ff155574",
X"ff2e0981",
X"06ef3880",
X"70595d88",
X"7f085f5a",
X"7c811e70",
X"81ff0660",
X"13703370",
X"af327030",
X"a0732771",
X"80250751",
X"51525b53",
X"5f575574",
X"80d83876",
X"ae2e0981",
X"06833881",
X"55777a27",
X"75075574",
X"802e9f38",
X"79883270",
X"3078ae32",
X"70307073",
X"079f2a53",
X"51575156",
X"75ac3888",
X"588b5aff",
X"ab39ff9f",
X"17557499",
X"268938e0",
X"177081ff",
X"06585577",
X"81197081",
X"ff06721c",
X"535a5755",
X"767534ff",
X"87397c1e",
X"7f0c8055",
X"76a02683",
X"38815574",
X"8b1a347a",
X"51fc913f",
X"83e08008",
X"80f538a0",
X"547a2270",
X"852b83e0",
X"06545590",
X"1b08527b",
X"5194d13f",
X"83e08008",
X"5783e080",
X"08818238",
X"7b335574",
X"802e80f5",
X"388b1c33",
X"70832a70",
X"81065156",
X"5674b438",
X"8b7c841d",
X"0883e080",
X"08595b5b",
X"58ff1858",
X"77ff2e9a",
X"38797081",
X"055b3379",
X"7081055b",
X"33717131",
X"52565675",
X"802ee238",
X"86397580",
X"2ebc387a",
X"51fbf43f",
X"ff863983",
X"e0800856",
X"83e08008",
X"802ea938",
X"83e08008",
X"832e0981",
X"0680de38",
X"841b088b",
X"11335155",
X"7480d238",
X"845680cd",
X"398356ec",
X"39815680",
X"c4397656",
X"841b088b",
X"11335155",
X"74b7388b",
X"1c337084",
X"2a708106",
X"51565774",
X"802ed538",
X"951c3394",
X"1d337198",
X"2b71902b",
X"079b1f33",
X"7f9a0533",
X"71882b07",
X"72077f88",
X"050c5a58",
X"5658fcda",
X"397583e0",
X"800c903d",
X"0d04f83d",
X"0d7a7c59",
X"57825483",
X"fe537752",
X"765192e0",
X"3f835683",
X"e0800880",
X"ec388117",
X"33773371",
X"882b0756",
X"56825674",
X"82d4d52e",
X"09810680",
X"d4387554",
X"b6537752",
X"765192b4",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"ac388254",
X"80d25377",
X"52765192",
X"8b3f83e0",
X"80089838",
X"81173377",
X"3371882b",
X"0783e080",
X"08525656",
X"748182c6",
X"2e833881",
X"567583e0",
X"800c8a3d",
X"0d04ec3d",
X"0d665980",
X"0b83e098",
X"0c785678",
X"802e83e8",
X"3891a53f",
X"83e08008",
X"81065582",
X"567483d8",
X"38747553",
X"8e3d7053",
X"5858fec2",
X"3f83e080",
X"0881ff06",
X"5675812e",
X"09810680",
X"d4389054",
X"83be5374",
X"52765191",
X"973f83e0",
X"800880c9",
X"388e3d33",
X"5574802e",
X"80c93802",
X"bb053302",
X"8405ba05",
X"3371982b",
X"71902b07",
X"028c05b9",
X"05337088",
X"2b720794",
X"3d337107",
X"70587c57",
X"54525d57",
X"5956fde6",
X"3f83e080",
X"0881ff06",
X"5675832e",
X"09810686",
X"38815682",
X"db397580",
X"2e863887",
X"5682d139",
X"a4548d53",
X"77527651",
X"90ae3f81",
X"5683e080",
X"0882bd38",
X"02ba0533",
X"028405b9",
X"05337188",
X"2b07585c",
X"76ab3802",
X"80ca0533",
X"02840580",
X"c9053371",
X"982b7190",
X"2b07963d",
X"3370882b",
X"72070294",
X"0580c705",
X"33710754",
X"525d5758",
X"5602b305",
X"33777129",
X"028805b2",
X"0533028c",
X"05b10533",
X"71882b07",
X"701c708c",
X"1f0c5e59",
X"57585c8d",
X"3d33821a",
X"3402b505",
X"338f3d33",
X"71882b07",
X"595b7784",
X"1a2302b7",
X"05330284",
X"05b60533",
X"71882b07",
X"565b74ab",
X"380280c6",
X"05330284",
X"0580c505",
X"3371982b",
X"71902b07",
X"953d3370",
X"882b7207",
X"02940580",
X"c3053371",
X"07515253",
X"575d5b74",
X"76317731",
X"78842a8f",
X"3d335471",
X"71315356",
X"5698803f",
X"83e08008",
X"82057088",
X"1b0c709f",
X"f6268105",
X"575583ff",
X"f6752783",
X"38835675",
X"79347583",
X"2e098106",
X"af380280",
X"d2053302",
X"840580d1",
X"05337198",
X"2b71902b",
X"07983d33",
X"70882b72",
X"07029405",
X"80cf0533",
X"7107901f",
X"0c525d57",
X"59568639",
X"761a901a",
X"0c841922",
X"8c1a0818",
X"71842a05",
X"941b0c5c",
X"800b811a",
X"347883e0",
X"980c8056",
X"7583e080",
X"0c963d0d",
X"04e93d0d",
X"83e09808",
X"56865475",
X"802e81a6",
X"38800b81",
X"1734993d",
X"e011466a",
X"54c01153",
X"ec0551f6",
X"cf3f83e0",
X"80085483",
X"e0800881",
X"8538893d",
X"33547380",
X"2e933802",
X"ab053370",
X"842a7081",
X"06515555",
X"73802e86",
X"38835480",
X"e53902b5",
X"05338f3d",
X"3371982b",
X"71902b07",
X"028c05bb",
X"05330290",
X"05ba0533",
X"71882b07",
X"7207a01b",
X"0c029005",
X"bf053302",
X"9405be05",
X"3371982b",
X"71902b07",
X"029c05bd",
X"05337088",
X"2b720799",
X"3d337107",
X"7f9c050c",
X"5283e080",
X"08981f0c",
X"565a5252",
X"53575957",
X"810b8117",
X"3483e080",
X"08547383",
X"e0800c99",
X"3d0d04f5",
X"3d0d7d60",
X"028805ba",
X"05227283",
X"e098085b",
X"5d5a5c5c",
X"807b2386",
X"5676802e",
X"81e03881",
X"17338106",
X"55855674",
X"802e81d2",
X"389c1708",
X"98180831",
X"55747827",
X"87387483",
X"ffff0658",
X"77802e81",
X"ae389817",
X"087083ff",
X"06565674",
X"80ca3882",
X"1733ff05",
X"76892a06",
X"7081ff06",
X"5a5578a0",
X"38758738",
X"a0170855",
X"8d39a417",
X"0851efe0",
X"3f83e080",
X"08558175",
X"2780f838",
X"74a4180c",
X"a4170851",
X"f28d3f83",
X"e0800880",
X"2e80e438",
X"83e08008",
X"19a8180c",
X"98170883",
X"ff068480",
X"71317083",
X"ffff0658",
X"51557776",
X"27833877",
X"56755498",
X"170883ff",
X"0653a817",
X"08527955",
X"7b83387b",
X"5574518a",
X"d33f83e0",
X"8008a438",
X"98170816",
X"98180c75",
X"1a787731",
X"7083ffff",
X"067d2279",
X"05525a56",
X"5a747b23",
X"fece3980",
X"56883980",
X"0b811834",
X"81567583",
X"e0800c8d",
X"3d0d04fa",
X"3d0d7883",
X"e0980855",
X"56865573",
X"802e81dc",
X"38811433",
X"81065385",
X"5572802e",
X"81ce389c",
X"14085372",
X"76278338",
X"72569814",
X"0857800b",
X"98150c75",
X"802e81a9",
X"38821433",
X"70892b56",
X"5376802e",
X"b5387452",
X"ff165192",
X"ee3f83e0",
X"8008ff18",
X"76547053",
X"585392df",
X"3f83e080",
X"08732696",
X"38743070",
X"78067098",
X"170c7771",
X"31a41708",
X"52585153",
X"8939a014",
X"0870a416",
X"0c537476",
X"27b43872",
X"51edc13f",
X"83e08008",
X"53810b83",
X"e0800827",
X"80cb3883",
X"e0800888",
X"15082780",
X"c03883e0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c9399814",
X"08167098",
X"160c7352",
X"56efc83f",
X"83e08008",
X"802e9638",
X"821433ff",
X"0576892a",
X"0683e080",
X"0805a815",
X"0c805588",
X"39800b81",
X"15348155",
X"7483e080",
X"0c883d0d",
X"04ee3d0d",
X"64568655",
X"83e09808",
X"802e80f6",
X"38943df4",
X"1184180c",
X"6654d405",
X"527551f1",
X"973f83e0",
X"80085583",
X"e0800880",
X"cf38893d",
X"33547380",
X"2ebc3802",
X"ab053370",
X"842a7081",
X"06515555",
X"84557380",
X"2ebc3802",
X"b505338f",
X"3d337198",
X"2b71902b",
X"07028c05",
X"bb053302",
X"9005ba05",
X"3371882b",
X"07720788",
X"1b0c5357",
X"59577551",
X"eed23f83",
X"e0800855",
X"74832e09",
X"81068338",
X"84557483",
X"e0800c94",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405d",
X"865683e0",
X"9808802e",
X"849b389e",
X"3df40584",
X"1e0c7e98",
X"387c51ee",
X"973f83e0",
X"80085684",
X"84398141",
X"82803983",
X"4181fb39",
X"933d7f96",
X"05415980",
X"7f829505",
X"5f567560",
X"81ff0534",
X"8341901d",
X"08762e81",
X"dd38a054",
X"7c227085",
X"2b83e006",
X"5458901d",
X"08527851",
X"86ae3f83",
X"e0800841",
X"83e08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"e8387b81",
X"bf065574",
X"8f2480dd",
X"389a1933",
X"557480d5",
X"389c1933",
X"5574802e",
X"80cb38f3",
X"1e70585e",
X"8156758b",
X"2e098106",
X"85388e56",
X"8b39759a",
X"2e098106",
X"83389c56",
X"75197070",
X"81055233",
X"7133811a",
X"821a5f5b",
X"525b5574",
X"86387977",
X"34853980",
X"df773477",
X"7b57577a",
X"a02e0981",
X"06c03881",
X"567b81e5",
X"32703070",
X"9f2a5151",
X"557bae2e",
X"93387480",
X"2e8e3861",
X"832a7081",
X"06515574",
X"802e9738",
X"7c51ecf7",
X"3f83e080",
X"084183e0",
X"80088738",
X"901d08fe",
X"a5388060",
X"3475802e",
X"88387d52",
X"7f5183b1",
X"3f60802e",
X"8638800b",
X"901e0c60",
X"5660832e",
X"09810688",
X"38800b90",
X"1e0c8539",
X"6081d238",
X"891f5790",
X"1d08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347c51ea",
X"fe3f83e0",
X"80085683",
X"e0800883",
X"2e098106",
X"8838800b",
X"901e0c80",
X"56961f33",
X"55748a38",
X"891f5296",
X"1f5181b1",
X"3f7583e0",
X"800c9e3d",
X"0d04fd3d",
X"0d757753",
X"54733351",
X"70893871",
X"33517080",
X"2ea13873",
X"33723352",
X"53727127",
X"8538ff51",
X"94397073",
X"27853881",
X"518b3981",
X"14811353",
X"54d33980",
X"517083e0",
X"800c853d",
X"0d04fd3d",
X"0d757754",
X"54723370",
X"81ff0652",
X"5270802e",
X"a3387181",
X"ff068114",
X"ffbf1253",
X"54527099",
X"268938a0",
X"127081ff",
X"06535171",
X"74708105",
X"5634d239",
X"80743485",
X"3d0d04ff",
X"bd3d0d80",
X"c63d0852",
X"a53d7052",
X"54ffb33f",
X"80c73d08",
X"52853d70",
X"5253ffa6",
X"3f725273",
X"51fedf3f",
X"80c53d0d",
X"04fe3d0d",
X"74765353",
X"71708105",
X"53335170",
X"73708105",
X"553470f0",
X"38843d0d",
X"04fe3d0d",
X"74528072",
X"33525370",
X"732e8d38",
X"81128114",
X"71335354",
X"5270f538",
X"7283e080",
X"0c843d0d",
X"04fc3d0d",
X"76557483",
X"e680082e",
X"af388053",
X"745187cd",
X"3f83e080",
X"0881ff06",
X"ff147081",
X"ff067230",
X"709f2a51",
X"52555354",
X"72802e84",
X"3871dd38",
X"73fe3874",
X"83e6800c",
X"863d0d04",
X"ff3d0dff",
X"0b83e680",
X"0c84af3f",
X"81518791",
X"3f83e080",
X"0881ff06",
X"5271ee38",
X"81d63f71",
X"83e0800c",
X"833d0d04",
X"fc3d0d76",
X"028405a2",
X"05220288",
X"05a60522",
X"7a545555",
X"55ff823f",
X"72802ea0",
X"3883e694",
X"14337570",
X"81055734",
X"81147083",
X"ffff06ff",
X"157083ff",
X"ff065652",
X"5552dd39",
X"800b83e0",
X"800c863d",
X"0d04fc3d",
X"0d76787a",
X"11565355",
X"80537174",
X"2e933872",
X"15517033",
X"83e69413",
X"34811281",
X"145452ea",
X"39800b83",
X"e0800c86",
X"3d0d04fd",
X"3d0d9054",
X"83e68008",
X"5187803f",
X"83e08008",
X"81ff06ff",
X"15713071",
X"30707307",
X"9f2a729f",
X"2a065255",
X"52555372",
X"db38853d",
X"0d04ff3d",
X"0d83e68c",
X"081083e6",
X"84080780",
X"fce80852",
X"710c833d",
X"0d04800b",
X"83e68c0c",
X"e13f0481",
X"0b83e68c",
X"0cd83f04",
X"ed3f0471",
X"83e6880c",
X"04803d0d",
X"8051f43f",
X"810b83e6",
X"8c0c810b",
X"83e6840c",
X"ffb83f82",
X"3d0d0480",
X"3d0d7230",
X"70740780",
X"2583e684",
X"0c51ffa2",
X"3f823d0d",
X"04fe3d0d",
X"02930533",
X"80fcec08",
X"54730c80",
X"fce80852",
X"71087081",
X"06515170",
X"f7387208",
X"7081ff06",
X"83e0800c",
X"51843d0d",
X"04803d0d",
X"81ff51cd",
X"3f83e080",
X"0881ff06",
X"83e0800c",
X"823d0d04",
X"ff3d0d74",
X"902b7407",
X"80fcdc08",
X"52710c83",
X"3d0d0404",
X"fb3d0d78",
X"0284059f",
X"05337098",
X"2b555755",
X"7280259b",
X"387580ff",
X"06568052",
X"80f751e0",
X"3f83e080",
X"0881ff06",
X"54738126",
X"80ff3880",
X"51fee03f",
X"ff9f3f81",
X"51fed83f",
X"ff973f75",
X"51fee63f",
X"74982a51",
X"fedf3f74",
X"902a7081",
X"ff065253",
X"fed33f74",
X"882a7081",
X"ff065253",
X"fec73f74",
X"81ff0651",
X"febf3f81",
X"557580c0",
X"2e098106",
X"86388195",
X"558d3975",
X"80c82e09",
X"81068438",
X"81875574",
X"51fe9e3f",
X"8a55fec5",
X"3f83e080",
X"0881ff06",
X"70982b54",
X"54728025",
X"8c38ff15",
X"7081ff06",
X"565374e2",
X"387383e0",
X"800c873d",
X"0d04fa3d",
X"0dfdbe3f",
X"8051fdd3",
X"3f8a54fe",
X"903fff14",
X"7081ff06",
X"555373f3",
X"38737453",
X"5580c051",
X"fea63f83",
X"e0800881",
X"ff065473",
X"812e0981",
X"0682a138",
X"83aa5280",
X"c851fe8c",
X"3f83e080",
X"0881ff06",
X"5372812e",
X"09810681",
X"a9387454",
X"873d7411",
X"5456fdc5",
X"3f83e080",
X"08733481",
X"147081ff",
X"06555383",
X"7427e538",
X"029a0533",
X"5372812e",
X"09810681",
X"db38029b",
X"05335380",
X"ce905472",
X"81aa2e8e",
X"3881c939",
X"80e451ff",
X"9fbe3fff",
X"14547380",
X"2e81b938",
X"820a5281",
X"e951fda4",
X"3f83e080",
X"0881ff06",
X"5372dd38",
X"725280fa",
X"51fd913f",
X"83e08008",
X"81ff0653",
X"72819138",
X"72547316",
X"53fcd23f",
X"83e08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e83887",
X"3d337086",
X"2a708106",
X"5154548c",
X"557280e4",
X"38845580",
X"df397452",
X"81e951fc",
X"cb3f83e0",
X"800881ff",
X"06538255",
X"81e95681",
X"73278638",
X"735580c1",
X"5680ce90",
X"548b3980",
X"e451ff9e",
X"af3fff14",
X"5473802e",
X"a9388052",
X"7551fc98",
X"3f83e080",
X"0881ff06",
X"5372e038",
X"84805280",
X"d051fc84",
X"3f83e080",
X"0881ff06",
X"5372802e",
X"83388055",
X"7483e690",
X"348051fa",
X"fe3ffbbd",
X"3f883d0d",
X"04fb3d0d",
X"7754800b",
X"83e69033",
X"70832a70",
X"81065155",
X"57557275",
X"2e098106",
X"85387389",
X"2b547352",
X"80d151fb",
X"bb3f83e0",
X"800881ff",
X"065372bd",
X"3882b8c0",
X"54fafe3f",
X"83e08008",
X"81ff0653",
X"7281ff2e",
X"09810689",
X"38ff1454",
X"73e7389f",
X"397281fe",
X"2e098106",
X"963883ea",
X"945283e6",
X"9451fae8",
X"3fface3f",
X"facb3f83",
X"39815580",
X"51fa803f",
X"fabf3f74",
X"81ff0683",
X"e0800c87",
X"3d0d04fb",
X"3d0d7783",
X"e6945654",
X"8151f9e3",
X"3f83e690",
X"3370832a",
X"70810651",
X"54567285",
X"3873892b",
X"54735280",
X"d851fab4",
X"3f83e080",
X"0881ff06",
X"537280e5",
X"3881ff51",
X"f9cb3f81",
X"fe51f9c5",
X"3f848053",
X"74708105",
X"563351f9",
X"b83fff13",
X"7083ffff",
X"06515372",
X"eb387251",
X"f9a73f72",
X"51f9a23f",
X"f9cb3f83",
X"e080089f",
X"0653a788",
X"5472852e",
X"8d389a39",
X"80e451ff",
X"9be63fff",
X"1454f9ad",
X"3f83e080",
X"0881ff2e",
X"843873e8",
X"388051f8",
X"da3ff999",
X"3f800b83",
X"e0800c87",
X"3d0d0483",
X"e08c0802",
X"83e08c0c",
X"fd3d0d80",
X"5383e08c",
X"088c0508",
X"5283e08c",
X"08880508",
X"5183d43f",
X"83e08008",
X"7083e080",
X"0c54853d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cfd",
X"3d0d8153",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"83a13f83",
X"e0800870",
X"83e0800c",
X"54853d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cf93d",
X"0d800b83",
X"e08c08fc",
X"050c83e0",
X"8c088805",
X"088025b9",
X"3883e08c",
X"08880508",
X"3083e08c",
X"0888050c",
X"800b83e0",
X"8c08f405",
X"0c83e08c",
X"08fc0508",
X"8a38810b",
X"83e08c08",
X"f4050c83",
X"e08c08f4",
X"050883e0",
X"8c08fc05",
X"0c83e08c",
X"088c0508",
X"8025b938",
X"83e08c08",
X"8c050830",
X"83e08c08",
X"8c050c80",
X"0b83e08c",
X"08f0050c",
X"83e08c08",
X"fc05088a",
X"38810b83",
X"e08c08f0",
X"050c83e0",
X"8c08f005",
X"0883e08c",
X"08fc050c",
X"805383e0",
X"8c088c05",
X"085283e0",
X"8c088805",
X"085181df",
X"3f83e080",
X"087083e0",
X"8c08f805",
X"0c5483e0",
X"8c08fc05",
X"08802e90",
X"3883e08c",
X"08f80508",
X"3083e08c",
X"08f8050c",
X"83e08c08",
X"f8050870",
X"83e0800c",
X"54893d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cfb3d",
X"0d800b83",
X"e08c08fc",
X"050c83e0",
X"8c088805",
X"08802599",
X"3883e08c",
X"08880508",
X"3083e08c",
X"0888050c",
X"810b83e0",
X"8c08fc05",
X"0c83e08c",
X"088c0508",
X"80259038",
X"83e08c08",
X"8c050830",
X"83e08c08",
X"8c050c81",
X"5383e08c",
X"088c0508",
X"5283e08c",
X"08880508",
X"51bd3f83",
X"e0800870",
X"83e08c08",
X"f8050c54",
X"83e08c08",
X"fc050880",
X"2e903883",
X"e08c08f8",
X"05083083",
X"e08c08f8",
X"050c83e0",
X"8c08f805",
X"087083e0",
X"800c5487",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"fd3d0d81",
X"0b83e08c",
X"08fc050c",
X"800b83e0",
X"8c08f805",
X"0c83e08c",
X"088c0508",
X"83e08c08",
X"88050827",
X"b93883e0",
X"8c08fc05",
X"08802eae",
X"38800b83",
X"e08c088c",
X"050824a2",
X"3883e08c",
X"088c0508",
X"1083e08c",
X"088c050c",
X"83e08c08",
X"fc050810",
X"83e08c08",
X"fc050cff",
X"b83983e0",
X"8c08fc05",
X"08802e80",
X"e13883e0",
X"8c088c05",
X"0883e08c",
X"08880508",
X"26ad3883",
X"e08c0888",
X"050883e0",
X"8c088c05",
X"083183e0",
X"8c088805",
X"0c83e08c",
X"08f80508",
X"83e08c08",
X"fc050807",
X"83e08c08",
X"f8050c83",
X"e08c08fc",
X"0508812a",
X"83e08c08",
X"fc050c83",
X"e08c088c",
X"0508812a",
X"83e08c08",
X"8c050cff",
X"953983e0",
X"8c089005",
X"08802e93",
X"3883e08c",
X"08880508",
X"7083e08c",
X"08f4050c",
X"51913983",
X"e08c08f8",
X"05087083",
X"e08c08f4",
X"050c5183",
X"e08c08f4",
X"050883e0",
X"800c853d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cff",
X"3d0d800b",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"05088106",
X"ff117009",
X"7083e08c",
X"088c0508",
X"0683e08c",
X"08fc0508",
X"1183e08c",
X"08fc050c",
X"83e08c08",
X"88050881",
X"2a83e08c",
X"0888050c",
X"83e08c08",
X"8c050810",
X"83e08c08",
X"8c050c51",
X"51515183",
X"e08c0888",
X"0508802e",
X"8438ffab",
X"3983e08c",
X"08fc0508",
X"7083e080",
X"0c51833d",
X"0d83e08c",
X"0c04fc3d",
X"0d767079",
X"7b555555",
X"558f7227",
X"8c387275",
X"07830651",
X"70802ea9",
X"38ff1252",
X"71ff2e98",
X"38727081",
X"05543374",
X"70810556",
X"34ff1252",
X"71ff2e09",
X"8106ea38",
X"7483e080",
X"0c863d0d",
X"04745172",
X"70840554",
X"08717084",
X"05530c72",
X"70840554",
X"08717084",
X"05530c72",
X"70840554",
X"08717084",
X"05530c72",
X"70840554",
X"08717084",
X"05530cf0",
X"1252718f",
X"26c93883",
X"72279538",
X"72708405",
X"54087170",
X"8405530c",
X"fc125271",
X"8326ed38",
X"7054ff81",
X"39000000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"000009a7",
X"000009e8",
X"00000a0a",
X"00000a28",
X"00000a28",
X"00000a28",
X"00000a28",
X"00000a97",
X"00000ac7",
X"70704740",
X"9c704268",
X"9c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"43617274",
X"72696467",
X"6520386b",
X"2073696d",
X"706c6500",
X"45786974",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"25732025",
X"73000000",
X"2e2e0000",
X"2f000000",
X"41545200",
X"58464400",
X"58455800",
X"524f4d00",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"6e616d65",
X"20000000",
X"25303278",
X"00000000",
X"00000000",
X"00000000",
X"00003cbc",
X"00003cc0",
X"00003cc8",
X"00003cd4",
X"00003ce0",
X"00003cec",
X"00003cf8",
X"00003cfc",
X"0001d20f",
X"0001d400",
X"0001d401",
X"0001d409",
X"0001d010",
X"0001d301",
X"0001d300",
X"0001d20a",
X"0001d01b",
X"0001d016",
X"0001d019",
X"0001d018",
X"0001d017",
X"0001d01a",
X"0001d403",
X"0001d402",
X"0001d40e",
X"0004007c",
X"00040078",
X"00040074",
X"00040068",
X"00040060",
X"0004005c",
X"00040058",
X"00040054",
X"00040050",
X"0004004c",
X"00040048",
X"00040044",
X"00040040",
X"00040034",
X"00040030",
X"0004002c",
X"00040028",
X"00040024",
X"00040020",
X"0004001c",
X"00040018",
X"00040014",
X"00040010",
X"0004000c",
X"00040008",
X"00040004",
X"00040000",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"69383030",
X"00000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
