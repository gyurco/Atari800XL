
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81d3",
X"e4738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81da",
X"fc0c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757580f3",
X"d52d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7580f394",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80dc8304",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"775193c4",
X"3f83c080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3381db84",
X"0b81db84",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"52775192",
X"f33f83c0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583c0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"55b3a83f",
X"83c08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"811451b2",
X"c03f83c0",
X"80083070",
X"83c08008",
X"07802583",
X"c0800c53",
X"863d0d04",
X"fc3d0d76",
X"70525599",
X"e03f83c0",
X"80085481",
X"5383c080",
X"0880c738",
X"745199a3",
X"3f83c080",
X"080b0b81",
X"d8f85383",
X"c0800852",
X"53ff8f3f",
X"83c08008",
X"a5380b0b",
X"81d8fc52",
X"7251fefe",
X"3f83c080",
X"0894380b",
X"0b81d980",
X"527251fe",
X"ed3f83c0",
X"8008802e",
X"83388154",
X"73537283",
X"c0800c86",
X"3d0d04fd",
X"3d0d7570",
X"525498f9",
X"3f815383",
X"c0800898",
X"38735198",
X"c23f83c0",
X"b0085283",
X"c0800851",
X"feb43f83",
X"c0800853",
X"7283c080",
X"0c853d0d",
X"04df3d0d",
X"a43d0870",
X"525e8ee7",
X"3f83c080",
X"0833953d",
X"56547396",
X"3881de94",
X"527451b1",
X"9a3f9a39",
X"7d527851",
X"91e83f84",
X"e3397d51",
X"8ecd3f83",
X"c0800852",
X"74518dfd",
X"3f804380",
X"42804180",
X"4083c0b8",
X"0852943d",
X"70525d94",
X"d03f83c0",
X"80085980",
X"0b83c080",
X"08555b83",
X"c080087b",
X"2e943881",
X"1b74525b",
X"97d23f83",
X"c0800854",
X"83c08008",
X"ee38805a",
X"ff5f7909",
X"709f2c7b",
X"065b547a",
X"7a248438",
X"ff1b5af6",
X"1a700970",
X"9f2c7206",
X"7bff125a",
X"5a525555",
X"80752595",
X"38765197",
X"973f83c0",
X"800876ff",
X"18585557",
X"738024ed",
X"38747f2e",
X"873880c2",
X"fa3f745f",
X"78ff1b70",
X"585d5880",
X"7a259538",
X"775196ec",
X"3f83c080",
X"0876ff18",
X"58555873",
X"8024ed38",
X"800b83c7",
X"d00c800b",
X"83c8940c",
X"0b0b81d9",
X"84518bbe",
X"3f81800b",
X"83c8940c",
X"0b0b81d9",
X"8c518bae",
X"3fa80b83",
X"c7d00c76",
X"802e80e8",
X"3883c7d0",
X"08777932",
X"70307072",
X"07802570",
X"872b83c8",
X"940c5156",
X"78535656",
X"969f3f83",
X"c0800880",
X"2e8a380b",
X"0b81d994",
X"518af33f",
X"765195df",
X"3f83c080",
X"08520b0b",
X"81daa051",
X"8ae03f76",
X"5195e53f",
X"83c08008",
X"83c7d008",
X"55577574",
X"258638a8",
X"1656f739",
X"7583c7d0",
X"0c86f076",
X"24ff9438",
X"87980b83",
X"c7d00c77",
X"802eb738",
X"7751959b",
X"3f83c080",
X"08785255",
X"95bb3f0b",
X"0b81d99c",
X"5483c080",
X"088f3887",
X"39807634",
X"81d8390b",
X"0b81d998",
X"54745373",
X"520b0b81",
X"d8ec5189",
X"f93f8054",
X"0b0b81da",
X"f85189ee",
X"3f811454",
X"73a82e09",
X"8106ed38",
X"868da051",
X"beef3f80",
X"52903d70",
X"525780e1",
X"d33f8352",
X"765180e1",
X"cb3f6281",
X"91386180",
X"2e80fd38",
X"7b5473ff",
X"2e963878",
X"802e818c",
X"38785194",
X"b73f83c0",
X"8008ff15",
X"5559e739",
X"78802e80",
X"f7387851",
X"94b33f83",
X"c0800880",
X"2efbfd38",
X"785193fb",
X"3f83c080",
X"08520b0b",
X"81d8f451",
X"abda3f83",
X"c08008a3",
X"387c51ad",
X"923f83c0",
X"80085574",
X"ff165654",
X"807425ae",
X"38741d70",
X"33555673",
X"af2efec5",
X"38e93978",
X"5193ba3f",
X"83c08008",
X"527c51ac",
X"ca3f8f39",
X"7f882960",
X"10057a05",
X"61055afb",
X"fd396280",
X"2efbbe38",
X"80527651",
X"80e0a93f",
X"a33d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"842a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"a80b9088",
X"b834b80b",
X"9088b834",
X"7083c080",
X"0c823d0d",
X"04803d0d",
X"9088b833",
X"7081ff06",
X"70852a81",
X"32708106",
X"51515151",
X"70802e8d",
X"38980b90",
X"88b834b8",
X"0b9088b8",
X"347083c0",
X"800c823d",
X"0d04930b",
X"9088bc34",
X"ff0b9088",
X"a83404ff",
X"3d0d028f",
X"05335280",
X"0b9088bc",
X"348a51bc",
X"b43fdf3f",
X"80f80b90",
X"88a03480",
X"0b908888",
X"34fa1252",
X"71908880",
X"34800b90",
X"88983471",
X"90889034",
X"9088b852",
X"807234b8",
X"7234833d",
X"0d04803d",
X"0d028b05",
X"33517090",
X"88b434fe",
X"bf3f83c0",
X"8008802e",
X"f638823d",
X"0d04803d",
X"0d853980",
X"c6873ffe",
X"d83f83c0",
X"8008802e",
X"f2389088",
X"b4337081",
X"ff0683c0",
X"800c5182",
X"3d0d0480",
X"3d0da30b",
X"9088bc34",
X"ff0b9088",
X"a8349088",
X"b851a871",
X"34b87134",
X"823d0d04",
X"803d0d90",
X"88bc3370",
X"81c00670",
X"30708025",
X"83c0800c",
X"51515182",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067083",
X"2a813270",
X"81065151",
X"51517080",
X"2ee838b0",
X"0b9088b8",
X"34b80b90",
X"88b83482",
X"3d0d0480",
X"3d0d9080",
X"ac088106",
X"83c0800c",
X"823d0d04",
X"fd3d0d75",
X"77545480",
X"73259438",
X"73708105",
X"55335281",
X"d9a05185",
X"a13fff13",
X"53e93985",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"80dea93f",
X"83c08008",
X"7a27ed38",
X"74802e80",
X"e0387452",
X"755180de",
X"933f83c0",
X"80087553",
X"76525480",
X"de963f83",
X"c080087a",
X"53755256",
X"80ddf93f",
X"83c08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"c08008c2",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9c",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fbfd3f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd13f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbad3f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83c0900c",
X"7183c094",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383c090",
X"085283c0",
X"940851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"99e65351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fd3d",
X"0d757052",
X"54a3c43f",
X"83c08008",
X"14537274",
X"2e9238ff",
X"13703353",
X"5371af2e",
X"098106ee",
X"38811353",
X"7283c080",
X"0c853d0d",
X"04fd3d0d",
X"75777053",
X"5454c73f",
X"83c08008",
X"732ea138",
X"83c08008",
X"733152ff",
X"125271ff",
X"2e8f3872",
X"70810554",
X"33747081",
X"055634eb",
X"39ff1454",
X"80743485",
X"3d0d0480",
X"3d0d7251",
X"ff903f82",
X"3d0d0471",
X"83c0800c",
X"04803d0d",
X"72518071",
X"34810bbc",
X"120c800b",
X"80c0120c",
X"823d0d04",
X"800b83c2",
X"e408248a",
X"38a4ae3f",
X"ff0b83c2",
X"e40c800b",
X"83c0800c",
X"04ff3d0d",
X"735283c0",
X"c008722e",
X"8d38d93f",
X"71519699",
X"3f7183c0",
X"c00c833d",
X"0d04f43d",
X"0d7e6062",
X"5c5a5581",
X"54bc1508",
X"81913874",
X"51cf3f79",
X"58807a25",
X"80f73883",
X"c3940870",
X"892a5783",
X"ff067884",
X"80723156",
X"56577378",
X"25833873",
X"557583c2",
X"e4082e84",
X"38ff893f",
X"83c2e408",
X"8025a638",
X"75892b51",
X"98dc3f83",
X"c394088f",
X"3dfc1155",
X"5c548152",
X"f81b5196",
X"c63f7614",
X"83c3940c",
X"7583c2e4",
X"0c745376",
X"527851a2",
X"df3f83c0",
X"800883c3",
X"94081683",
X"c3940c78",
X"7631761b",
X"5b595677",
X"8024ff8b",
X"38617a71",
X"0c547554",
X"75802e83",
X"38815473",
X"83c0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"9b3f7651",
X"feaf3f86",
X"3dfc0553",
X"78527751",
X"95e93f79",
X"75710c54",
X"83c08008",
X"5483c080",
X"08802e83",
X"38815473",
X"83c0800c",
X"863d0d04",
X"fe3d0d75",
X"83c2e408",
X"53538072",
X"24893871",
X"732e8438",
X"fdd63f74",
X"51fdea3f",
X"725197ae",
X"3f83c080",
X"085283c0",
X"8008802e",
X"83388152",
X"7183c080",
X"0c843d0d",
X"04803d0d",
X"7280c011",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d72bc11",
X"0883c080",
X"0c51823d",
X"0d0480c4",
X"0b83c080",
X"0c04fd3d",
X"0d757771",
X"54705355",
X"539f9c3f",
X"82c81308",
X"bc150c82",
X"c0130880",
X"c0150cfc",
X"eb3f7351",
X"93ab3f73",
X"83c0c00c",
X"83c08008",
X"5383c080",
X"08802e83",
X"38815372",
X"83c0800c",
X"853d0d04",
X"fd3d0d75",
X"775553fc",
X"bf3f7280",
X"2ea538bc",
X"13085273",
X"519ea63f",
X"83c08008",
X"8f387752",
X"7251ff9a",
X"3f83c080",
X"08538a39",
X"82cc1308",
X"53d83981",
X"537283c0",
X"800c853d",
X"0d04fe3d",
X"0dff0b83",
X"c2e40c74",
X"83c0c40c",
X"7583c2e0",
X"0c9f933f",
X"83c08008",
X"81ff0652",
X"81537199",
X"3883c2fc",
X"518e943f",
X"83c08008",
X"5283c080",
X"08802e83",
X"38725271",
X"537283c0",
X"800c843d",
X"0d04fa3d",
X"0d787a82",
X"c4120882",
X"c4120870",
X"72245956",
X"56575773",
X"732e0981",
X"06913880",
X"c0165280",
X"c017519c",
X"973f83c0",
X"80085574",
X"83c0800c",
X"883d0d04",
X"f63d0d7c",
X"5b807b71",
X"5c54577a",
X"772e8c38",
X"811a82cc",
X"1408545a",
X"72f63880",
X"5980d939",
X"7a548157",
X"80707b7b",
X"315a5755",
X"ff185374",
X"732580c1",
X"3882cc14",
X"08527351",
X"ff8c3f80",
X"0b83c080",
X"0825a138",
X"82cc1408",
X"82cc1108",
X"82cc160c",
X"7482cc12",
X"0c537580",
X"2e863872",
X"82cc170c",
X"72548057",
X"7382cc15",
X"08811757",
X"5556ffb8",
X"39811959",
X"800bff1b",
X"54547873",
X"25833881",
X"54768132",
X"70750651",
X"5372ff90",
X"388c3d0d",
X"04f73d0d",
X"7b7d5a5a",
X"82d05283",
X"c2e00851",
X"80d1b13f",
X"83c08008",
X"57f9e13f",
X"795283c2",
X"e85195b5",
X"3f83c080",
X"08548053",
X"83c08008",
X"732e0981",
X"06828338",
X"83c0c408",
X"0b0b81d8",
X"f4537052",
X"569bd43f",
X"0b0b81d8",
X"f45280c0",
X"16519bc7",
X"3f75bc17",
X"0c7382c0",
X"170c810b",
X"82c4170c",
X"810b82c8",
X"170c7382",
X"cc170cff",
X"1782d017",
X"55578191",
X"3983c0d0",
X"3370822a",
X"70810651",
X"54557281",
X"80387481",
X"2a810658",
X"7780f638",
X"74842a81",
X"0682c415",
X"0c83c0d0",
X"33810682",
X"c8150c79",
X"5273519a",
X"ee3f7351",
X"9b853f83",
X"c0800814",
X"53af7370",
X"81055534",
X"72bc150c",
X"83c0d152",
X"72519acf",
X"3f83c0c8",
X"0882c015",
X"0c83c0de",
X"5280c014",
X"519abc3f",
X"78802e8d",
X"38735178",
X"2d83c080",
X"08802e99",
X"387782cc",
X"150c7580",
X"2e863873",
X"82cc170c",
X"7382d015",
X"ff195955",
X"5676802e",
X"9b3883c0",
X"c85283c2",
X"e85194ab",
X"3f83c080",
X"088a3883",
X"c0d13353",
X"72fed238",
X"78802e89",
X"3883c0c4",
X"0851fcb8",
X"3f83c0c4",
X"08537283",
X"c0800c8b",
X"3d0d04ff",
X"3d0d8052",
X"7351fdb5",
X"3f833d0d",
X"04f03d0d",
X"62705254",
X"f6903f83",
X"c0800874",
X"53873d70",
X"535555f6",
X"b03ff790",
X"3f7351d3",
X"3f635374",
X"5283c080",
X"0851fab8",
X"3f923d0d",
X"047183c0",
X"800c0480",
X"c01283c0",
X"800c0480",
X"3d0d7282",
X"c0110883",
X"c0800c51",
X"823d0d04",
X"803d0d72",
X"82cc1108",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"7282c411",
X"0883c080",
X"0c51823d",
X"0d04f93d",
X"0d7983c0",
X"98085757",
X"81772781",
X"96387688",
X"17082781",
X"8e387533",
X"5574822e",
X"89387483",
X"2eb33880",
X"fe397454",
X"761083fe",
X"06537688",
X"2a8c1708",
X"0552893d",
X"fc055199",
X"c13f83c0",
X"800880df",
X"38029d05",
X"33893d33",
X"71882b07",
X"565680d1",
X"39845476",
X"822b83fc",
X"06537687",
X"2a8c1708",
X"0552893d",
X"fc055199",
X"913f83c0",
X"8008b038",
X"029f0533",
X"0284059e",
X"05337198",
X"2b71902b",
X"07028c05",
X"9d053370",
X"882b7207",
X"8d3d3371",
X"80fffffe",
X"80060751",
X"52535758",
X"56833981",
X"557483c0",
X"800c893d",
X"0d04fb3d",
X"0d83c098",
X"08fe1988",
X"1208fe05",
X"55565480",
X"56747327",
X"8d388214",
X"33757129",
X"94160805",
X"57537583",
X"c0800c87",
X"3d0d04fc",
X"3d0d7652",
X"800b83c0",
X"98087033",
X"51525370",
X"832e0981",
X"06913895",
X"12339413",
X"3371982b",
X"71902b07",
X"5555519b",
X"12339a13",
X"3371882b",
X"07740783",
X"c0800c55",
X"863d0d04",
X"fc3d0d76",
X"83c09808",
X"55558075",
X"23881508",
X"5372812e",
X"88388814",
X"08732685",
X"388152b2",
X"39729038",
X"73335271",
X"832e0981",
X"06853890",
X"14085372",
X"8c160c72",
X"802e8d38",
X"7251fed6",
X"3f83c080",
X"08528539",
X"90140852",
X"7190160c",
X"80527183",
X"c0800c86",
X"3d0d04fa",
X"3d0d7883",
X"c0980871",
X"22810570",
X"83ffff06",
X"57545755",
X"73802e88",
X"38901508",
X"53728638",
X"835280e7",
X"39738f06",
X"527180da",
X"38811390",
X"160c8c15",
X"08537290",
X"38830b84",
X"17225752",
X"73762780",
X"c638bf39",
X"821633ff",
X"0574842a",
X"065271b2",
X"387251fc",
X"b13f8152",
X"7183c080",
X"0827a838",
X"835283c0",
X"80088817",
X"08279c38",
X"83c08008",
X"8c160c83",
X"c0800851",
X"fdbc3f83",
X"c0800890",
X"160c7375",
X"23805271",
X"83c0800c",
X"883d0d04",
X"f23d0d60",
X"6264585e",
X"5b753355",
X"74a02e09",
X"81068838",
X"81167044",
X"56ef3962",
X"70335656",
X"74af2e09",
X"81068438",
X"81164380",
X"0b881c0c",
X"62703351",
X"55749f26",
X"91387a51",
X"fdd23f83",
X"c0800856",
X"807d3483",
X"8139933d",
X"841c0870",
X"58595f8a",
X"55a07670",
X"81055834",
X"ff155574",
X"ff2e0981",
X"06ef3880",
X"705a5c88",
X"7f085f5a",
X"7b811d70",
X"81ff0660",
X"13703370",
X"af327030",
X"a0732771",
X"80250751",
X"51525b53",
X"5e575574",
X"80e73876",
X"ae2e0981",
X"06833881",
X"55787a27",
X"75075574",
X"802e9f38",
X"79883270",
X"3078ae32",
X"70307073",
X"079f2a53",
X"51575156",
X"75bb3888",
X"598b5aff",
X"ab397698",
X"2b557480",
X"25873881",
X"d2f41733",
X"57ff9f17",
X"55749926",
X"8938e017",
X"7081ff06",
X"58557881",
X"1a7081ff",
X"06721b53",
X"5b575576",
X"7534fef8",
X"397b1e7f",
X"0c805576",
X"a0268338",
X"8155748b",
X"19347a51",
X"fc823f83",
X"c0800880",
X"f538a054",
X"7a227085",
X"2b83e006",
X"5455901b",
X"08527c51",
X"93cc3f83",
X"c0800857",
X"83c08008",
X"8181387c",
X"33557480",
X"2e80f438",
X"8b1d3370",
X"832a7081",
X"06515656",
X"74b4388b",
X"7d841d08",
X"83c08008",
X"595b5b58",
X"ff185877",
X"ff2e9a38",
X"79708105",
X"5b337970",
X"81055b33",
X"71713152",
X"56567580",
X"2ee23886",
X"3975802e",
X"96387a51",
X"fbe53fff",
X"863983c0",
X"80085683",
X"c08008b6",
X"38833976",
X"56841b08",
X"8b113351",
X"5574a738",
X"8b1d3370",
X"842a7081",
X"06515656",
X"74893883",
X"56943981",
X"5690397c",
X"51fa943f",
X"83c08008",
X"881c0cfd",
X"81397583",
X"c0800c90",
X"3d0d04f8",
X"3d0d7a7c",
X"59578254",
X"83fe5377",
X"52765192",
X"913f8356",
X"83c08008",
X"80ec3881",
X"17337733",
X"71882b07",
X"56568256",
X"7482d4d5",
X"2e098106",
X"80d43875",
X"54b65377",
X"52765191",
X"e53f83c0",
X"80089838",
X"81173377",
X"3371882b",
X"0783c080",
X"08525656",
X"748182c6",
X"2eac3882",
X"5480d253",
X"77527651",
X"91bc3f83",
X"c0800898",
X"38811733",
X"77337188",
X"2b0783c0",
X"80085256",
X"56748182",
X"c62e8338",
X"81567583",
X"c0800c8a",
X"3d0d04eb",
X"3d0d675a",
X"800b83c0",
X"980c90de",
X"3f83c080",
X"08810655",
X"82567483",
X"ef387475",
X"538f3d70",
X"535759fe",
X"ca3f83c0",
X"800881ff",
X"06577681",
X"2e098106",
X"80d43890",
X"5483be53",
X"74527551",
X"90d03f83",
X"c0800880",
X"c9388f3d",
X"33557480",
X"2e80c938",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"0770587b",
X"575e525e",
X"575957fd",
X"ee3f83c0",
X"800881ff",
X"06577683",
X"2e098106",
X"86388156",
X"82f23976",
X"802e8638",
X"865682e8",
X"39a4548d",
X"53785275",
X"518fe73f",
X"815683c0",
X"800882d4",
X"3802be05",
X"33028405",
X"bd053371",
X"882b0759",
X"5d77ab38",
X"0280ce05",
X"33028405",
X"80cd0533",
X"71982b71",
X"902b0797",
X"3d337088",
X"2b720702",
X"940580cb",
X"05337107",
X"54525e57",
X"595602b7",
X"05337871",
X"29028805",
X"b6053302",
X"8c05b505",
X"3371882b",
X"07701d70",
X"7f8c050c",
X"5f595759",
X"5d8e3d33",
X"821b3402",
X"b9053390",
X"3d337188",
X"2b075a5c",
X"78841b23",
X"02bb0533",
X"028405ba",
X"05337188",
X"2b07565c",
X"74ab3802",
X"80ca0533",
X"02840580",
X"c9053371",
X"982b7190",
X"2b07963d",
X"3370882b",
X"72070294",
X"0580c705",
X"33710751",
X"5253575e",
X"5c747631",
X"78317984",
X"2a903d33",
X"54717131",
X"53565680",
X"c2963f83",
X"c0800882",
X"0570881c",
X"0c83c080",
X"08e08a05",
X"56567483",
X"dffe2683",
X"38825783",
X"fff67627",
X"85388357",
X"89398656",
X"76802e80",
X"db38767a",
X"3476832e",
X"098106b0",
X"380280d6",
X"05330284",
X"0580d505",
X"3371982b",
X"71902b07",
X"993d3370",
X"882b7207",
X"02940580",
X"d3053371",
X"077f9005",
X"0c525e57",
X"58568639",
X"771b901b",
X"0c841a22",
X"8c1b0819",
X"71842a05",
X"941c0c5d",
X"800b811b",
X"347983c0",
X"980c8056",
X"7583c080",
X"0c973d0d",
X"04e93d0d",
X"83c09808",
X"56855475",
X"802e8182",
X"38800b81",
X"1734993d",
X"e011466a",
X"548a3d70",
X"5458ec05",
X"51f6e53f",
X"83c08008",
X"5483c080",
X"0880df38",
X"893d3354",
X"73802e91",
X"3802ab05",
X"3370842a",
X"81065155",
X"74802e86",
X"38835480",
X"c1397651",
X"f4893f83",
X"c08008a0",
X"170c02bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"3371079c",
X"1c0c5278",
X"981b0c53",
X"56595781",
X"0b811734",
X"74547383",
X"c0800c99",
X"3d0d04f5",
X"3d0d7d7f",
X"617283c0",
X"98085a5d",
X"5d595c80",
X"7b0c8557",
X"75802e81",
X"e0388116",
X"33810655",
X"84577480",
X"2e81d238",
X"91397481",
X"17348639",
X"800b8117",
X"34815781",
X"c0399c16",
X"08981708",
X"31557478",
X"27833874",
X"5877802e",
X"81a93898",
X"16087083",
X"ff065657",
X"7480cf38",
X"821633ff",
X"0577892a",
X"067081ff",
X"065a5578",
X"a0387687",
X"38a01608",
X"558d39a4",
X"160851f0",
X"e93f83c0",
X"80085581",
X"7527ffa8",
X"3874a417",
X"0ca41608",
X"51f2833f",
X"83c08008",
X"5583c080",
X"08802eff",
X"893883c0",
X"800819a8",
X"170c9816",
X"0883ff06",
X"84807131",
X"51557775",
X"27833877",
X"557483ff",
X"ff065498",
X"160883ff",
X"0653a816",
X"08527957",
X"7b83387b",
X"5776518a",
X"8d3f83c0",
X"8008fed0",
X"38981608",
X"1598170c",
X"741a7876",
X"317c0817",
X"7d0c595a",
X"fed33980",
X"577683c0",
X"800c8d3d",
X"0d04fa3d",
X"0d7883c0",
X"98085556",
X"85557380",
X"2e81e138",
X"81143381",
X"06538455",
X"72802e81",
X"d3389c14",
X"08537276",
X"27833872",
X"56981408",
X"57800b98",
X"150c7580",
X"2e81b738",
X"82143370",
X"892b5653",
X"76802eb5",
X"387452ff",
X"1651bd98",
X"3f83c080",
X"08ff1876",
X"54705358",
X"53bd893f",
X"83c08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed83f83",
X"c0800853",
X"810b83c0",
X"8008278b",
X"38881408",
X"83c08008",
X"26883880",
X"0b811534",
X"b03983c0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc73f",
X"83c08008",
X"8c3883c0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683c0",
X"800805a8",
X"150c8055",
X"7483c080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83c09808",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1d13f",
X"83c08008",
X"5583c080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef7",
X"3f83c080",
X"0888170c",
X"7551efa8",
X"3f83c080",
X"08557483",
X"c0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683c0",
X"9808802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f73f83c0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"86983f83",
X"c0800841",
X"83c08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"ede13f83",
X"c0800841",
X"83c08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"83a53f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f23f83c0",
X"80088332",
X"70307072",
X"079f2c83",
X"c0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"81b13f75",
X"83c0800c",
X"9e3d0d04",
X"fd3d0d75",
X"77535473",
X"33517089",
X"38713351",
X"70802ea1",
X"38733372",
X"33525372",
X"71278538",
X"ff519439",
X"70732785",
X"3881518b",
X"39811481",
X"135354d3",
X"39805170",
X"83c0800c",
X"853d0d04",
X"fd3d0d75",
X"77545472",
X"337081ff",
X"06525270",
X"802ea338",
X"7181ff06",
X"8114ffbf",
X"12535452",
X"70992689",
X"38a01270",
X"81ff0653",
X"51717470",
X"81055634",
X"d2398074",
X"34853d0d",
X"04ffbd3d",
X"0d80c63d",
X"0852a53d",
X"705254ff",
X"b33f80c7",
X"3d085285",
X"3d705253",
X"ffa63f72",
X"527351fe",
X"df3f80c5",
X"3d0d04fe",
X"3d0d7476",
X"53537170",
X"81055333",
X"51707370",
X"81055534",
X"70f03884",
X"3d0d04fe",
X"3d0d7452",
X"80723352",
X"5370732e",
X"8d388112",
X"81147133",
X"53545270",
X"f5387283",
X"c0800c84",
X"3d0d04fc",
X"3d0d7655",
X"7483c3a8",
X"082eaf38",
X"80537451",
X"87c13f83",
X"c0800881",
X"ff06ff14",
X"7081ff06",
X"7230709f",
X"2a515255",
X"53547280",
X"2e843871",
X"dd3873fe",
X"387483c3",
X"a80c863d",
X"0d04ff3d",
X"0dff0b83",
X"c3a80c84",
X"a53f8151",
X"87853f83",
X"c0800881",
X"ff065271",
X"ee3881d3",
X"3f7183c0",
X"800c833d",
X"0d04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"823f7280",
X"2ea03883",
X"c3bc1433",
X"75708105",
X"57348114",
X"7083ffff",
X"06ff1570",
X"83ffff06",
X"56525552",
X"dd39800b",
X"83c0800c",
X"863d0d04",
X"fc3d0d76",
X"787a1156",
X"53558053",
X"71742e93",
X"38721551",
X"703383c3",
X"bc133481",
X"12811454",
X"52ea3980",
X"0b83c080",
X"0c863d0d",
X"04fd3d0d",
X"905483c3",
X"a8085186",
X"f43f83c0",
X"800881ff",
X"06ff1571",
X"30713070",
X"73079f2a",
X"729f2a06",
X"52555255",
X"5372db38",
X"853d0d04",
X"803d0d83",
X"c3b40810",
X"83c3ac08",
X"079080a8",
X"0c823d0d",
X"04800b83",
X"c3b40ce4",
X"3f04810b",
X"83c3b40c",
X"db3f04ed",
X"3f047183",
X"c3b00c04",
X"803d0d80",
X"51f43f81",
X"0b83c3b4",
X"0c810b83",
X"c3ac0cff",
X"bb3f823d",
X"0d04803d",
X"0d723070",
X"74078025",
X"83c3ac0c",
X"51ffa53f",
X"823d0d04",
X"803d0d02",
X"8b053390",
X"80a40c90",
X"80a80870",
X"81065151",
X"70f53890",
X"80a40870",
X"81ff0683",
X"c0800c51",
X"823d0d04",
X"803d0d81",
X"ff51d13f",
X"83c08008",
X"81ff0683",
X"c0800c82",
X"3d0d0480",
X"3d0d7390",
X"2b730790",
X"80b40c82",
X"3d0d0404",
X"fb3d0d78",
X"0284059f",
X"05337098",
X"2b555755",
X"7280259b",
X"387580ff",
X"06568052",
X"80f751e0",
X"3f83c080",
X"0881ff06",
X"54738126",
X"80ff3880",
X"51fee73f",
X"ffa23f81",
X"51fedf3f",
X"ff9a3f75",
X"51feed3f",
X"74982a51",
X"fee63f74",
X"902a7081",
X"ff065253",
X"feda3f74",
X"882a7081",
X"ff065253",
X"fece3f74",
X"81ff0651",
X"fec63f81",
X"557580c0",
X"2e098106",
X"86388195",
X"558d3975",
X"80c82e09",
X"81068438",
X"81875574",
X"51fea53f",
X"8a55fec8",
X"3f83c080",
X"0881ff06",
X"70982b54",
X"54728025",
X"8c38ff15",
X"7081ff06",
X"565374e2",
X"387383c0",
X"800c873d",
X"0d04fa3d",
X"0dfdc53f",
X"8051fdda",
X"3f8a54fe",
X"933fff14",
X"7081ff06",
X"555373f3",
X"38737453",
X"5580c051",
X"fea63f83",
X"c0800881",
X"ff065473",
X"812e0981",
X"06829f38",
X"83aa5280",
X"c851fe8c",
X"3f83c080",
X"0881ff06",
X"5372812e",
X"09810681",
X"a8387454",
X"873d7411",
X"5456fdc8",
X"3f83c080",
X"08733481",
X"147081ff",
X"06555383",
X"7427e538",
X"029a0533",
X"5372812e",
X"09810681",
X"d938029b",
X"05335380",
X"ce905472",
X"81aa2e8d",
X"3881c739",
X"80e4518a",
X"cc3fff14",
X"5473802e",
X"81b83882",
X"0a5281e9",
X"51fda53f",
X"83c08008",
X"81ff0653",
X"72de3872",
X"5280fa51",
X"fd923f83",
X"c0800881",
X"ff065372",
X"81903872",
X"54731653",
X"fcd63f83",
X"c0800873",
X"34811470",
X"81ff0655",
X"53837427",
X"e838873d",
X"3370862a",
X"70810651",
X"54548c55",
X"7280e338",
X"845580de",
X"39745281",
X"e951fccc",
X"3f83c080",
X"0881ff06",
X"53825581",
X"e9568173",
X"27863873",
X"5580c156",
X"80ce9054",
X"8a3980e4",
X"5189be3f",
X"ff145473",
X"802ea938",
X"80527551",
X"fc9a3f83",
X"c0800881",
X"ff065372",
X"e1388480",
X"5280d051",
X"fc863f83",
X"c0800881",
X"ff065372",
X"802e8338",
X"80557483",
X"c3b83480",
X"51fb873f",
X"fbc23f88",
X"3d0d04fb",
X"3d0d7754",
X"800b83c3",
X"b8337083",
X"2a708106",
X"51555755",
X"72752e09",
X"81068538",
X"73892b54",
X"735280d1",
X"51fbbd3f",
X"83c08008",
X"81ff0653",
X"72bd3882",
X"b8c054fb",
X"833f83c0",
X"800881ff",
X"06537281",
X"ff2e0981",
X"068938ff",
X"145473e7",
X"389f3972",
X"81fe2e09",
X"81069638",
X"83c7bc52",
X"83c3bc51",
X"faed3ffa",
X"d33ffad0",
X"3f833981",
X"558051fa",
X"893ffac4",
X"3f7481ff",
X"0683c080",
X"0c873d0d",
X"04fb3d0d",
X"7783c3bc",
X"56548151",
X"f9ec3f83",
X"c3b83370",
X"832a7081",
X"06515456",
X"72853873",
X"892b5473",
X"5280d851",
X"fab63f83",
X"c0800881",
X"ff065372",
X"80e43881",
X"ff51f9d4",
X"3f81fe51",
X"f9ce3f84",
X"80537470",
X"81055633",
X"51f9c13f",
X"ff137083",
X"ffff0651",
X"5372eb38",
X"7251f9b0",
X"3f7251f9",
X"ab3ff9d0",
X"3f83c080",
X"089f0653",
X"a7885472",
X"852e8c38",
X"993980e4",
X"5186f63f",
X"ff1454f9",
X"b33f83c0",
X"800881ff",
X"2e843873",
X"e9388051",
X"f8e43ff9",
X"9f3f800b",
X"83c0800c",
X"873d0d04",
X"7183c7c0",
X"0c888080",
X"0b83c7bc",
X"0c848080",
X"0b83c7c4",
X"0c04fd3d",
X"0d777017",
X"557705ff",
X"1a535371",
X"ff2e9438",
X"73708105",
X"55335170",
X"73708105",
X"5534ff12",
X"52e93985",
X"3d0d04fc",
X"3d0d87a6",
X"81557433",
X"83c7c834",
X"a05483a0",
X"805383c7",
X"c0085283",
X"c7bc0851",
X"ffb83fa0",
X"5483a480",
X"5383c7c0",
X"085283c7",
X"bc0851ff",
X"a53f9054",
X"83a88053",
X"83c7c008",
X"5283c7bc",
X"0851ff92",
X"3fa05380",
X"5283c7c4",
X"0883a080",
X"055185ce",
X"3fa05380",
X"5283c7c4",
X"0883a480",
X"055185be",
X"3f905380",
X"5283c7c4",
X"0883a880",
X"055185ae",
X"3fff7534",
X"83a08054",
X"805383c7",
X"c0085283",
X"c7c40851",
X"fecc3f80",
X"d0805483",
X"b0805383",
X"c7c00852",
X"83c7c408",
X"51feb73f",
X"86e13fa2",
X"54805383",
X"c7c4088c",
X"80055281",
X"dbf851fe",
X"a13f860b",
X"87a88334",
X"800b87a8",
X"8234800b",
X"87a09a34",
X"af0b87a0",
X"9634bf0b",
X"87a09734",
X"800b87a0",
X"98349f0b",
X"87a09934",
X"800b87a0",
X"9b34e00b",
X"87a88934",
X"a20b87a8",
X"8034830b",
X"87a48f34",
X"820b87a8",
X"8134863d",
X"0d04fd3d",
X"0d83a080",
X"54805383",
X"c7c40852",
X"83c7c008",
X"51fdbf3f",
X"80d08054",
X"83b08053",
X"83c7c408",
X"5283c7c0",
X"0851fdaa",
X"3fa05483",
X"a0805383",
X"c7c40852",
X"83c7c008",
X"51fd973f",
X"a05483a4",
X"805383c7",
X"c4085283",
X"c7c00851",
X"fd843f90",
X"5483a880",
X"5383c7c4",
X"085283c7",
X"c00851fc",
X"f13f83c7",
X"c83387a6",
X"8134853d",
X"0d04803d",
X"0d908090",
X"08810683",
X"c0800c82",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe067607",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"812c8106",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fd06",
X"76100772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087082",
X"2cbf0683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fe8306",
X"76822b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"882c8706",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f1ff",
X"0676882b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"708b2cbf",
X"0683c080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870f8",
X"8fff0676",
X"8b2b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087091",
X"2cbf0683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fc87ff",
X"ff067691",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870992c",
X"810683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"ffbf0a06",
X"76992b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80800870",
X"882c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"70892c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708a2c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708b",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8c2cbf06",
X"83c0800c",
X"51823d0d",
X"04fe3d0d",
X"7481e629",
X"872a9080",
X"a00c843d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"81055434",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727084",
X"05540cff",
X"1151f039",
X"843d0d04",
X"fe3d0d84",
X"80805380",
X"5288800a",
X"51ffb33f",
X"81808053",
X"80528280",
X"0a51c63f",
X"843d0d04",
X"803d0d81",
X"51fbfc3f",
X"72802e90",
X"388051fd",
X"fe3fcd3f",
X"83c7cc33",
X"51fdf43f",
X"8151fc8d",
X"3f8051fc",
X"883f8051",
X"fbd93f82",
X"3d0d04fd",
X"3d0d7552",
X"805480ff",
X"72258838",
X"810bff80",
X"135354ff",
X"bf125170",
X"99268638",
X"e012529e",
X"39ff9f12",
X"51997127",
X"9538d012",
X"e0137054",
X"54518971",
X"2788388f",
X"73278338",
X"80527380",
X"2e853881",
X"80125271",
X"81ff0683",
X"c0800c85",
X"3d0d0480",
X"3d0d84d8",
X"c0518071",
X"70810553",
X"347084e0",
X"c02e0981",
X"06f03882",
X"3d0d04fe",
X"3d0d0297",
X"053351ff",
X"863f83c0",
X"800881ff",
X"0683c7d0",
X"08545280",
X"73249b38",
X"83c89008",
X"137283c8",
X"94080753",
X"53717334",
X"83c7d008",
X"810583c7",
X"d00c843d",
X"0d04fa3d",
X"0d82800a",
X"1b558057",
X"883dfc05",
X"54795374",
X"527851cb",
X"d33f883d",
X"0d04fe3d",
X"0d83c7e8",
X"08527451",
X"d2b73f83",
X"c080088c",
X"38765375",
X"5283c7e8",
X"0851c73f",
X"843d0d04",
X"fe3d0d83",
X"c7e80853",
X"75527451",
X"ccf63f83",
X"c080088d",
X"38775376",
X"5283c7e8",
X"0851ffa2",
X"3f843d0d",
X"04fe3d0d",
X"83c7e808",
X"51cbea3f",
X"83c08008",
X"8180802e",
X"09810688",
X"3883c180",
X"80539b39",
X"83c7e808",
X"51cbce3f",
X"83c08008",
X"80d0802e",
X"09810693",
X"3883c1b0",
X"805383c0",
X"80085283",
X"c7e80851",
X"fed83f84",
X"3d0d0480",
X"3d0df9e4",
X"3f83c080",
X"08842981",
X"dc9c0570",
X"0883c080",
X"0c51823d",
X"0d04ed3d",
X"0d804480",
X"43804280",
X"4180705a",
X"5bfdd03f",
X"800b83c7",
X"d00c800b",
X"83c8940c",
X"81d9ec51",
X"c6b83f81",
X"800b83c8",
X"940c81d9",
X"f051c6aa",
X"3f80d00b",
X"83c7d00c",
X"7830707a",
X"07802570",
X"872b83c8",
X"940c5155",
X"f8d53f83",
X"c0800852",
X"81d9f851",
X"c6843f80",
X"f80b83c7",
X"d00c7881",
X"32703070",
X"72078025",
X"70872b83",
X"c8940c51",
X"5656feef",
X"3f83c080",
X"085281da",
X"8451c5da",
X"3f81a00b",
X"83c7d00c",
X"78823270",
X"30707207",
X"80257087",
X"2b83c894",
X"0c515683",
X"c7e80852",
X"56c6f43f",
X"83c08008",
X"5281da8c",
X"51c5ab3f",
X"81f00b83",
X"c7d00c81",
X"0b83c7d4",
X"5b5883c7",
X"d0088219",
X"7a327030",
X"70720780",
X"2570872b",
X"83c8940c",
X"51578e3d",
X"7055ff1b",
X"54575757",
X"9aa73f79",
X"7084055b",
X"0851c6ab",
X"3f745483",
X"c0800853",
X"775281da",
X"9451c4de",
X"3fa81783",
X"c7d00c81",
X"18587785",
X"2e098106",
X"ffb03883",
X"900b83c7",
X"d00c7887",
X"32703070",
X"72078025",
X"70872b83",
X"c8940c51",
X"5656f7fb",
X"3f81daa4",
X"5583c080",
X"08802e8e",
X"3883c7e4",
X"0851c5d7",
X"3f83c080",
X"08557452",
X"81daac51",
X"c48c3f83",
X"e00b83c7",
X"d00c7888",
X"32703070",
X"72078025",
X"70872b83",
X"c8940c51",
X"5781dab8",
X"5255c3ea",
X"3f868da0",
X"51f8f63f",
X"8052913d",
X"7052559b",
X"db3f8352",
X"74519bd4",
X"3f635574",
X"82fc3861",
X"19597880",
X"25853874",
X"59903988",
X"79258538",
X"88598739",
X"78882682",
X"db387882",
X"2b5581d4",
X"f4150804",
X"f5e93f83",
X"c0800861",
X"57557581",
X"2e098106",
X"893883c0",
X"80081055",
X"903975ff",
X"2e098106",
X"883883c0",
X"8008812c",
X"55907525",
X"85389055",
X"88397480",
X"24833881",
X"557451f5",
X"c33f8290",
X"39f5d53f",
X"83c08008",
X"61055574",
X"80258538",
X"80558839",
X"87752583",
X"38875574",
X"51f5ce3f",
X"81ee3960",
X"87386280",
X"2e81e538",
X"83c0b408",
X"83c0b00c",
X"8bdf0b83",
X"c0b80c83",
X"c7e80851",
X"ffb4ee3f",
X"fadf3f81",
X"c7396056",
X"80762599",
X"388af80b",
X"83c0b80c",
X"83c7c815",
X"70085255",
X"ffb4ce3f",
X"74085291",
X"39758025",
X"913883c7",
X"c8150851",
X"c3bf3f80",
X"52fd1951",
X"b8396280",
X"2e818d38",
X"83c7c815",
X"700883c7",
X"d408720c",
X"83c7d40c",
X"fd1a7053",
X"51558c94",
X"3f83c080",
X"08568051",
X"8c8a3f83",
X"c0800852",
X"745188a2",
X"3f755280",
X"51889b3f",
X"80d63960",
X"55807525",
X"b83883c0",
X"bc0883c0",
X"b00c8bdf",
X"0b83c0b8",
X"0c83c7e4",
X"0851ffb3",
X"d83f83c7",
X"e40851ff",
X"b0f23f83",
X"c0800881",
X"ff067052",
X"55f4d93f",
X"74802e9c",
X"388155a0",
X"39748025",
X"933883c7",
X"e40851c2",
X"b03f8051",
X"f4be3f84",
X"39628738",
X"7a802efa",
X"84388055",
X"7483c080",
X"0c953d0d",
X"04fe3d0d",
X"83c88051",
X"80f3e83f",
X"83c7f051",
X"80f3e03f",
X"f4da3f83",
X"c0800880",
X"2e863880",
X"51818b39",
X"f4df3f83",
X"c0800880",
X"ff38f4ff",
X"3f83c080",
X"08802eb9",
X"388151f2",
X"8e3f8051",
X"f4953fef",
X"823f800b",
X"83c7d00c",
X"f99c3f83",
X"c0800853",
X"ff0b83c7",
X"d00cf0ee",
X"3f7280cc",
X"3883c7cc",
X"3351f3ef",
X"3f7251f1",
X"de3f80c1",
X"39f4a73f",
X"83c08008",
X"802eb638",
X"8151f1cb",
X"3f8051f3",
X"d23feebf",
X"3f8af80b",
X"83c0b80c",
X"83c7d408",
X"51ffb1f9",
X"3fff0b83",
X"c7d00cf0",
X"a93f83c7",
X"d4085280",
X"5186873f",
X"8151f598",
X"3f843d0d",
X"04fb3d0d",
X"805283c8",
X"805180e2",
X"ee3f8152",
X"83c7f051",
X"80e2e43f",
X"800b83c7",
X"cc349080",
X"80528684",
X"808051c4",
X"c53f83c0",
X"80088193",
X"3889be3f",
X"81ddfc51",
X"c9853f83",
X"c0800855",
X"9c800a54",
X"80c08053",
X"81dac052",
X"83c08008",
X"51f6d93f",
X"83c7e808",
X"5381dad0",
X"527451c3",
X"cf3f83c0",
X"80088438",
X"f6e73f83",
X"c7ec0853",
X"81dadc52",
X"7451c3b8",
X"3f83c080",
X"08b53887",
X"3dfc0554",
X"84808053",
X"86a88080",
X"5283c7ec",
X"0851c1c4",
X"3f83c080",
X"08933875",
X"8480802e",
X"09810689",
X"38810b83",
X"c7cc3487",
X"39800b83",
X"c7cc3483",
X"c7cc3351",
X"f1e93f81",
X"51f3d53f",
X"92fa3f81",
X"51f3cd3f",
X"8151fd81",
X"3ffa3983",
X"c08c0802",
X"83c08c0c",
X"fb3d0d02",
X"81dae80b",
X"83c0b40c",
X"81daec0b",
X"83c0ac0c",
X"81daf00b",
X"83c0bc0c",
X"83c08c08",
X"fc050c80",
X"0b83c7d4",
X"0b83c08c",
X"08f8050c",
X"83c08c08",
X"f4050cc1",
X"d53f83c0",
X"80088605",
X"fc0683c0",
X"8c08f005",
X"0c0283c0",
X"8c08f005",
X"08310d83",
X"3d7083c0",
X"8c08f805",
X"08708405",
X"83c08c08",
X"f8050c0c",
X"51ffbe9d",
X"3f83c08c",
X"08f40508",
X"810583c0",
X"8c08f405",
X"0c83c08c",
X"08f40508",
X"872e0981",
X"06ffac38",
X"86948080",
X"51eae93f",
X"ff0b83c7",
X"d00c800b",
X"83c8940c",
X"84d8c00b",
X"83c8900c",
X"8151ee93",
X"3f8151ee",
X"b83f8051",
X"eeb33f81",
X"51eed93f",
X"8151efae",
X"3f8251ee",
X"fc3f8051",
X"efd23f80",
X"51effc3f",
X"80d0e752",
X"8051ffbb",
X"d63ffccd",
X"3f83c08c",
X"08fc0508",
X"0d800b83",
X"c0800c87",
X"3d0d83c0",
X"8c0c0480",
X"3d0d81ff",
X"51800b83",
X"c8a01234",
X"ff115170",
X"f438823d",
X"0d04ff3d",
X"0d737033",
X"53518111",
X"33713471",
X"81123483",
X"3d0d04fb",
X"3d0d7779",
X"56568070",
X"71555552",
X"717525ac",
X"38721670",
X"33701470",
X"81ff0655",
X"51515171",
X"74278938",
X"81127081",
X"ff065351",
X"71811470",
X"83ffff06",
X"55525474",
X"7324d638",
X"7183c080",
X"0c873d0d",
X"04fb3d0d",
X"7756ffb5",
X"823f83c0",
X"8008802e",
X"f53883ca",
X"bc088605",
X"7081ff06",
X"5253ffb3",
X"823f810b",
X"9088d434",
X"9088d433",
X"7081ff06",
X"51537286",
X"38f9da3f",
X"ef398055",
X"74167582",
X"2b545490",
X"88c01333",
X"74348115",
X"5574852e",
X"098106e8",
X"38810b90",
X"88d43475",
X"3383c8a0",
X"34811633",
X"83c8a134",
X"82163383",
X"c8a23483",
X"163383c8",
X"a3348452",
X"83c8a051",
X"febd3f83",
X"c0800881",
X"ff068417",
X"33575372",
X"762e0981",
X"068d38ff",
X"b3ae3f83",
X"c0800880",
X"2e9a3883",
X"cabc08a8",
X"2e098106",
X"8938860b",
X"83cabc0c",
X"8739a80b",
X"83cabc0c",
X"80e451ee",
X"ac3f873d",
X"0d04f43d",
X"0d7e6059",
X"55805d80",
X"75822b71",
X"83cac012",
X"0c83cad4",
X"175b5b57",
X"76793477",
X"772e83b8",
X"38765277",
X"51ffbce4",
X"3f8e3dfc",
X"05549053",
X"83caa852",
X"7751ffbc",
X"9f3f7c56",
X"75902e09",
X"81068394",
X"3883caa8",
X"51fd973f",
X"83caaa51",
X"fd903f83",
X"caac51fd",
X"893f7683",
X"cab80c77",
X"51ffb9eb",
X"3f81d8fc",
X"5283c080",
X"0851ffa9",
X"913f83c0",
X"8008812e",
X"09810680",
X"d4387683",
X"cad00c82",
X"0b83caa8",
X"34ff960b",
X"83caa934",
X"7751ffbc",
X"b03f83c0",
X"80085583",
X"c0800877",
X"25883883",
X"c080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583caaa",
X"347483ca",
X"ab347683",
X"caac34ff",
X"800b83ca",
X"ad348190",
X"3983caa8",
X"3383caa9",
X"3371882b",
X"07565b74",
X"83ffff2e",
X"09810680",
X"e838fe80",
X"0b83cad0",
X"0c810b83",
X"cab80cff",
X"0b83caa8",
X"34ff0b83",
X"caa93477",
X"51ffbbbd",
X"3f83c080",
X"0883cad8",
X"0c83c080",
X"085583c0",
X"80088025",
X"883883c0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83caaa34",
X"7483caab",
X"347683ca",
X"ac34ff80",
X"0b83caad",
X"34810b83",
X"cab734a5",
X"39748596",
X"2e098106",
X"80fe3875",
X"83cad00c",
X"7751ffba",
X"f13f83ca",
X"b73383c0",
X"80080755",
X"7483cab7",
X"3483cab7",
X"33810655",
X"74802e83",
X"38845783",
X"caac3383",
X"caad3371",
X"882b0756",
X"5c748180",
X"2e098106",
X"a13883ca",
X"aa3383ca",
X"ab337188",
X"2b07565b",
X"ad807527",
X"87387682",
X"07579c39",
X"76810757",
X"96397482",
X"802e0981",
X"06873876",
X"83075787",
X"397481ff",
X"268a3877",
X"83cac01b",
X"0c767934",
X"8e3d0d04",
X"803d0d72",
X"842983ca",
X"c0057008",
X"83c0800c",
X"51823d0d",
X"04fe3d0d",
X"800b83ca",
X"a40c800b",
X"83caa00c",
X"ff0b83c8",
X"9c0ca80b",
X"83cabc0c",
X"ae51ffad",
X"ce3f800b",
X"83cac054",
X"52807370",
X"8405550c",
X"81125271",
X"842e0981",
X"06ef3884",
X"3d0d04fe",
X"3d0d7402",
X"84059605",
X"22535371",
X"802e9738",
X"72708105",
X"543351ff",
X"add83fff",
X"127083ff",
X"ff065152",
X"e639843d",
X"0d04fe3d",
X"0d029205",
X"225382ac",
X"51e9be3f",
X"80c351ff",
X"adb43f81",
X"9651e9b1",
X"3f725283",
X"c8a051ff",
X"b23f7252",
X"83c8a051",
X"f8f13f83",
X"c0800881",
X"ff0651ff",
X"ad903f84",
X"3d0d04ff",
X"b13d0d80",
X"d13df805",
X"51f99a3f",
X"83caa408",
X"810583ca",
X"a40c80cf",
X"3d33cf11",
X"7081ff06",
X"51565674",
X"832688ed",
X"38758f06",
X"ff055675",
X"83c89c08",
X"2e9b3875",
X"83269638",
X"7583c89c",
X"0c758429",
X"83cac005",
X"70085355",
X"7551fa96",
X"3f807624",
X"88c93875",
X"842983ca",
X"c0055574",
X"08802e88",
X"ba3883c8",
X"9c088429",
X"83cac005",
X"70080288",
X"0582b905",
X"33525b55",
X"7480d22e",
X"84b13874",
X"80d22490",
X"3874bf2e",
X"9c387480",
X"d02e81d7",
X"3887f839",
X"7480d32e",
X"80d23874",
X"80d72e81",
X"c63887e7",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055656",
X"ffac8c3f",
X"80c151ff",
X"abc43ff6",
X"ea3f860b",
X"83c8a034",
X"815283c8",
X"a051ffac",
X"e73f8151",
X"fde43f74",
X"8938860b",
X"83cabc0c",
X"8739a80b",
X"83cabc0c",
X"ffabd83f",
X"80c151ff",
X"ab903ff6",
X"b63f900b",
X"83cab733",
X"81065656",
X"74802e83",
X"38985683",
X"caac3383",
X"caad3371",
X"882b0756",
X"59748180",
X"2e098106",
X"9c3883ca",
X"aa3383ca",
X"ab337188",
X"2b075657",
X"ad807527",
X"8c387581",
X"80075685",
X"3975a007",
X"567583c8",
X"a034ff0b",
X"83c8a134",
X"e00b83c8",
X"a234800b",
X"83c8a334",
X"845283c8",
X"a051ffab",
X"db3f8451",
X"869e3902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"5659ffaa",
X"ca3f7951",
X"ffb5b73f",
X"83c08008",
X"802e8b38",
X"80ce51ff",
X"a9f43f85",
X"f23980c1",
X"51ffa9ea",
X"3fffaadf",
X"3fffa992",
X"3f83cad0",
X"08588375",
X"259b3883",
X"caac3383",
X"caad3371",
X"882b07fc",
X"1771297a",
X"05838005",
X"5a51578d",
X"39748180",
X"2918ff80",
X"05588180",
X"57805676",
X"762e9338",
X"ffa9c33f",
X"83c08008",
X"83c8a017",
X"34811656",
X"ea39ffa9",
X"b13f83c0",
X"800881ff",
X"06775383",
X"c8a05256",
X"f4d93f83",
X"c0800881",
X"ff065575",
X"752e0981",
X"06818a38",
X"ffa9b03f",
X"80c151ff",
X"a8e83fff",
X"a9dd3f77",
X"527951ff",
X"b3c63f80",
X"5e80d13d",
X"fdf40554",
X"765383c8",
X"a0527951",
X"ffb1d33f",
X"0282b905",
X"33558158",
X"7480d72e",
X"098106bd",
X"3880d13d",
X"fdf00554",
X"76538f3d",
X"70537a52",
X"59ffb2d8",
X"3f805676",
X"762ea238",
X"751983c8",
X"a0173371",
X"33707232",
X"70307080",
X"2570307e",
X"06811d5d",
X"5e515151",
X"525b55db",
X"3982ac51",
X"e3f73f77",
X"802e8638",
X"80c35184",
X"3980ce51",
X"ffa7e33f",
X"ffa8d83f",
X"ffa78b3f",
X"83dd3902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"59558070",
X"5d59ffa7",
X"fe3f80c1",
X"51ffa7b6",
X"3f83cab8",
X"08792e82",
X"de3883ca",
X"d80880fc",
X"055580fd",
X"52745187",
X"bb3f83c0",
X"80085b77",
X"8224b238",
X"ff187087",
X"2b83ffff",
X"800681dc",
X"bc0583c8",
X"a0595755",
X"81805575",
X"70810557",
X"33777081",
X"055934ff",
X"157081ff",
X"06515574",
X"ea38828d",
X"397782e8",
X"2e81ab38",
X"7782e92e",
X"09810681",
X"b23881da",
X"f451ffad",
X"b93f7858",
X"77873270",
X"30707207",
X"80257a8a",
X"32703070",
X"72078025",
X"73075354",
X"5a515755",
X"75802e97",
X"38787826",
X"9238a00b",
X"83c8a01a",
X"34811970",
X"81ff065a",
X"55eb3981",
X"187081ff",
X"0659558a",
X"7827ffbc",
X"388f5883",
X"c89b1833",
X"83c8a019",
X"34ff1870",
X"81ff0659",
X"55778426",
X"ea389058",
X"800b83c8",
X"a0193481",
X"187081ff",
X"0670982b",
X"52595574",
X"8025e938",
X"80c6557a",
X"858f2484",
X"3880c255",
X"7483c8a0",
X"3480f10b",
X"83c8a334",
X"810b83c8",
X"a4347a83",
X"c8a1347a",
X"882c5574",
X"83c8a234",
X"80cb3982",
X"f0782580",
X"c4387780",
X"fd29fd97",
X"d3055279",
X"51ffaff4",
X"3f80d13d",
X"fdec0554",
X"80fd5383",
X"c8a05279",
X"51ffafac",
X"3f7b8119",
X"59567580",
X"fc248338",
X"78587788",
X"2c557483",
X"c99d3477",
X"83c99e34",
X"7583c99f",
X"34818059",
X"80cc3983",
X"cad00857",
X"8378259b",
X"3883caac",
X"3383caad",
X"3371882b",
X"07fc1a71",
X"29790583",
X"80055951",
X"598d3977",
X"81802917",
X"ff800557",
X"81805976",
X"527951ff",
X"af823f80",
X"d13dfdec",
X"05547853",
X"83c8a052",
X"7951ffae",
X"bb3f7851",
X"f6b83fff",
X"a4f53fff",
X"a3a83f8b",
X"3983caa0",
X"08810583",
X"caa00c80",
X"d13d0d04",
X"f6d93ffc",
X"39fc3d0d",
X"76787184",
X"2983cac0",
X"05700851",
X"53535370",
X"9e3880ce",
X"723480cf",
X"0b811334",
X"80ce0b82",
X"133480c5",
X"0b831334",
X"70841334",
X"80e73983",
X"cad41333",
X"5480d272",
X"3473822a",
X"70810651",
X"5180cf53",
X"70843880",
X"d7537281",
X"1334a00b",
X"82133473",
X"83065170",
X"812e9e38",
X"70812488",
X"3870802e",
X"8f389f39",
X"70822e92",
X"3870832e",
X"92389339",
X"80d8558e",
X"3980d355",
X"893980cd",
X"55843980",
X"c4557483",
X"133480c4",
X"0b841334",
X"800b8513",
X"34863d0d",
X"04fc3d0d",
X"76558075",
X"0c800b84",
X"160c800b",
X"88160c80",
X"0b8c160c",
X"83c88051",
X"80dcc43f",
X"83c7f051",
X"80dcbc3f",
X"87a68033",
X"7081ff06",
X"5152de80",
X"3f71812a",
X"81327281",
X"32718106",
X"71810631",
X"84180c54",
X"5471832a",
X"81327282",
X"2a813271",
X"81067181",
X"0631770c",
X"535387a0",
X"90337009",
X"81068817",
X"0c5283c0",
X"8008802e",
X"80c23883",
X"c0800881",
X"2a708106",
X"83c08008",
X"81063184",
X"170c5283",
X"c0800883",
X"2a83c080",
X"08822a71",
X"81067181",
X"0631770c",
X"535383c0",
X"8008842a",
X"81068816",
X"0c83c080",
X"08852a81",
X"068c160c",
X"863d0d04",
X"fe3d0d74",
X"76545271",
X"51febe3f",
X"72812ea2",
X"38817326",
X"8d387282",
X"2ea83872",
X"832e9c38",
X"e6397108",
X"e2388412",
X"08dd3888",
X"1208d838",
X"a5398812",
X"08812e9e",
X"38913988",
X"1208812e",
X"95387108",
X"91388412",
X"088c388c",
X"1208812e",
X"098106ff",
X"b238843d",
X"0d04fc3d",
X"0d767853",
X"54815380",
X"55873971",
X"10731054",
X"52737226",
X"5172802e",
X"a7387080",
X"2e863871",
X"8025e838",
X"72802e98",
X"38717426",
X"89387372",
X"31757407",
X"56547281",
X"2a72812a",
X"5353e539",
X"73517883",
X"38745170",
X"83c0800c",
X"863d0d04",
X"fe3d0d80",
X"53755274",
X"51ffa33f",
X"843d0d04",
X"fe3d0d81",
X"53755274",
X"51ff933f",
X"843d0d04",
X"fb3d0d77",
X"79555580",
X"56747625",
X"86387430",
X"55815673",
X"80258838",
X"73307681",
X"32575480",
X"53735274",
X"51fee73f",
X"83c08008",
X"5475802e",
X"873883c0",
X"80083054",
X"7383c080",
X"0c873d0d",
X"04fa3d0d",
X"787a5755",
X"80577477",
X"25863874",
X"30558157",
X"759f2c54",
X"81537574",
X"32743152",
X"7451feaa",
X"3f83c080",
X"08547680",
X"2e873883",
X"c0800830",
X"547383c0",
X"800c883d",
X"0d04fb3d",
X"0d780284",
X"059f0533",
X"5556800b",
X"81d78456",
X"5381732b",
X"74065271",
X"802e8338",
X"81527470",
X"82055622",
X"7073902b",
X"0790809c",
X"0c518113",
X"5372882e",
X"098106d9",
X"38805383",
X"cae01333",
X"517081ff",
X"2eb23870",
X"1081d5a4",
X"05702255",
X"51807317",
X"70337010",
X"81d5a405",
X"70225151",
X"51525273",
X"712e9138",
X"81125271",
X"862e0981",
X"06f13873",
X"90809c0c",
X"81135372",
X"862e0981",
X"06ffb838",
X"80537216",
X"70335151",
X"7081ff2e",
X"94387010",
X"81d5a405",
X"70227084",
X"80800790",
X"809c0c51",
X"51811353",
X"72862e09",
X"8106d738",
X"80537216",
X"51703383",
X"cae01434",
X"81135372",
X"862e0981",
X"06ec3887",
X"3d0d0404",
X"ff3d0d74",
X"0284058f",
X"05335252",
X"70883871",
X"9080940c",
X"8e397081",
X"2e098106",
X"86387190",
X"80980c83",
X"3d0d04fb",
X"3d0d029f",
X"05337998",
X"2b70982c",
X"7c982b70",
X"982c83ca",
X"fc157033",
X"70982b70",
X"982c5158",
X"5c5a5155",
X"51545470",
X"732e0981",
X"06943883",
X"cadc1433",
X"70982b70",
X"982c5152",
X"5670722e",
X"b1387275",
X"347183ca",
X"dc153483",
X"cadd3383",
X"cafd3371",
X"982b7190",
X"2b0783ca",
X"dc337088",
X"2b720783",
X"cafc3371",
X"079080b8",
X"0c525953",
X"5452873d",
X"0d04fe3d",
X"0d748111",
X"33713371",
X"882b0783",
X"c0800c53",
X"51843d0d",
X"0483cae8",
X"3383c080",
X"0c04f53d",
X"0d02bb05",
X"33028405",
X"bf053302",
X"880580c3",
X"0533028c",
X"0580c605",
X"22665c5a",
X"5e5c567a",
X"557b5489",
X"53a1527d",
X"5180d0c0",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8d3d0d04",
X"83c08c08",
X"0283c08c",
X"0cf53d0d",
X"83c08c08",
X"88050883",
X"c08c088f",
X"053383c0",
X"8c089205",
X"22028c05",
X"73900583",
X"c08c08e8",
X"050c83c0",
X"8c08f805",
X"0c83c08c",
X"08f0050c",
X"83c08c08",
X"ec050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"f0050883",
X"c08c08e0",
X"050c83c0",
X"8c08fc05",
X"0c83c08c",
X"08f00508",
X"89278a38",
X"890b83c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"860587ff",
X"fc0683c0",
X"8c08e005",
X"0c0283c0",
X"8c08e005",
X"08310d85",
X"3d705583",
X"c08c08ec",
X"05085483",
X"c08c08f0",
X"05085383",
X"c08c08f4",
X"05085283",
X"c08c08e4",
X"050c80d9",
X"f23f83c0",
X"800881ff",
X"0683c08c",
X"08e40508",
X"83c08c08",
X"ec050c83",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08802e8c",
X"3883c08c",
X"08f80508",
X"0d89c839",
X"83c08c08",
X"f0050880",
X"2e89a638",
X"83c08c08",
X"ec050881",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"842ea938",
X"840b83c0",
X"8c08e005",
X"082588c7",
X"3883c08c",
X"08e00508",
X"852e859b",
X"3883c08c",
X"08e00508",
X"a12e87ad",
X"3888ac39",
X"800b83c0",
X"8c08ec05",
X"08850533",
X"83c08c08",
X"e0050c83",
X"c08c08fc",
X"050c83c0",
X"8c08e005",
X"08832e09",
X"81068883",
X"3883c08c",
X"08e80508",
X"81053383",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08812687",
X"e638810b",
X"83c08c08",
X"e0050880",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08fc050c",
X"83c08c08",
X"ec050882",
X"053383c0",
X"8c08e005",
X"08870534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088b0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08e005",
X"088c0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088d0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08e005",
X"088e0523",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088a0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"08057094",
X"0508fcff",
X"ff067194",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08ec0508",
X"86053383",
X"c08c08e0",
X"050c83c0",
X"8c08f405",
X"0c83c08c",
X"08e00508",
X"83c08c08",
X"fc05082e",
X"098106b6",
X"3883c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08fc0508",
X"83c08c08",
X"e005088b",
X"053483c0",
X"8c08ec05",
X"08870533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508812e",
X"8f3883c0",
X"8c08e005",
X"08822eb7",
X"38848c39",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"820b83c0",
X"8c08e005",
X"088a0534",
X"83d93983",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c83",
X"c08c08fc",
X"050883c0",
X"8c08e005",
X"088a0534",
X"83a13983",
X"c08c08fc",
X"0508802e",
X"83953883",
X"c08c08ec",
X"05088305",
X"33830683",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08832e09",
X"810682f3",
X"3883c08c",
X"08ec0508",
X"82053370",
X"982b83c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"83c08c08",
X"e0050880",
X"2582cc38",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"83c08c08",
X"ec050886",
X"053383c0",
X"8c08e005",
X"0880d605",
X"3483c08c",
X"08e00508",
X"840583c0",
X"8c08ec05",
X"08820533",
X"8f0683c0",
X"8c08e405",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"e4050883",
X"c08c08e0",
X"05083483",
X"c08c08ec",
X"05088405",
X"3383c08c",
X"08e00508",
X"81053480",
X"0b83c08c",
X"08e00508",
X"82053483",
X"c08c08e0",
X"050808ff",
X"83ff0682",
X"800783c0",
X"8c08e005",
X"080c83c0",
X"8c08e805",
X"08810533",
X"810583c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"83c08c08",
X"e8050881",
X"05348183",
X"3983c08c",
X"08fc0508",
X"802e80f7",
X"3883c08c",
X"08ec0508",
X"86053383",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08a22e09",
X"810680d7",
X"3883c08c",
X"08ec0508",
X"88053383",
X"c08c08ec",
X"05088705",
X"33718280",
X"290583c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c52",
X"83c08c08",
X"e4050c83",
X"c08c08f4",
X"050c83c0",
X"8c08e405",
X"0883c08c",
X"08e00508",
X"88052383",
X"c08c08ec",
X"05083383",
X"c08c08f0",
X"05087131",
X"7083ffff",
X"0683c08c",
X"08f0050c",
X"83c08c08",
X"e0050c83",
X"c08c08ec",
X"05080583",
X"c08c08ec",
X"050cf6d0",
X"3983c08c",
X"08f80508",
X"0d83c08c",
X"08f00508",
X"83c08c08",
X"e0050c83",
X"c08c08f8",
X"05080d83",
X"c08c08e0",
X"050883c0",
X"800c8d3d",
X"0d83c08c",
X"0c0483c0",
X"8c080283",
X"c08c0ce6",
X"3d0d83c0",
X"8c088805",
X"08028405",
X"83c08c08",
X"e8050c83",
X"c08c08d4",
X"050c800b",
X"83cb8434",
X"83c08c08",
X"d4050890",
X"0583c08c",
X"08c0050c",
X"800b83c0",
X"8c08c005",
X"0834800b",
X"83c08c08",
X"c0050881",
X"0534800b",
X"83c08c08",
X"c4050c83",
X"c08c08c4",
X"050880d8",
X"2983c08c",
X"08c00508",
X"0583c08c",
X"08ffb405",
X"0c800b83",
X"c08c08ff",
X"b4050880",
X"d8050c83",
X"c08c08ff",
X"b4050884",
X"0583c08c",
X"08ffb405",
X"0c83c08c",
X"08c40508",
X"83c08c08",
X"ffb40508",
X"34880b83",
X"c08c08ff",
X"b4050881",
X"0534800b",
X"83c08c08",
X"ffb40508",
X"82053483",
X"c08c08ff",
X"b4050808",
X"ffa1ff06",
X"a0800783",
X"c08c08ff",
X"b405080c",
X"83c08c08",
X"c4050881",
X"057081ff",
X"0683c08c",
X"08c4050c",
X"83c08c08",
X"ffb4050c",
X"810b83c0",
X"8c08c405",
X"0827fedb",
X"3883c08c",
X"08ec0570",
X"5483c08c",
X"08c8050c",
X"925283c0",
X"8c08d405",
X"085180cd",
X"993f83c0",
X"800881ff",
X"067083c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"05088dea",
X"3883c08c",
X"08f40551",
X"f18c3f83",
X"c0800883",
X"ffff0683",
X"c08c08f6",
X"055283c0",
X"8c08e405",
X"0cf0f33f",
X"83c08008",
X"83ffff06",
X"83c08c08",
X"fd053383",
X"c08c08ff",
X"b8050883",
X"c08c08c4",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08c40508",
X"83c08c08",
X"ffbc0508",
X"2780fe38",
X"83c08c08",
X"c8050854",
X"83c08c08",
X"c4050853",
X"895283c0",
X"8c08d405",
X"085180cc",
X"9e3f83c0",
X"800881ff",
X"0683c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"0880f238",
X"83c08c08",
X"ee0551ef",
X"f13f83c0",
X"800883ff",
X"ff065383",
X"c08c08c4",
X"05085283",
X"c08c08d4",
X"050851f0",
X"b33f83c0",
X"8c08c405",
X"08810570",
X"81ff0683",
X"c08c08c4",
X"050c83c0",
X"8c08ffb4",
X"050cfef1",
X"3983c08c",
X"08c00508",
X"81053383",
X"c08c08ff",
X"b4050c81",
X"db0b83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb4",
X"0508802e",
X"8be03894",
X"3983c08c",
X"08ffb805",
X"0883c08c",
X"08ffbc05",
X"0c8bcb39",
X"83c08c08",
X"f1053352",
X"83c08c08",
X"d4050851",
X"80cb9c3f",
X"800b83c0",
X"8c08c005",
X"08810533",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"c4050c83",
X"c08c08c4",
X"050883c0",
X"8c08ffb4",
X"05082789",
X"e63883c0",
X"8c08c405",
X"0880d829",
X"7083c08c",
X"08c00508",
X"05708805",
X"70830533",
X"83c08c08",
X"cc050c83",
X"c08c08c8",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08d805",
X"0c83c08c",
X"08cc0508",
X"87a63883",
X"c08c08c8",
X"05082202",
X"84057186",
X"0587fffc",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08dc050c",
X"83c08c08",
X"ffb8050c",
X"0283c08c",
X"08ffb405",
X"08310d89",
X"3d705983",
X"c08c08ff",
X"b8050858",
X"83c08c08",
X"ffbc0508",
X"87053357",
X"83c08c08",
X"ffb4050c",
X"a25583c0",
X"8c08cc05",
X"08548653",
X"81815283",
X"c08c08d4",
X"050851be",
X"933f83c0",
X"800881ff",
X"0683c08c",
X"08d0050c",
X"83c08c08",
X"d0050881",
X"c13883c0",
X"8c08ffbc",
X"05089605",
X"5383c08c",
X"08ffb805",
X"085283c0",
X"8c08ffb4",
X"050851a1",
X"c63f83c0",
X"800881ff",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb405",
X"08802e81",
X"853883c0",
X"8c08ffbc",
X"05089405",
X"83c08c08",
X"ffbc0508",
X"96053370",
X"862a83c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08cc05",
X"0c83c08c",
X"08ffb405",
X"08832e09",
X"810680c6",
X"3883c08c",
X"08ffb405",
X"0883c08c",
X"08c80508",
X"82053483",
X"cae83370",
X"810583c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb4",
X"050883ca",
X"e83483c0",
X"8c08ffb8",
X"050883c0",
X"8c08cc05",
X"083483c0",
X"8c08dc05",
X"080d83c0",
X"8c08d005",
X"0881ff06",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"fbff3883",
X"c08c08d8",
X"050883c0",
X"8c08c005",
X"08058805",
X"70820533",
X"5183c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb405",
X"08832e09",
X"810680e3",
X"3883c08c",
X"08ffb805",
X"0883c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb405",
X"08810570",
X"81ff0651",
X"83c08c08",
X"ffb4050c",
X"810b83c0",
X"8c08ffb4",
X"050827dd",
X"38800b83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b4050881",
X"057081ff",
X"065183c0",
X"8c08ffb4",
X"050c970b",
X"83c08c08",
X"ffb40508",
X"27dd3883",
X"c08c08e4",
X"050880f9",
X"32703070",
X"80255151",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"e0050891",
X"2e098106",
X"80f93883",
X"c08c08ff",
X"b4050880",
X"2e80ec38",
X"83c08c08",
X"c4050880",
X"e238850b",
X"83c08c08",
X"c00508a6",
X"0534a00b",
X"83c08c08",
X"c00508a7",
X"0534850b",
X"83c08c08",
X"c00508a8",
X"053480c0",
X"0b83c08c",
X"08c00508",
X"a9053486",
X"0b83c08c",
X"08c00508",
X"aa053490",
X"0b83c08c",
X"08c00508",
X"ab053486",
X"0b83c08c",
X"08c00508",
X"ac0534a0",
X"0b83c08c",
X"08c00508",
X"ad053483",
X"c08c08e4",
X"050889d8",
X"32703070",
X"80255151",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"e0050883",
X"edec2e09",
X"810680f6",
X"38817083",
X"c08c08ff",
X"b4050806",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb40508",
X"802e80ce",
X"3883c08c",
X"08c40508",
X"80c43884",
X"0b83c08c",
X"08c00508",
X"aa053480",
X"c00b83c0",
X"8c08c005",
X"08ab0534",
X"840b83c0",
X"8c08c005",
X"08ac0534",
X"900b83c0",
X"8c08c005",
X"08ad0534",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"c005088c",
X"053483c0",
X"8c08e405",
X"0880f932",
X"70307080",
X"25515183",
X"c08c08ff",
X"b4050c83",
X"c08c08e0",
X"0508862e",
X"09810680",
X"c3388170",
X"83c08c08",
X"ffb40508",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb405",
X"08802e9c",
X"3883c08c",
X"08c40508",
X"933883c0",
X"8c08ffb8",
X"050883c0",
X"8c08c005",
X"088d0534",
X"83c08c08",
X"c4050880",
X"d82983c0",
X"8c08c005",
X"08057084",
X"05708305",
X"3383c08c",
X"08ffb405",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"ffbc050c",
X"80588057",
X"83c08c08",
X"ffb40508",
X"56805580",
X"548a53a1",
X"5283c08c",
X"08d40508",
X"51b78d3f",
X"83c08008",
X"81ff0670",
X"30709f2a",
X"5183c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"08a02e8c",
X"3883c08c",
X"08ffb405",
X"08f6c238",
X"83c08c08",
X"ffbc0508",
X"8b053383",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b4050880",
X"2eb33883",
X"c08c08c8",
X"05088305",
X"3383c08c",
X"08ffb405",
X"0c805880",
X"5783c08c",
X"08ffb405",
X"08568055",
X"80548b53",
X"a15283c0",
X"8c08d405",
X"0851b688",
X"3f83c08c",
X"08c40508",
X"81057081",
X"ff0683c0",
X"8c08c005",
X"08810533",
X"5283c08c",
X"08c4050c",
X"83c08c08",
X"ffb4050c",
X"f6893980",
X"0b83c08c",
X"08c4050c",
X"83c08c08",
X"c4050880",
X"d82983c0",
X"8c08d405",
X"0805709a",
X"053383c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb4",
X"0508822e",
X"098106a9",
X"3883cb84",
X"56815580",
X"5483c08c",
X"08ffb405",
X"085383c0",
X"8c08ffb8",
X"05089705",
X"335283c0",
X"8c08d405",
X"0851e48a",
X"3f83c08c",
X"08c40508",
X"81057081",
X"ff0683c0",
X"8c08c405",
X"0c83c08c",
X"08ffb405",
X"0c810b83",
X"c08c08c4",
X"050827fe",
X"fb38810b",
X"83c08c08",
X"c0050834",
X"800b83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08e805",
X"080d83c0",
X"8c08ffbc",
X"050883c0",
X"800c9c3d",
X"0d83c08c",
X"0c04f53d",
X"0d901e57",
X"800b8118",
X"33545978",
X"7327819d",
X"387880d8",
X"29178a11",
X"33545472",
X"832e0981",
X"0680f838",
X"9414335b",
X"a98c3f83",
X"c080085a",
X"80567581",
X"c4291a87",
X"11335454",
X"72802e80",
X"c0387308",
X"81d5982e",
X"098106b5",
X"38807459",
X"557480d8",
X"29189a11",
X"33545472",
X"832e0981",
X"069238a4",
X"14703354",
X"547a7327",
X"8738ff13",
X"53727434",
X"81157081",
X"ff065653",
X"817527d1",
X"38811670",
X"81ff0657",
X"538f7627",
X"ffa43883",
X"cae833ff",
X"05537283",
X"cae83481",
X"197081ff",
X"06811933",
X"5e5a537b",
X"7926fee5",
X"38800b83",
X"c0800c8d",
X"3d0d0483",
X"c08c0802",
X"83c08c0c",
X"e63d0d83",
X"c08c0888",
X"05080284",
X"05719005",
X"70337083",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08c8",
X"050c83c0",
X"8c08dc05",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"ffa40508",
X"802e94b5",
X"38800b83",
X"c08c08c8",
X"05088105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08d4050c",
X"83c08c08",
X"d4050883",
X"c08c08ff",
X"a4050825",
X"93fd3883",
X"c08c08d4",
X"050880d8",
X"2983c08c",
X"08c80508",
X"05840570",
X"86053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"a4050880",
X"2e938938",
X"a6b23f83",
X"c08c08ff",
X"b8050880",
X"d4050883",
X"c0800826",
X"92f23802",
X"83c08c08",
X"ffb80508",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08d8",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08fc05",
X"2383c08c",
X"08ffa405",
X"08860583",
X"fc0683c0",
X"8c08ffa4",
X"050c0283",
X"c08c08ff",
X"a4050831",
X"0d853d70",
X"5583c08c",
X"08fc0554",
X"83c08c08",
X"ffb80508",
X"5383c08c",
X"08e00508",
X"5283c08c",
X"08c0050c",
X"ae8a3f83",
X"c0800881",
X"ff0683c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"050891bb",
X"3883c08c",
X"08ffb805",
X"08870533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e80d5",
X"3883c08c",
X"08ffb805",
X"08860533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"822e0981",
X"06b33883",
X"c08c08fc",
X"052283c0",
X"8c08ffa4",
X"050c870b",
X"83c08c08",
X"ffa40508",
X"27973883",
X"c08c08c0",
X"05088205",
X"5283c08c",
X"08c00508",
X"3351dba6",
X"3f83c08c",
X"08ffb805",
X"08860533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"832e0981",
X"0690a438",
X"83c08c08",
X"ffb80508",
X"92057082",
X"053383c0",
X"8c08fc05",
X"2283c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08c4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffa80508",
X"268fe438",
X"800b83c0",
X"8c08e405",
X"0c800b83",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"b0050810",
X"83c08c08",
X"05f80583",
X"c08c08ff",
X"b0050884",
X"2983c08c",
X"08ffb005",
X"08100583",
X"c08c08c4",
X"05080570",
X"84057033",
X"83c08c08",
X"c0050805",
X"703383c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffbc",
X"05082383",
X"c08c08ff",
X"a8050881",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508902e",
X"098106be",
X"3883c08c",
X"08ffa805",
X"083383c0",
X"8c08c005",
X"08058105",
X"70337082",
X"802983c0",
X"8c08ffb4",
X"05080551",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffbc05",
X"082383c0",
X"8c08ffac",
X"05088605",
X"2283c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa805",
X"08a23883",
X"c08c08ff",
X"ac050888",
X"052283c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"050881ff",
X"2e80e538",
X"83c08c08",
X"ffbc0508",
X"227083c0",
X"8c08ffa8",
X"05083170",
X"82802971",
X"3183c08c",
X"08ffac05",
X"08880522",
X"7083c08c",
X"08ffa805",
X"08317073",
X"355383c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c5183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"bc050823",
X"83c08c08",
X"ffb00508",
X"81057081",
X"ff0683c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa4",
X"050c810b",
X"83c08c08",
X"ffb00508",
X"27fce038",
X"83c08c08",
X"f8052283",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a40508bf",
X"26913883",
X"c08c08e4",
X"05088207",
X"83c08c08",
X"e4050c81",
X"c00b83c0",
X"8c08ffa4",
X"05082791",
X"3883c08c",
X"08e40508",
X"810783c0",
X"8c08e405",
X"0c83c08c",
X"08fa0522",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"bf269138",
X"83c08c08",
X"e4050888",
X"0783c08c",
X"08e4050c",
X"81c00b83",
X"c08c08ff",
X"a4050827",
X"913883c0",
X"8c08e405",
X"08840783",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffb00508",
X"1083c08c",
X"08c40508",
X"05709005",
X"703383c0",
X"8c08c005",
X"08057033",
X"72810533",
X"70720651",
X"535183c0",
X"8c08ffa8",
X"050c5183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e9b3890",
X"0b83c08c",
X"08ffb005",
X"082b83c0",
X"8c08e405",
X"080783c0",
X"8c08e405",
X"0c83c08c",
X"08ffb005",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a4050c97",
X"0b83c08c",
X"08ffb005",
X"0827fef4",
X"3883c08c",
X"08ffb805",
X"08900533",
X"83c08c08",
X"e4050883",
X"c08c08ff",
X"b4050c83",
X"c08c08c4",
X"050c83c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffb8",
X"05088c05",
X"082e83ff",
X"3883c08c",
X"08ffb405",
X"0883c08c",
X"08ffb805",
X"088c050c",
X"83c08c08",
X"ffb80508",
X"89053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e83b938",
X"83c08c08",
X"e40583c0",
X"8c08ffb4",
X"05088f06",
X"83c08c08",
X"e4050c83",
X"c08c08cc",
X"050c800b",
X"83c08c08",
X"f0050c80",
X"0b83c08c",
X"08f40523",
X"800b81d7",
X"943383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffbc",
X"05082e82",
X"d33883c0",
X"8c08f005",
X"81d7940b",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"d0050c83",
X"c08c08ff",
X"ac050833",
X"83c08c08",
X"ffac0508",
X"81053381",
X"722b8172",
X"2b077083",
X"c08c08ff",
X"b4050806",
X"5283c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffa805",
X"082e0981",
X"0681be38",
X"83c08c08",
X"ffbc0508",
X"852680f6",
X"3883c08c",
X"08ffac05",
X"08820533",
X"7081ff06",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa40508",
X"802e80ca",
X"3883c08c",
X"08ffbc05",
X"0883c08c",
X"08ffbc05",
X"08810570",
X"81ff0683",
X"c08c08d0",
X"05087305",
X"5383c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb005",
X"0883c08c",
X"08ffa405",
X"083483c0",
X"8c08ffac",
X"05088305",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e9d",
X"38810b83",
X"c08c08ff",
X"a405082b",
X"83c08c08",
X"cc050808",
X"0783c08c",
X"08cc0508",
X"0c83c08c",
X"08ffac05",
X"08840570",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa405",
X"08fdc838",
X"83c08c08",
X"f0055280",
X"51d0c33f",
X"83c08c08",
X"e4050852",
X"83c08c08",
X"c4050851",
X"d1fe3f83",
X"c08c08fb",
X"05337081",
X"800a2981",
X"0a057098",
X"2c5583c0",
X"8c08ffa4",
X"050c83c0",
X"8c08f905",
X"33708180",
X"0a29810a",
X"0570982c",
X"5583c08c",
X"08ffa405",
X"0c83c08c",
X"08c40508",
X"5383c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa805",
X"0cd1d43f",
X"83c08c08",
X"ffb80508",
X"88053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e84e038",
X"83c08c08",
X"ffb80508",
X"90053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050881",
X"2684c038",
X"807081d7",
X"c80b81d7",
X"c80b8105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffb405",
X"082e81ae",
X"3883c08c",
X"08ffac05",
X"08842983",
X"c08c08ff",
X"a8050805",
X"703383c0",
X"8c08c005",
X"08057033",
X"72810533",
X"70720651",
X"535183c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"aa38810b",
X"83c08c08",
X"ffac0508",
X"2b83c08c",
X"08ffb405",
X"08077083",
X"ffff0683",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"ac050881",
X"057081ff",
X"0681d7c8",
X"71842971",
X"05708105",
X"33515383",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a40508fe",
X"d43883c0",
X"8c08ffb8",
X"05088a05",
X"2283c08c",
X"08c0050c",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"c005082e",
X"82ad3880",
X"0b83c08c",
X"08e8050c",
X"800b83c0",
X"8c08ec05",
X"23807083",
X"c08c08e8",
X"0583c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffb005",
X"0c81af39",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffac0508",
X"2c708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e80",
X"e73883c0",
X"8c08ffb0",
X"050883c0",
X"8c08ffb0",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ffbc0508",
X"730583c0",
X"8c08ffb8",
X"05089005",
X"3383c08c",
X"08ffac05",
X"08842905",
X"535383c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050881d7",
X"ca053383",
X"c08c08ff",
X"a4050834",
X"83c08c08",
X"ffac0508",
X"81057081",
X"ff0683c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa4",
X"050c8f0b",
X"83c08c08",
X"ffac0508",
X"2783c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb005",
X"0885268c",
X"3883c08c",
X"08ffa405",
X"08fea938",
X"83c08c08",
X"e8055280",
X"51caf33f",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffb80508",
X"8a052383",
X"c08c08ff",
X"b8050880",
X"d2053383",
X"c08c08ff",
X"b8050880",
X"d4050805",
X"83c08c08",
X"ffb80508",
X"80d4050c",
X"83c08c08",
X"d805080d",
X"83c08c08",
X"d4050881",
X"800a2981",
X"800a0570",
X"982c83c0",
X"8c08c805",
X"08810533",
X"83c08c08",
X"ffa8050c",
X"5183c08c",
X"08d4050c",
X"83c08c08",
X"ffa80508",
X"83c08c08",
X"d4050824",
X"ec853880",
X"0b83c08c",
X"08ffa805",
X"0c83c08c",
X"08dc0508",
X"0d83c08c",
X"08ffa805",
X"0883c080",
X"0c9c3d0d",
X"83c08c0c",
X"04f33d0d",
X"02bf0533",
X"02840580",
X"c3053383",
X"cb84335a",
X"5b597980",
X"2e8d3878",
X"78065776",
X"802e8e38",
X"81893978",
X"78065776",
X"802e80ff",
X"3883cb84",
X"33707a07",
X"58587988",
X"38780970",
X"79065157",
X"7683cb84",
X"3492973f",
X"83c08008",
X"5e805c8f",
X"5d7d1c87",
X"11335858",
X"76802e80",
X"c1387708",
X"81d5982e",
X"098106b6",
X"38805b81",
X"5a7d1c70",
X"1c9a1133",
X"59595976",
X"822e0981",
X"06943883",
X"cb845681",
X"55805476",
X"53971833",
X"527851cb",
X"c53fff1a",
X"80d81c5c",
X"5a798025",
X"d038ff1d",
X"81c41d5d",
X"5d7c8025",
X"ffa7388f",
X"3d0d04e9",
X"3d0d696c",
X"02880580",
X"ea05225c",
X"5a5b8070",
X"71415e58",
X"ff78797a",
X"7b7c7d46",
X"4c4a4540",
X"5d436299",
X"3d346202",
X"840580dd",
X"05347779",
X"2280ffff",
X"06544572",
X"79237978",
X"2e888738",
X"7a708105",
X"5c337084",
X"2a718c06",
X"70822a5a",
X"56568306",
X"ff1b7083",
X"ffff065c",
X"54568054",
X"75742e91",
X"387a7081",
X"055c33ff",
X"1b7083ff",
X"ff065c54",
X"54817627",
X"9b387381",
X"ff067b70",
X"81055d33",
X"55748280",
X"2905ff1b",
X"7083ffff",
X"065c5454",
X"827627aa",
X"387383ff",
X"ff067b70",
X"81055d33",
X"70902b72",
X"077d7081",
X"055f3370",
X"982b7207",
X"fe1f7083",
X"ffff0640",
X"52525252",
X"54547e80",
X"2e80c438",
X"7686f738",
X"748a2e09",
X"81069438",
X"811f7081",
X"ff06811e",
X"7081ff06",
X"5f524053",
X"86dc3974",
X"8c2e0981",
X"0686d338",
X"ff1f7081",
X"ff06ff1e",
X"7081ff06",
X"5f524053",
X"7b632586",
X"bd38ff43",
X"86b83976",
X"812e83bb",
X"38768124",
X"89387680",
X"2e8d3886",
X"a5397682",
X"2e84a638",
X"869c39f8",
X"15537284",
X"26849538",
X"72842981",
X"d8880553",
X"72080464",
X"802e80cd",
X"38782283",
X"80800653",
X"72838080",
X"2e098106",
X"bc388056",
X"756427a4",
X"38751e70",
X"83ffff06",
X"77101b90",
X"1172832a",
X"58515751",
X"53737534",
X"72870681",
X"712b5153",
X"72811634",
X"81167081",
X"ff065753",
X"977627cc",
X"387f8407",
X"40800b99",
X"3d435661",
X"16703370",
X"982b7098",
X"2c515151",
X"53807324",
X"80fb3860",
X"73291e70",
X"83ffff06",
X"7a228380",
X"80065258",
X"53728380",
X"802e0981",
X"0680de38",
X"60883270",
X"30707207",
X"80256390",
X"32703070",
X"72078025",
X"73075354",
X"58515553",
X"73802ebd",
X"38768706",
X"5372b638",
X"75842976",
X"10057911",
X"84117983",
X"2a575751",
X"53737534",
X"60811634",
X"65861423",
X"66881423",
X"7587387f",
X"8107408d",
X"3975812e",
X"09810685",
X"387f8207",
X"40811670",
X"81ff0657",
X"53817627",
X"fee53863",
X"61291e70",
X"83ffff06",
X"5f538070",
X"4642ff02",
X"840580dd",
X"0534ff0b",
X"993d3483",
X"f539811c",
X"7081ff06",
X"5d538042",
X"73812e09",
X"81068e38",
X"7781800a",
X"2981800a",
X"055880d3",
X"3973802e",
X"89387382",
X"2e098106",
X"8d387c81",
X"800a2981",
X"800a055d",
X"a439815f",
X"83b839ff",
X"1c7081ff",
X"065d537b",
X"63258338",
X"ff437c80",
X"2e92387c",
X"81800a29",
X"81ff0a05",
X"5d7c982c",
X"5d839339",
X"77802e92",
X"38778180",
X"0a2981ff",
X"0a055877",
X"982c5882",
X"fd397753",
X"839e3974",
X"892680f4",
X"38748429",
X"81d89c05",
X"53720804",
X"73872e82",
X"e1387385",
X"2e82db38",
X"73882e82",
X"d538738c",
X"2e82cf38",
X"73892e09",
X"81068638",
X"814582c2",
X"3973812e",
X"09810682",
X"b9386280",
X"2582b338",
X"7b982b70",
X"982c5143",
X"82a83973",
X"83ffff06",
X"46829f39",
X"7383ffff",
X"06478296",
X"397381ff",
X"0641828e",
X"3973811a",
X"34828739",
X"7381ff06",
X"4481ff39",
X"7e5382a0",
X"3974812e",
X"81e33874",
X"81248938",
X"74802e8d",
X"3881e739",
X"74822e81",
X"d83881de",
X"3974567b",
X"83388156",
X"74537386",
X"2e098106",
X"97387581",
X"06537280",
X"2e8e3878",
X"2282ffff",
X"06fe8080",
X"0753b639",
X"7b833881",
X"5373822e",
X"09810697",
X"38728106",
X"5372802e",
X"8e387822",
X"81ffff06",
X"81808007",
X"5393397b",
X"9638fc14",
X"53728126",
X"8e387822",
X"ff808007",
X"53727923",
X"80e53980",
X"5573812e",
X"09810683",
X"38735577",
X"5377802e",
X"89387481",
X"06537280",
X"ca3872d0",
X"15545572",
X"81268338",
X"81557780",
X"2eb93874",
X"81065372",
X"802eb038",
X"78228380",
X"80065372",
X"8380802e",
X"0981069f",
X"3873b02e",
X"09810687",
X"3861993d",
X"34913973",
X"b12e0981",
X"06893861",
X"02840580",
X"dd053461",
X"8105538c",
X"39617431",
X"81055384",
X"39611453",
X"7283ffff",
X"064279f7",
X"fb387d83",
X"2a537282",
X"1a347822",
X"83808006",
X"53728380",
X"802e0981",
X"06883881",
X"537f872e",
X"83388053",
X"7283c080",
X"0c993d0d",
X"04fd3d0d",
X"75831133",
X"82123371",
X"982b7190",
X"2b078114",
X"3370882b",
X"72077533",
X"710783c0",
X"800c5253",
X"54565452",
X"853d0d04",
X"f63d0d02",
X"b7053302",
X"8405bb05",
X"33028805",
X"bf05335b",
X"5b5b8058",
X"80577888",
X"2b7a0756",
X"80557a54",
X"8153a352",
X"7c5192cc",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8c3d0d04",
X"f63d0d02",
X"b7053302",
X"8405bb05",
X"33028805",
X"bf05335b",
X"5b5b8058",
X"80577888",
X"2b7a0756",
X"80557a54",
X"8353a352",
X"7c519290",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8c3d0d04",
X"f73d0d02",
X"b3053302",
X"8405b605",
X"22605a58",
X"56805580",
X"54805381",
X"a3527b51",
X"91e23f83",
X"c0800881",
X"ff0683c0",
X"800c8b3d",
X"0d04ee3d",
X"0d649011",
X"5c5c807b",
X"34800b84",
X"1c0c800b",
X"881c3481",
X"0b891c34",
X"880b8a1c",
X"34800b8b",
X"1c34881b",
X"08c10681",
X"07881c0c",
X"8f3d7054",
X"5d88527b",
X"519beb3f",
X"83c08008",
X"81ff0670",
X"5b597881",
X"a938903d",
X"335e81db",
X"5a7d892e",
X"09810681",
X"99387c53",
X"92527b51",
X"9bc43f83",
X"c0800881",
X"ff06705b",
X"59788182",
X"387c5888",
X"577856a9",
X"55785486",
X"5381a052",
X"7b5190d0",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"80e03802",
X"ba05337b",
X"347c5478",
X"537d527b",
X"519bac3f",
X"83c08008",
X"81ff0670",
X"5b597880",
X"c13802bd",
X"0533527b",
X"519bc43f",
X"83c08008",
X"81ff0670",
X"5b5978aa",
X"38817b33",
X"5a5a7979",
X"26993880",
X"54795388",
X"527b51fd",
X"bb3f811a",
X"7081ff06",
X"7c33525b",
X"59e43981",
X"0b881c34",
X"805a7983",
X"c0800c94",
X"3d0d0480",
X"0b83c080",
X"0c04f93d",
X"0d790284",
X"05ab0533",
X"8e3d7054",
X"585858ff",
X"beb03f8a",
X"3d8a0551",
X"ffbea73f",
X"7551fc8d",
X"3f83c080",
X"08848681",
X"2ebe3883",
X"c0800884",
X"86812699",
X"3883c080",
X"08848280",
X"2e80e638",
X"83c08008",
X"8482812e",
X"9f3881b4",
X"3983c080",
X"0880c082",
X"832e80f4",
X"3883c080",
X"0880c086",
X"832e80e8",
X"38819939",
X"83c09c33",
X"55805674",
X"762e0981",
X"06818b38",
X"74547653",
X"91527751",
X"fbd63f74",
X"54765390",
X"527751fb",
X"cb3f7454",
X"76538452",
X"7751fbfc",
X"3f810b83",
X"c09c3481",
X"b15680de",
X"39805476",
X"53915277",
X"51fba93f",
X"80547653",
X"90527751",
X"fb9e3f80",
X"0b83c09c",
X"34765287",
X"18335197",
X"963fb539",
X"80547653",
X"94527751",
X"fb823f80",
X"54765390",
X"527751fa",
X"f73f7551",
X"ffbcdb3f",
X"83c08008",
X"892a8106",
X"53765287",
X"18335190",
X"cd3f800b",
X"83c09c34",
X"80567583",
X"c0800c89",
X"3d0d04f2",
X"3d0d6090",
X"115a5880",
X"0b881a33",
X"71595656",
X"74762e82",
X"a53882ac",
X"3f841908",
X"83c08008",
X"26829538",
X"78335a81",
X"0b8e3d23",
X"903df811",
X"55f40553",
X"99185277",
X"518ae53f",
X"83c08008",
X"81ff0670",
X"57557477",
X"2e098106",
X"81d93886",
X"39745681",
X"d2398156",
X"82578e3d",
X"33770655",
X"74802ebb",
X"38800b8d",
X"3d34903d",
X"f0055484",
X"53755277",
X"51facd3f",
X"83c08008",
X"81ff0655",
X"749d387b",
X"53755277",
X"51fce73f",
X"83c08008",
X"81ff0655",
X"7481b12e",
X"818b3874",
X"ffb33876",
X"1081fc06",
X"81177081",
X"ff065856",
X"57877627",
X"ffa83881",
X"56757a26",
X"80eb3880",
X"0b8d3d34",
X"8c3d7055",
X"57845375",
X"527751f9",
X"f73f83c0",
X"800881ff",
X"06557480",
X"c1387651",
X"ffbad73f",
X"83c08008",
X"82870655",
X"7482812e",
X"098106aa",
X"3802ae05",
X"33810755",
X"74028405",
X"ae05347b",
X"53755277",
X"51fbeb3f",
X"83c08008",
X"81ff0655",
X"7481b12e",
X"903874fe",
X"b8388116",
X"7081ff06",
X"5755ff91",
X"39805675",
X"81ff0656",
X"973f83c0",
X"80088fd0",
X"05841a0c",
X"75577683",
X"c0800c90",
X"3d0d0404",
X"9080a008",
X"83c0800c",
X"04ff3d0d",
X"7387e829",
X"51ff91b9",
X"3f833d0d",
X"040483cb",
X"880b83c0",
X"800c04fd",
X"3d0d7577",
X"5454800b",
X"83cae834",
X"728a3890",
X"90800b84",
X"150c9039",
X"72812e09",
X"81068838",
X"9098800b",
X"84150c84",
X"140883cb",
X"800c800b",
X"88150c80",
X"0b8c150c",
X"83cb8008",
X"53820b87",
X"80143481",
X"51ff9e3f",
X"83cb8008",
X"53800b88",
X"143483cb",
X"80085381",
X"0b878014",
X"3483cb80",
X"0853800b",
X"8c143483",
X"cb800853",
X"800ba414",
X"34917434",
X"800b83c0",
X"a034800b",
X"83c0a434",
X"800b83c0",
X"a8348054",
X"7381c429",
X"83cb8c05",
X"53800b83",
X"14348114",
X"7081ff06",
X"55538f74",
X"27e63885",
X"3d0d04fe",
X"3d0d7476",
X"82113370",
X"bf068171",
X"2bff0556",
X"51515253",
X"90712783",
X"38ff5276",
X"51717123",
X"83cb8008",
X"51871333",
X"90123480",
X"0b83c0a4",
X"34800b83",
X"c0a83488",
X"13338a14",
X"33525271",
X"802eaa38",
X"7081ff06",
X"51845270",
X"83387052",
X"7183c0a4",
X"348a1333",
X"70307080",
X"25842b70",
X"88075151",
X"52537083",
X"c0a83490",
X"397081ff",
X"06517083",
X"38985271",
X"83c0a834",
X"800b83c0",
X"800c843d",
X"0d04f13d",
X"0d616568",
X"028c0580",
X"cb053302",
X"900580ce",
X"05220294",
X"0580d605",
X"22424041",
X"5a4040fd",
X"8b3f83c0",
X"8008a788",
X"055b8070",
X"715b5b52",
X"83943983",
X"cb800851",
X"7d941234",
X"83c0a433",
X"81075580",
X"7054567f",
X"862680ea",
X"387f8429",
X"81d8d005",
X"83cb8008",
X"53517008",
X"04800b84",
X"1334a139",
X"77337030",
X"70802583",
X"71315151",
X"52537084",
X"13348d39",
X"810b8413",
X"34b83983",
X"0b841334",
X"81705456",
X"ad39810b",
X"841334a2",
X"39773370",
X"30708025",
X"83713151",
X"51525370",
X"84133480",
X"78335252",
X"70833881",
X"52717834",
X"81537488",
X"075583c0",
X"a83383cb",
X"80085257",
X"810b81d0",
X"123483cb",
X"80085181",
X"0b819012",
X"347e802e",
X"ae387280",
X"2ea9387e",
X"ff1e5254",
X"7083ffff",
X"06537283",
X"ffff2e97",
X"38737081",
X"05553383",
X"cb800853",
X"517081c0",
X"1334ff13",
X"51de3983",
X"cb8008a8",
X"11335351",
X"76881234",
X"83cb8008",
X"51747134",
X"81ff5291",
X"3983cb80",
X"08a01133",
X"70810651",
X"5253708f",
X"38fafd3f",
X"7a83c080",
X"0826e638",
X"81883981",
X"0ba01434",
X"83cb8008",
X"a8113380",
X"ff067078",
X"07525351",
X"70802e80",
X"ed387186",
X"2a708106",
X"51517080",
X"2e913880",
X"78335253",
X"70833881",
X"53727834",
X"80e03971",
X"842a7081",
X"06515170",
X"802e9b38",
X"81197083",
X"ffff067d",
X"30709f2a",
X"51525a51",
X"787c2e09",
X"8106af38",
X"a4397183",
X"2a708106",
X"51517080",
X"2e933881",
X"1a7081ff",
X"065b5179",
X"832e0981",
X"0690388a",
X"3971a306",
X"5170802e",
X"85387151",
X"9239f9e4",
X"3f7a83c0",
X"800826fc",
X"e2387181",
X"bf065170",
X"83c0800c",
X"913d0d04",
X"f63d0d02",
X"b3053302",
X"8405b705",
X"33028805",
X"ba052259",
X"5959800b",
X"8c3d348c",
X"3dfc0556",
X"80558054",
X"76537752",
X"7851fbf2",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8c3d0d04",
X"f33d0d7f",
X"6264028c",
X"0580c205",
X"22722281",
X"1533425f",
X"415e5959",
X"8078237d",
X"53783352",
X"8151ffa0",
X"3f83c080",
X"0881ff06",
X"5675802e",
X"86387554",
X"81ad3983",
X"cb8008a8",
X"1133821b",
X"3370862a",
X"70810673",
X"982b5351",
X"575c5657",
X"79802583",
X"38815673",
X"762e8738",
X"81f05481",
X"8239818c",
X"17337081",
X"ff067922",
X"7d713190",
X"2b70902c",
X"7009709f",
X"2c720670",
X"52525351",
X"53575754",
X"75742483",
X"38755574",
X"84808029",
X"fc808005",
X"70902c51",
X"5574ff2e",
X"943883cb",
X"80088180",
X"11335154",
X"737c7081",
X"055e34db",
X"39772276",
X"05547378",
X"23790970",
X"9f2a7081",
X"06821c33",
X"81bf0671",
X"862b0751",
X"51515473",
X"821a347c",
X"76268a38",
X"7722547a",
X"7426febb",
X"38805473",
X"83c0800c",
X"8f3d0d04",
X"f93d0d7a",
X"57800b89",
X"3d23893d",
X"fc055376",
X"527951f8",
X"da3f83c0",
X"800881ff",
X"06705755",
X"7496387c",
X"547b5388",
X"3d225276",
X"51fde53f",
X"83c08008",
X"81ff0656",
X"7583c080",
X"0c893d0d",
X"04f03d0d",
X"62660288",
X"0580ce05",
X"22415d5e",
X"80028405",
X"80d20522",
X"7f810533",
X"ff115a5d",
X"5a5d81da",
X"5876bf26",
X"80e93878",
X"802e80e1",
X"387a5878",
X"7b278338",
X"7858821e",
X"3370872a",
X"585a7692",
X"3d34923d",
X"fc055677",
X"557b547e",
X"537d3352",
X"8251f8de",
X"3f83c080",
X"0881ff06",
X"5d800b92",
X"3d33585a",
X"76802e83",
X"38815a82",
X"1e3380ff",
X"067a872b",
X"07577682",
X"1f347c91",
X"38787831",
X"7083ffff",
X"06791e5e",
X"5a57ff9b",
X"397c5877",
X"83c0800c",
X"923d0d04",
X"f83d0d7b",
X"028405b2",
X"05225858",
X"800b8a3d",
X"238a3dfc",
X"05537752",
X"7a51f6f7",
X"3f83c080",
X"0881ff06",
X"70575574",
X"96387d54",
X"7653893d",
X"22527751",
X"feaf3f83",
X"c0800881",
X"ff065675",
X"83c0800c",
X"8a3d0d04",
X"ec3d0d66",
X"6e028805",
X"80df0533",
X"028c0580",
X"e3053302",
X"900580e7",
X"05330294",
X"0580eb05",
X"33029805",
X"80ee0522",
X"4143415f",
X"5c405702",
X"80f20522",
X"963d2396",
X"3df00553",
X"84177053",
X"775259f6",
X"863f83c0",
X"800881ff",
X"06587781",
X"e538777a",
X"81800658",
X"40807725",
X"83388140",
X"79943d34",
X"7b028405",
X"80c90534",
X"7c028405",
X"80ca0534",
X"7d028405",
X"80cb0534",
X"7a953d34",
X"7a882a57",
X"76028405",
X"80cd0534",
X"953d2257",
X"76028405",
X"80ce0534",
X"76882a57",
X"76028405",
X"80cf0534",
X"77923d34",
X"963dec11",
X"57578855",
X"f4175492",
X"3d225377",
X"527751f6",
X"953f83c0",
X"800881ff",
X"06587780",
X"ed387e80",
X"2e80cb38",
X"923d2279",
X"0858587f",
X"802e9c38",
X"76818080",
X"07790c7e",
X"54963dfc",
X"05537783",
X"ffff0652",
X"7851f9fc",
X"3f993976",
X"82808007",
X"790c7e54",
X"953d2253",
X"7783ffff",
X"06527851",
X"fc8f3f83",
X"c0800881",
X"ff065877",
X"9d38923d",
X"22538052",
X"7f307080",
X"25847131",
X"535157f9",
X"873f83c0",
X"800881ff",
X"06587783",
X"c0800c96",
X"3d0d04f6",
X"3d0d7c02",
X"8405b705",
X"335b5b80",
X"58805780",
X"56805579",
X"54855380",
X"527a51fd",
X"a33f83c0",
X"800881ff",
X"06597885",
X"3879871c",
X"347883c0",
X"800c8c3d",
X"0d04f93d",
X"0d02a705",
X"33028405",
X"ab053302",
X"8805af05",
X"33585957",
X"800b83cb",
X"8f335454",
X"72742e9f",
X"38811470",
X"81ff0655",
X"53738f26",
X"81b63873",
X"81c42983",
X"cb8c0583",
X"11335153",
X"72e33873",
X"81c42983",
X"cb880555",
X"800b8716",
X"34768816",
X"34758a16",
X"34778916",
X"3480750c",
X"83cb8008",
X"8c160c80",
X"0b841634",
X"880b8516",
X"34800b86",
X"16348415",
X"08ffa1ff",
X"06a08007",
X"84160c81",
X"147081ff",
X"06535374",
X"51febc3f",
X"83c08008",
X"81ff0670",
X"55537280",
X"cd388a39",
X"7308750c",
X"725480c2",
X"397281dd",
X"f0555681",
X"ddf00880",
X"2eb23875",
X"84291470",
X"08765370",
X"08515454",
X"722d83c0",
X"800881ff",
X"06537280",
X"2ece3881",
X"167081ff",
X"0681ddf0",
X"71842911",
X"53565753",
X"7208d038",
X"80547383",
X"c0800c89",
X"3d0d04f9",
X"3d0d7957",
X"800b8418",
X"0883cb80",
X"0c58f088",
X"3f881708",
X"83c08008",
X"2783ed38",
X"effa3f83",
X"c0800881",
X"0588180c",
X"83cb8008",
X"b8113370",
X"81ff0651",
X"51547381",
X"2ea43873",
X"81248838",
X"73782e8a",
X"38b83973",
X"822e9538",
X"b1397633",
X"81f00654",
X"73902ea6",
X"38917734",
X"a1397358",
X"763381f0",
X"06547390",
X"2e098106",
X"9138efa8",
X"3f83c080",
X"0881c805",
X"8c180ca0",
X"77348056",
X"7581c429",
X"83cb8f11",
X"33555573",
X"802eaa38",
X"83cb8815",
X"70085654",
X"74802e9d",
X"38881508",
X"802e9638",
X"8c140883",
X"cb80082e",
X"09810689",
X"38735188",
X"15085473",
X"2d811670",
X"81ff0657",
X"548f7627",
X"ffba3876",
X"335473b0",
X"2e819938",
X"73b0248f",
X"3873912e",
X"ab3873a0",
X"2e80f538",
X"82a63973",
X"80d02e81",
X"e4387380",
X"d0248b38",
X"7380c02e",
X"81993882",
X"8f397381",
X"802e81fb",
X"38828539",
X"80567581",
X"c42983cb",
X"8c118311",
X"33565955",
X"73802ea8",
X"3883cb88",
X"15700856",
X"5474802e",
X"9b388c14",
X"0883cb80",
X"082e0981",
X"068e3873",
X"51841508",
X"54732d80",
X"0b831934",
X"81167081",
X"ff065754",
X"8f7627ff",
X"b9389277",
X"3481b539",
X"edc23f8c",
X"170883c0",
X"80082781",
X"a738b077",
X"3481a139",
X"83cb8008",
X"54800b8c",
X"153483cb",
X"80085484",
X"0b881534",
X"80c07734",
X"ed963f83",
X"c08008b2",
X"058c180c",
X"80fa39ed",
X"873f8c17",
X"0883c080",
X"082780ec",
X"3883cb80",
X"0854810b",
X"8c153483",
X"cb800854",
X"800b8815",
X"3483cb80",
X"0854880b",
X"a01534ec",
X"db3f83c0",
X"80089405",
X"8c180c80",
X"d07734bc",
X"3983cb80",
X"08a01133",
X"70832a70",
X"81065151",
X"55557380",
X"2ea63888",
X"0ba01634",
X"ecae3f8c",
X"170883c0",
X"80082794",
X"38ff8077",
X"348e3977",
X"53805280",
X"51fa8b3f",
X"ff907734",
X"83cb8008",
X"a0113370",
X"832a7081",
X"06515155",
X"5573802e",
X"8638880b",
X"a0163489",
X"3d0d04f6",
X"3d0d02b3",
X"05330284",
X"05b70533",
X"5b5b800b",
X"83cb8c70",
X"84127274",
X"5d59575b",
X"58568315",
X"33537280",
X"2e80f338",
X"7333537a",
X"732e0981",
X"0680e738",
X"81143353",
X"79732e09",
X"810680da",
X"38805574",
X"81c42983",
X"cb900570",
X"33831b33",
X"58555373",
X"762e0981",
X"068a3881",
X"13335273",
X"51ff9c3f",
X"81157081",
X"ff065653",
X"8f7527d3",
X"38800b83",
X"cb881970",
X"08565455",
X"73752e91",
X"38725184",
X"14085372",
X"2d83c080",
X"0881ff06",
X"55800b83",
X"18347453",
X"a0398116",
X"81c41981",
X"c41781c4",
X"1781c41d",
X"81c41c5c",
X"5d575759",
X"568f7625",
X"fee83880",
X"537283c0",
X"800c8c3d",
X"0d04f83d",
X"0d02ae05",
X"227d5957",
X"80568155",
X"80548653",
X"8180527a",
X"51f5953f",
X"83c08008",
X"81ff0683",
X"c0800c8a",
X"3d0d04f7",
X"3d0d02b2",
X"05220284",
X"05b70533",
X"605a5b57",
X"80568255",
X"79548653",
X"8180527b",
X"51f4e53f",
X"83c08008",
X"81ff0683",
X"c0800c8b",
X"3d0d04f8",
X"3d0d02af",
X"05335980",
X"58805780",
X"56805578",
X"54895380",
X"527a51f4",
X"bb3f83c0",
X"800881ff",
X"0683c080",
X"0c8a3d0d",
X"04000000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002b20",
X"00002b61",
X"00002b83",
X"00002baa",
X"00002baa",
X"00002baa",
X"00002baa",
X"00002c1b",
X"00002c6d",
X"000041aa",
X"000049ee",
X"00004aa7",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3f00",
X"0c0c4000",
X"0a0a4100",
X"0b0b4100",
X"07074100",
X"0a0b4300",
X"080b4200",
X"04044500",
X"05054400",
X"06060004",
X"08080004",
X"09090004",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"00005733",
X"00005a3a",
X"00005846",
X"00005a3a",
X"00005883",
X"000058d4",
X"00005913",
X"0000591c",
X"00005a3a",
X"00005a3a",
X"00005a3a",
X"00005a3a",
X"00005925",
X"0000592d",
X"00005934",
X"00005b3a",
X"00005c33",
X"00005d47",
X"0000603d",
X"00006058",
X"00006044",
X"00006058",
X"0000605f",
X"0000606a",
X"00006071",
X"25732025",
X"73000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"66726565",
X"7a65722e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"6e616d65",
X"20000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00006ca8",
X"00006cac",
X"00006cb4",
X"00006cc0",
X"00006ccc",
X"00006cd8",
X"00006ce4",
X"00006ce8",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00006c44",
X"00006a98",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"69383030",
X"00000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
