---------------------------------------------------------------------------
-- (c) 2013 mark watson
-- I am happy for anyone to use this for non-commercial use.
-- If my vhdl files are used commercially or otherwise sold,
-- please contact me for explicit permission at scrameta (gmail).
-- This applies for source and binary form and derived works.
---------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY gtia_palette IS
PORT 
( 
	ATARI_COLOUR : IN STD_LOGIC_VECTOR(7 downto 0);
	PAL : IN STD_LOGIC;
	
	R_next : OUT STD_LOGIC_VECTOR(7 downto 0);
	G_next : OUT STD_LOGIC_VECTOR(7 downto 0);
	B_next : OUT STD_LOGIC_VECTOR(7 downto 0)
);
END gtia_palette;

ARCHITECTURE vhdl OF gtia_palette IS
begin
		--altirra_pal_default.pal
		process(atari_colour)
		begin
			case atari_colour is
				when X"00" =>
					R_next <= X"00";
					G_next <= X"00";
					B_next <= X"00";
				when X"01" =>
					R_next <= X"11";
					G_next <= X"11";
					B_next <= X"11";
				when X"02" =>
					R_next <= X"22";
					G_next <= X"22";
					B_next <= X"22";
				when X"03" =>
					R_next <= X"33";
					G_next <= X"33";
					B_next <= X"33";
				when X"04" =>
					R_next <= X"44";
					G_next <= X"44";
					B_next <= X"44";
				when X"05" =>
					R_next <= X"55";
					G_next <= X"55";
					B_next <= X"55";
				when X"06" =>
					R_next <= X"66";
					G_next <= X"66";
					B_next <= X"66";
				when X"07" =>
					R_next <= X"77";
					G_next <= X"77";
					B_next <= X"77";
				when X"08" =>
					R_next <= X"88";
					G_next <= X"88";
					B_next <= X"88";
				when X"09" =>
					R_next <= X"99";
					G_next <= X"99";
					B_next <= X"99";
				when X"0a" =>
					R_next <= X"aa";
					G_next <= X"aa";
					B_next <= X"aa";
				when X"0b" =>
					R_next <= X"bb";
					G_next <= X"bb";
					B_next <= X"bb";
				when X"0c" =>
					R_next <= X"cc";
					G_next <= X"cc";
					B_next <= X"cc";
				when X"0d" =>
					R_next <= X"dd";
					G_next <= X"dd";
					B_next <= X"dd";
				when X"0e" =>
					R_next <= X"ee";
					G_next <= X"ee";
					B_next <= X"ee";
				when X"0f" =>
					R_next <= X"ff";
					G_next <= X"ff";
					B_next <= X"ff";
				when X"10" =>
					R_next <= X"3f";
					G_next <= X"00";
					B_next <= X"00";
				when X"11" =>
					R_next <= X"50";
					G_next <= X"05";
					B_next <= X"00";
				when X"12" =>
					R_next <= X"61";
					G_next <= X"16";
					B_next <= X"00";
				when X"13" =>
					R_next <= X"72";
					G_next <= X"27";
					B_next <= X"00";
				when X"14" =>
					R_next <= X"83";
					G_next <= X"38";
					B_next <= X"00";
				when X"15" =>
					R_next <= X"94";
					G_next <= X"49";
					B_next <= X"00";
				when X"16" =>
					R_next <= X"a5";
					G_next <= X"5a";
					B_next <= X"01";
				when X"17" =>
					R_next <= X"b6";
					G_next <= X"6b";
					B_next <= X"12";
				when X"18" =>
					R_next <= X"c7";
					G_next <= X"7c";
					B_next <= X"23";
				when X"19" =>
					R_next <= X"d8";
					G_next <= X"8d";
					B_next <= X"34";
				when X"1a" =>
					R_next <= X"e9";
					G_next <= X"9e";
					B_next <= X"45";
				when X"1b" =>
					R_next <= X"fa";
					G_next <= X"af";
					B_next <= X"56";
				when X"1c" =>
					R_next <= X"ff";
					G_next <= X"c0";
					B_next <= X"67";
				when X"1d" =>
					R_next <= X"ff";
					G_next <= X"d1";
					B_next <= X"78";
				when X"1e" =>
					R_next <= X"ff";
					G_next <= X"e2";
					B_next <= X"89";
				when X"1f" =>
					R_next <= X"ff";
					G_next <= X"f3";
					B_next <= X"9a";
				when X"20" =>
					R_next <= X"50";
					G_next <= X"00";
					B_next <= X"00";
				when X"21" =>
					R_next <= X"61";
					G_next <= X"00";
					B_next <= X"00";
				when X"22" =>
					R_next <= X"72";
					G_next <= X"03";
					B_next <= X"00";
				when X"23" =>
					R_next <= X"83";
					G_next <= X"14";
					B_next <= X"03";
				when X"24" =>
					R_next <= X"94";
					G_next <= X"25";
					B_next <= X"14";
				when X"25" =>
					R_next <= X"a5";
					G_next <= X"36";
					B_next <= X"25";
				when X"26" =>
					R_next <= X"b6";
					G_next <= X"47";
					B_next <= X"36";
				when X"27" =>
					R_next <= X"c7";
					G_next <= X"58";
					B_next <= X"47";
				when X"28" =>
					R_next <= X"d8";
					G_next <= X"69";
					B_next <= X"58";
				when X"29" =>
					R_next <= X"e9";
					G_next <= X"7a";
					B_next <= X"69";
				when X"2a" =>
					R_next <= X"fa";
					G_next <= X"8b";
					B_next <= X"7a";
				when X"2b" =>
					R_next <= X"ff";
					G_next <= X"9c";
					B_next <= X"8b";
				when X"2c" =>
					R_next <= X"ff";
					G_next <= X"ad";
					B_next <= X"9c";
				when X"2d" =>
					R_next <= X"ff";
					G_next <= X"be";
					B_next <= X"ad";
				when X"2e" =>
					R_next <= X"ff";
					G_next <= X"cf";
					B_next <= X"be";
				when X"2f" =>
					R_next <= X"ff";
					G_next <= X"e0";
					B_next <= X"cf";
				when X"30" =>
					R_next <= X"54";
					G_next <= X"00";
					B_next <= X"03";
				when X"31" =>
					R_next <= X"65";
					G_next <= X"00";
					B_next <= X"14";
				when X"32" =>
					R_next <= X"76";
					G_next <= X"00";
					B_next <= X"25";
				when X"33" =>
					R_next <= X"87";
					G_next <= X"08";
					B_next <= X"36";
				when X"34" =>
					R_next <= X"98";
					G_next <= X"19";
					B_next <= X"47";
				when X"35" =>
					R_next <= X"a9";
					G_next <= X"2a";
					B_next <= X"58";
				when X"36" =>
					R_next <= X"ba";
					G_next <= X"3b";
					B_next <= X"69";
				when X"37" =>
					R_next <= X"cb";
					G_next <= X"4c";
					B_next <= X"7a";
				when X"38" =>
					R_next <= X"dc";
					G_next <= X"5d";
					B_next <= X"8b";
				when X"39" =>
					R_next <= X"ed";
					G_next <= X"6e";
					B_next <= X"9c";
				when X"3a" =>
					R_next <= X"fe";
					G_next <= X"7f";
					B_next <= X"ad";
				when X"3b" =>
					R_next <= X"ff";
					G_next <= X"90";
					B_next <= X"be";
				when X"3c" =>
					R_next <= X"ff";
					G_next <= X"a1";
					B_next <= X"cf";
				when X"3d" =>
					R_next <= X"ff";
					G_next <= X"b2";
					B_next <= X"e0";
				when X"3e" =>
					R_next <= X"ff";
					G_next <= X"c3";
					B_next <= X"f1";
				when X"3f" =>
					R_next <= X"ff";
					G_next <= X"d4";
					B_next <= X"ff";
				when X"40" =>
					R_next <= X"4f";
					G_next <= X"00";
					B_next <= X"35";
				when X"41" =>
					R_next <= X"60";
					G_next <= X"00";
					B_next <= X"46";
				when X"42" =>
					R_next <= X"71";
					G_next <= X"00";
					B_next <= X"57";
				when X"43" =>
					R_next <= X"82";
					G_next <= X"01";
					B_next <= X"68";
				when X"44" =>
					R_next <= X"93";
					G_next <= X"12";
					B_next <= X"79";
				when X"45" =>
					R_next <= X"a4";
					G_next <= X"23";
					B_next <= X"8a";
				when X"46" =>
					R_next <= X"b5";
					G_next <= X"34";
					B_next <= X"9b";
				when X"47" =>
					R_next <= X"c6";
					G_next <= X"45";
					B_next <= X"ac";
				when X"48" =>
					R_next <= X"d7";
					G_next <= X"56";
					B_next <= X"bd";
				when X"49" =>
					R_next <= X"e8";
					G_next <= X"67";
					B_next <= X"ce";
				when X"4a" =>
					R_next <= X"f9";
					G_next <= X"78";
					B_next <= X"df";
				when X"4b" =>
					R_next <= X"ff";
					G_next <= X"89";
					B_next <= X"f0";
				when X"4c" =>
					R_next <= X"ff";
					G_next <= X"9a";
					B_next <= X"ff";
				when X"4d" =>
					R_next <= X"ff";
					G_next <= X"ab";
					B_next <= X"ff";
				when X"4e" =>
					R_next <= X"ff";
					G_next <= X"bc";
					B_next <= X"ff";
				when X"4f" =>
					R_next <= X"ff";
					G_next <= X"cd";
					B_next <= X"ff";
				when X"50" =>
					R_next <= X"3d";
					G_next <= X"00";
					B_next <= X"68";
				when X"51" =>
					R_next <= X"4e";
					G_next <= X"00";
					B_next <= X"79";
				when X"52" =>
					R_next <= X"5f";
					G_next <= X"00";
					B_next <= X"8a";
				when X"53" =>
					R_next <= X"70";
					G_next <= X"00";
					B_next <= X"9b";
				when X"54" =>
					R_next <= X"81";
					G_next <= X"11";
					B_next <= X"ac";
				when X"55" =>
					R_next <= X"92";
					G_next <= X"22";
					B_next <= X"bd";
				when X"56" =>
					R_next <= X"a3";
					G_next <= X"33";
					B_next <= X"ce";
				when X"57" =>
					R_next <= X"b4";
					G_next <= X"44";
					B_next <= X"df";
				when X"58" =>
					R_next <= X"c5";
					G_next <= X"55";
					B_next <= X"f0";
				when X"59" =>
					R_next <= X"d6";
					G_next <= X"66";
					B_next <= X"ff";
				when X"5a" =>
					R_next <= X"e7";
					G_next <= X"77";
					B_next <= X"ff";
				when X"5b" =>
					R_next <= X"f8";
					G_next <= X"88";
					B_next <= X"ff";
				when X"5c" =>
					R_next <= X"ff";
					G_next <= X"99";
					B_next <= X"ff";
				when X"5d" =>
					R_next <= X"ff";
					G_next <= X"aa";
					B_next <= X"ff";
				when X"5e" =>
					R_next <= X"ff";
					G_next <= X"bb";
					B_next <= X"ff";
				when X"5f" =>
					R_next <= X"ff";
					G_next <= X"cc";
					B_next <= X"ff";
				when X"60" =>
					R_next <= X"20";
					G_next <= X"00";
					B_next <= X"8b";
				when X"61" =>
					R_next <= X"31";
					G_next <= X"00";
					B_next <= X"9c";
				when X"62" =>
					R_next <= X"42";
					G_next <= X"00";
					B_next <= X"ad";
				when X"63" =>
					R_next <= X"53";
					G_next <= X"08";
					B_next <= X"be";
				when X"64" =>
					R_next <= X"64";
					G_next <= X"19";
					B_next <= X"cf";
				when X"65" =>
					R_next <= X"75";
					G_next <= X"2a";
					B_next <= X"e0";
				when X"66" =>
					R_next <= X"86";
					G_next <= X"3b";
					B_next <= X"f1";
				when X"67" =>
					R_next <= X"97";
					G_next <= X"4c";
					B_next <= X"ff";
				when X"68" =>
					R_next <= X"a8";
					G_next <= X"5d";
					B_next <= X"ff";
				when X"69" =>
					R_next <= X"b9";
					G_next <= X"6e";
					B_next <= X"ff";
				when X"6a" =>
					R_next <= X"ca";
					G_next <= X"7f";
					B_next <= X"ff";
				when X"6b" =>
					R_next <= X"db";
					G_next <= X"90";
					B_next <= X"ff";
				when X"6c" =>
					R_next <= X"ec";
					G_next <= X"a1";
					B_next <= X"ff";
				when X"6d" =>
					R_next <= X"fd";
					G_next <= X"b2";
					B_next <= X"ff";
				when X"6e" =>
					R_next <= X"ff";
					G_next <= X"c3";
					B_next <= X"ff";
				when X"6f" =>
					R_next <= X"ff";
					G_next <= X"d4";
					B_next <= X"ff";
				when X"70" =>
					R_next <= X"00";
					G_next <= X"00";
					B_next <= X"89";
				when X"71" =>
					R_next <= X"00";
					G_next <= X"08";
					B_next <= X"9a";
				when X"72" =>
					R_next <= X"00";
					G_next <= X"19";
					B_next <= X"ab";
				when X"73" =>
					R_next <= X"10";
					G_next <= X"2a";
					B_next <= X"bc";
				when X"74" =>
					R_next <= X"21";
					G_next <= X"3b";
					B_next <= X"cd";
				when X"75" =>
					R_next <= X"32";
					G_next <= X"4c";
					B_next <= X"de";
				when X"76" =>
					R_next <= X"43";
					G_next <= X"5d";
					B_next <= X"ef";
				when X"77" =>
					R_next <= X"54";
					G_next <= X"6e";
					B_next <= X"ff";
				when X"78" =>
					R_next <= X"65";
					G_next <= X"7f";
					B_next <= X"ff";
				when X"79" =>
					R_next <= X"76";
					G_next <= X"90";
					B_next <= X"ff";
				when X"7a" =>
					R_next <= X"87";
					G_next <= X"a1";
					B_next <= X"ff";
				when X"7b" =>
					R_next <= X"98";
					G_next <= X"b2";
					B_next <= X"ff";
				when X"7c" =>
					R_next <= X"a9";
					G_next <= X"c3";
					B_next <= X"ff";
				when X"7d" =>
					R_next <= X"ba";
					G_next <= X"d4";
					B_next <= X"ff";
				when X"7e" =>
					R_next <= X"cb";
					G_next <= X"e5";
					B_next <= X"ff";
				when X"7f" =>
					R_next <= X"dc";
					G_next <= X"f6";
					B_next <= X"ff";
				when X"80" =>
					R_next <= X"00";
					G_next <= X"0c";
					B_next <= X"65";
				when X"81" =>
					R_next <= X"00";
					G_next <= X"1d";
					B_next <= X"76";
				when X"82" =>
					R_next <= X"00";
					G_next <= X"2e";
					B_next <= X"87";
				when X"83" =>
					R_next <= X"00";
					G_next <= X"3f";
					B_next <= X"98";
				when X"84" =>
					R_next <= X"05";
					G_next <= X"50";
					B_next <= X"a9";
				when X"85" =>
					R_next <= X"16";
					G_next <= X"61";
					B_next <= X"ba";
				when X"86" =>
					R_next <= X"27";
					G_next <= X"72";
					B_next <= X"cb";
				when X"87" =>
					R_next <= X"38";
					G_next <= X"83";
					B_next <= X"dc";
				when X"88" =>
					R_next <= X"49";
					G_next <= X"94";
					B_next <= X"ed";
				when X"89" =>
					R_next <= X"5a";
					G_next <= X"a5";
					B_next <= X"fe";
				when X"8a" =>
					R_next <= X"6b";
					G_next <= X"b6";
					B_next <= X"ff";
				when X"8b" =>
					R_next <= X"7c";
					G_next <= X"c7";
					B_next <= X"ff";
				when X"8c" =>
					R_next <= X"8d";
					G_next <= X"d8";
					B_next <= X"ff";
				when X"8d" =>
					R_next <= X"9e";
					G_next <= X"e9";
					B_next <= X"ff";
				when X"8e" =>
					R_next <= X"af";
					G_next <= X"fa";
					B_next <= X"ff";
				when X"8f" =>
					R_next <= X"c0";
					G_next <= X"ff";
					B_next <= X"ff";
				when X"90" =>
					R_next <= X"00";
					G_next <= X"1f";
					B_next <= X"30";
				when X"91" =>
					R_next <= X"00";
					G_next <= X"30";
					B_next <= X"41";
				when X"92" =>
					R_next <= X"00";
					G_next <= X"41";
					B_next <= X"52";
				when X"93" =>
					R_next <= X"00";
					G_next <= X"52";
					B_next <= X"63";
				when X"94" =>
					R_next <= X"00";
					G_next <= X"63";
					B_next <= X"74";
				when X"95" =>
					R_next <= X"05";
					G_next <= X"74";
					B_next <= X"85";
				when X"96" =>
					R_next <= X"16";
					G_next <= X"85";
					B_next <= X"96";
				when X"97" =>
					R_next <= X"27";
					G_next <= X"96";
					B_next <= X"a7";
				when X"98" =>
					R_next <= X"38";
					G_next <= X"a7";
					B_next <= X"b8";
				when X"99" =>
					R_next <= X"49";
					G_next <= X"b8";
					B_next <= X"c9";
				when X"9a" =>
					R_next <= X"5a";
					G_next <= X"c9";
					B_next <= X"da";
				when X"9b" =>
					R_next <= X"6b";
					G_next <= X"da";
					B_next <= X"eb";
				when X"9c" =>
					R_next <= X"7c";
					G_next <= X"eb";
					B_next <= X"fc";
				when X"9d" =>
					R_next <= X"8d";
					G_next <= X"fc";
					B_next <= X"ff";
				when X"9e" =>
					R_next <= X"9e";
					G_next <= X"ff";
					B_next <= X"ff";
				when X"9f" =>
					R_next <= X"af";
					G_next <= X"ff";
					B_next <= X"ff";
				when X"a0" =>
					R_next <= X"00";
					G_next <= X"2b";
					B_next <= X"00";
				when X"a1" =>
					R_next <= X"00";
					G_next <= X"3c";
					B_next <= X"0e";
				when X"a2" =>
					R_next <= X"00";
					G_next <= X"4d";
					B_next <= X"1f";
				when X"a3" =>
					R_next <= X"00";
					G_next <= X"5e";
					B_next <= X"30";
				when X"a4" =>
					R_next <= X"00";
					G_next <= X"6f";
					B_next <= X"41";
				when X"a5" =>
					R_next <= X"01";
					G_next <= X"80";
					B_next <= X"52";
				when X"a6" =>
					R_next <= X"12";
					G_next <= X"91";
					B_next <= X"63";
				when X"a7" =>
					R_next <= X"23";
					G_next <= X"a2";
					B_next <= X"74";
				when X"a8" =>
					R_next <= X"34";
					G_next <= X"b3";
					B_next <= X"85";
				when X"a9" =>
					R_next <= X"45";
					G_next <= X"c4";
					B_next <= X"96";
				when X"aa" =>
					R_next <= X"56";
					G_next <= X"d5";
					B_next <= X"a7";
				when X"ab" =>
					R_next <= X"67";
					G_next <= X"e6";
					B_next <= X"b8";
				when X"ac" =>
					R_next <= X"78";
					G_next <= X"f7";
					B_next <= X"c9";
				when X"ad" =>
					R_next <= X"89";
					G_next <= X"ff";
					B_next <= X"da";
				when X"ae" =>
					R_next <= X"9a";
					G_next <= X"ff";
					B_next <= X"eb";
				when X"af" =>
					R_next <= X"ab";
					G_next <= X"ff";
					B_next <= X"fc";
				when X"b0" =>
					R_next <= X"00";
					G_next <= X"33";
					B_next <= X"00";
				when X"b1" =>
					R_next <= X"00";
					G_next <= X"44";
					B_next <= X"00";
				when X"b2" =>
					R_next <= X"00";
					G_next <= X"55";
					B_next <= X"00";
				when X"b3" =>
					R_next <= X"00";
					G_next <= X"66";
					B_next <= X"00";
				when X"b4" =>
					R_next <= X"07";
					G_next <= X"77";
					B_next <= X"00";
				when X"b5" =>
					R_next <= X"18";
					G_next <= X"88";
					B_next <= X"00";
				when X"b6" =>
					R_next <= X"29";
					G_next <= X"99";
					B_next <= X"00";
				when X"b7" =>
					R_next <= X"3a";
					G_next <= X"aa";
					B_next <= X"0f";
				when X"b8" =>
					R_next <= X"4b";
					G_next <= X"bb";
					B_next <= X"20";
				when X"b9" =>
					R_next <= X"5c";
					G_next <= X"cc";
					B_next <= X"31";
				when X"ba" =>
					R_next <= X"6d";
					G_next <= X"dd";
					B_next <= X"42";
				when X"bb" =>
					R_next <= X"7e";
					G_next <= X"ee";
					B_next <= X"53";
				when X"bc" =>
					R_next <= X"8f";
					G_next <= X"ff";
					B_next <= X"64";
				when X"bd" =>
					R_next <= X"a0";
					G_next <= X"ff";
					B_next <= X"75";
				when X"be" =>
					R_next <= X"b1";
					G_next <= X"ff";
					B_next <= X"86";
				when X"bf" =>
					R_next <= X"c2";
					G_next <= X"ff";
					B_next <= X"97";
				when X"c0" =>
					R_next <= X"00";
					G_next <= X"2b";
					B_next <= X"00";
				when X"c1" =>
					R_next <= X"00";
					G_next <= X"3c";
					B_next <= X"00";
				when X"c2" =>
					R_next <= X"02";
					G_next <= X"4d";
					B_next <= X"00";
				when X"c3" =>
					R_next <= X"13";
					G_next <= X"5e";
					B_next <= X"00";
				when X"c4" =>
					R_next <= X"24";
					G_next <= X"6f";
					B_next <= X"00";
				when X"c5" =>
					R_next <= X"35";
					G_next <= X"80";
					B_next <= X"00";
				when X"c6" =>
					R_next <= X"46";
					G_next <= X"91";
					B_next <= X"00";
				when X"c7" =>
					R_next <= X"57";
					G_next <= X"a2";
					B_next <= X"00";
				when X"c8" =>
					R_next <= X"68";
					G_next <= X"b3";
					B_next <= X"00";
				when X"c9" =>
					R_next <= X"79";
					G_next <= X"c4";
					B_next <= X"0e";
				when X"ca" =>
					R_next <= X"8a";
					G_next <= X"d5";
					B_next <= X"1f";
				when X"cb" =>
					R_next <= X"9b";
					G_next <= X"e6";
					B_next <= X"30";
				when X"cc" =>
					R_next <= X"ac";
					G_next <= X"f7";
					B_next <= X"41";
				when X"cd" =>
					R_next <= X"bd";
					G_next <= X"ff";
					B_next <= X"52";
				when X"ce" =>
					R_next <= X"ce";
					G_next <= X"ff";
					B_next <= X"63";
				when X"cf" =>
					R_next <= X"df";
					G_next <= X"ff";
					B_next <= X"74";
				when X"d0" =>
					R_next <= X"01";
					G_next <= X"1c";
					B_next <= X"00";
				when X"d1" =>
					R_next <= X"12";
					G_next <= X"2d";
					B_next <= X"00";
				when X"d2" =>
					R_next <= X"23";
					G_next <= X"3e";
					B_next <= X"00";
				when X"d3" =>
					R_next <= X"34";
					G_next <= X"4f";
					B_next <= X"00";
				when X"d4" =>
					R_next <= X"45";
					G_next <= X"60";
					B_next <= X"00";
				when X"d5" =>
					R_next <= X"56";
					G_next <= X"71";
					B_next <= X"00";
				when X"d6" =>
					R_next <= X"67";
					G_next <= X"82";
					B_next <= X"00";
				when X"d7" =>
					R_next <= X"78";
					G_next <= X"93";
					B_next <= X"00";
				when X"d8" =>
					R_next <= X"89";
					G_next <= X"a4";
					B_next <= X"00";
				when X"d9" =>
					R_next <= X"9a";
					G_next <= X"b5";
					B_next <= X"03";
				when X"da" =>
					R_next <= X"ab";
					G_next <= X"c6";
					B_next <= X"14";
				when X"db" =>
					R_next <= X"bc";
					G_next <= X"d7";
					B_next <= X"25";
				when X"dc" =>
					R_next <= X"cd";
					G_next <= X"e8";
					B_next <= X"36";
				when X"dd" =>
					R_next <= X"de";
					G_next <= X"f9";
					B_next <= X"47";
				when X"de" =>
					R_next <= X"ef";
					G_next <= X"ff";
					B_next <= X"58";
				when X"df" =>
					R_next <= X"ff";
					G_next <= X"ff";
					B_next <= X"69";
				when X"e0" =>
					R_next <= X"23";
					G_next <= X"09";
					B_next <= X"00";
				when X"e1" =>
					R_next <= X"34";
					G_next <= X"1a";
					B_next <= X"00";
				when X"e2" =>
					R_next <= X"45";
					G_next <= X"2b";
					B_next <= X"00";
				when X"e3" =>
					R_next <= X"56";
					G_next <= X"3c";
					B_next <= X"00";
				when X"e4" =>
					R_next <= X"67";
					G_next <= X"4d";
					B_next <= X"00";
				when X"e5" =>
					R_next <= X"78";
					G_next <= X"5e";
					B_next <= X"00";
				when X"e6" =>
					R_next <= X"89";
					G_next <= X"6f";
					B_next <= X"00";
				when X"e7" =>
					R_next <= X"9a";
					G_next <= X"80";
					B_next <= X"00";
				when X"e8" =>
					R_next <= X"ab";
					G_next <= X"91";
					B_next <= X"00";
				when X"e9" =>
					R_next <= X"bc";
					G_next <= X"a2";
					B_next <= X"10";
				when X"ea" =>
					R_next <= X"cd";
					G_next <= X"b3";
					B_next <= X"21";
				when X"eb" =>
					R_next <= X"de";
					G_next <= X"c4";
					B_next <= X"32";
				when X"ec" =>
					R_next <= X"ef";
					G_next <= X"d5";
					B_next <= X"43";
				when X"ed" =>
					R_next <= X"ff";
					G_next <= X"e6";
					B_next <= X"54";
				when X"ee" =>
					R_next <= X"ff";
					G_next <= X"f7";
					B_next <= X"65";
				when X"ef" =>
					R_next <= X"ff";
					G_next <= X"ff";
					B_next <= X"76";
				when X"f0" =>
					R_next <= X"3f";
					G_next <= X"00";
					B_next <= X"00";
				when X"f1" =>
					R_next <= X"50";
					G_next <= X"05";
					B_next <= X"00";
				when X"f2" =>
					R_next <= X"61";
					G_next <= X"16";
					B_next <= X"00";
				when X"f3" =>
					R_next <= X"72";
					G_next <= X"27";
					B_next <= X"00";
				when X"f4" =>
					R_next <= X"83";
					G_next <= X"38";
					B_next <= X"00";
				when X"f5" =>
					R_next <= X"94";
					G_next <= X"49";
					B_next <= X"00";
				when X"f6" =>
					R_next <= X"a5";
					G_next <= X"5a";
					B_next <= X"01";
				when X"f7" =>
					R_next <= X"b6";
					G_next <= X"6b";
					B_next <= X"12";
				when X"f8" =>
					R_next <= X"c7";
					G_next <= X"7c";
					B_next <= X"23";
				when X"f9" =>
					R_next <= X"d8";
					G_next <= X"8d";
					B_next <= X"34";
				when X"fa" =>
					R_next <= X"e9";
					G_next <= X"9e";
					B_next <= X"45";
				when X"fb" =>
					R_next <= X"fa";
					G_next <= X"af";
					B_next <= X"56";
				when X"fc" =>
					R_next <= X"ff";
					G_next <= X"c0";
					B_next <= X"67";
				when X"fd" =>
					R_next <= X"ff";
					G_next <= X"d1";
					B_next <= X"78";
				when X"fe" =>
					R_next <= X"ff";
					G_next <= X"e2";
					B_next <= X"89";
				when X"ff" =>
					R_next <= X"ff";
					G_next <= X"f3";
					B_next <= X"9a";
				when others =>
					--nop
			end case;

		if (pal = '0') then
		--altirra_ntsc_default.pal
			case atari_colour is
				when X"00" =>
					R_next <= X"00";
					G_next <= X"00";
					B_next <= X"00";
				when X"01" =>
					R_next <= X"11";
					G_next <= X"11";
					B_next <= X"11";
				when X"02" =>
					R_next <= X"22";
					G_next <= X"22";
					B_next <= X"22";
				when X"03" =>
					R_next <= X"33";
					G_next <= X"33";
					B_next <= X"33";
				when X"04" =>
					R_next <= X"44";
					G_next <= X"44";
					B_next <= X"44";
				when X"05" =>
					R_next <= X"55";
					G_next <= X"55";
					B_next <= X"55";
				when X"06" =>
					R_next <= X"66";
					G_next <= X"66";
					B_next <= X"66";
				when X"07" =>
					R_next <= X"77";
					G_next <= X"77";
					B_next <= X"77";
				when X"08" =>
					R_next <= X"88";
					G_next <= X"88";
					B_next <= X"88";
				when X"09" =>
					R_next <= X"99";
					G_next <= X"99";
					B_next <= X"99";
				when X"0a" =>
					R_next <= X"aa";
					G_next <= X"aa";
					B_next <= X"aa";
				when X"0b" =>
					R_next <= X"bb";
					G_next <= X"bb";
					B_next <= X"bb";
				when X"0c" =>
					R_next <= X"cc";
					G_next <= X"cc";
					B_next <= X"cc";
				when X"0d" =>
					R_next <= X"dd";
					G_next <= X"dd";
					B_next <= X"dd";
				when X"0e" =>
					R_next <= X"ee";
					G_next <= X"ee";
					B_next <= X"ee";
				when X"0f" =>
					R_next <= X"ff";
					G_next <= X"ff";
					B_next <= X"ff";
				when X"10" =>
					R_next <= X"09";
					G_next <= X"19";
					B_next <= X"00";
				when X"11" =>
					R_next <= X"1a";
					G_next <= X"2a";
					B_next <= X"00";
				when X"12" =>
					R_next <= X"2b";
					G_next <= X"3b";
					B_next <= X"00";
				when X"13" =>
					R_next <= X"3c";
					G_next <= X"4c";
					B_next <= X"00";
				when X"14" =>
					R_next <= X"4d";
					G_next <= X"5d";
					B_next <= X"00";
				when X"15" =>
					R_next <= X"5e";
					G_next <= X"6e";
					B_next <= X"00";
				when X"16" =>
					R_next <= X"6f";
					G_next <= X"7f";
					B_next <= X"00";
				when X"17" =>
					R_next <= X"80";
					G_next <= X"90";
					B_next <= X"00";
				when X"18" =>
					R_next <= X"91";
					G_next <= X"a1";
					B_next <= X"00";
				when X"19" =>
					R_next <= X"a2";
					G_next <= X"b2";
					B_next <= X"01";
				when X"1a" =>
					R_next <= X"b3";
					G_next <= X"c3";
					B_next <= X"12";
				when X"1b" =>
					R_next <= X"c4";
					G_next <= X"d4";
					B_next <= X"23";
				when X"1c" =>
					R_next <= X"d5";
					G_next <= X"e5";
					B_next <= X"34";
				when X"1d" =>
					R_next <= X"e6";
					G_next <= X"f6";
					B_next <= X"45";
				when X"1e" =>
					R_next <= X"f7";
					G_next <= X"ff";
					B_next <= X"56";
				when X"1f" =>
					R_next <= X"ff";
					G_next <= X"ff";
					B_next <= X"67";
				when X"20" =>
					R_next <= X"30";
					G_next <= X"00";
					B_next <= X"00";
				when X"21" =>
					R_next <= X"41";
					G_next <= X"11";
					B_next <= X"00";
				when X"22" =>
					R_next <= X"52";
					G_next <= X"22";
					B_next <= X"00";
				when X"23" =>
					R_next <= X"63";
					G_next <= X"33";
					B_next <= X"00";
				when X"24" =>
					R_next <= X"74";
					G_next <= X"44";
					B_next <= X"00";
				when X"25" =>
					R_next <= X"85";
					G_next <= X"55";
					B_next <= X"00";
				when X"26" =>
					R_next <= X"96";
					G_next <= X"66";
					B_next <= X"00";
				when X"27" =>
					R_next <= X"a7";
					G_next <= X"77";
					B_next <= X"00";
				when X"28" =>
					R_next <= X"b8";
					G_next <= X"88";
					B_next <= X"09";
				when X"29" =>
					R_next <= X"c9";
					G_next <= X"99";
					B_next <= X"1a";
				when X"2a" =>
					R_next <= X"da";
					G_next <= X"aa";
					B_next <= X"2b";
				when X"2b" =>
					R_next <= X"eb";
					G_next <= X"bb";
					B_next <= X"3c";
				when X"2c" =>
					R_next <= X"fc";
					G_next <= X"cc";
					B_next <= X"4d";
				when X"2d" =>
					R_next <= X"ff";
					G_next <= X"dd";
					B_next <= X"5e";
				when X"2e" =>
					R_next <= X"ff";
					G_next <= X"ee";
					B_next <= X"6f";
				when X"2f" =>
					R_next <= X"ff";
					G_next <= X"ff";
					B_next <= X"80";
				when X"30" =>
					R_next <= X"4b";
					G_next <= X"00";
					B_next <= X"00";
				when X"31" =>
					R_next <= X"5c";
					G_next <= X"00";
					B_next <= X"00";
				when X"32" =>
					R_next <= X"6d";
					G_next <= X"0a";
					B_next <= X"00";
				when X"33" =>
					R_next <= X"7e";
					G_next <= X"1b";
					B_next <= X"00";
				when X"34" =>
					R_next <= X"8f";
					G_next <= X"2c";
					B_next <= X"00";
				when X"35" =>
					R_next <= X"a0";
					G_next <= X"3d";
					B_next <= X"0d";
				when X"36" =>
					R_next <= X"b1";
					G_next <= X"4e";
					B_next <= X"1e";
				when X"37" =>
					R_next <= X"c2";
					G_next <= X"5f";
					B_next <= X"2f";
				when X"38" =>
					R_next <= X"d3";
					G_next <= X"70";
					B_next <= X"40";
				when X"39" =>
					R_next <= X"e4";
					G_next <= X"81";
					B_next <= X"51";
				when X"3a" =>
					R_next <= X"f5";
					G_next <= X"92";
					B_next <= X"62";
				when X"3b" =>
					R_next <= X"ff";
					G_next <= X"a3";
					B_next <= X"73";
				when X"3c" =>
					R_next <= X"ff";
					G_next <= X"b4";
					B_next <= X"84";
				when X"3d" =>
					R_next <= X"ff";
					G_next <= X"c5";
					B_next <= X"95";
				when X"3e" =>
					R_next <= X"ff";
					G_next <= X"d6";
					B_next <= X"a6";
				when X"3f" =>
					R_next <= X"ff";
					G_next <= X"e7";
					B_next <= X"b7";
				when X"40" =>
					R_next <= X"55";
					G_next <= X"00";
					B_next <= X"00";
				when X"41" =>
					R_next <= X"66";
					G_next <= X"00";
					B_next <= X"10";
				when X"42" =>
					R_next <= X"77";
					G_next <= X"00";
					B_next <= X"21";
				when X"43" =>
					R_next <= X"88";
					G_next <= X"08";
					B_next <= X"32";
				when X"44" =>
					R_next <= X"99";
					G_next <= X"19";
					B_next <= X"43";
				when X"45" =>
					R_next <= X"aa";
					G_next <= X"2a";
					B_next <= X"54";
				when X"46" =>
					R_next <= X"bb";
					G_next <= X"3b";
					B_next <= X"65";
				when X"47" =>
					R_next <= X"cc";
					G_next <= X"4c";
					B_next <= X"76";
				when X"48" =>
					R_next <= X"dd";
					G_next <= X"5d";
					B_next <= X"87";
				when X"49" =>
					R_next <= X"ee";
					G_next <= X"6e";
					B_next <= X"98";
				when X"4a" =>
					R_next <= X"ff";
					G_next <= X"7f";
					B_next <= X"a9";
				when X"4b" =>
					R_next <= X"ff";
					G_next <= X"90";
					B_next <= X"ba";
				when X"4c" =>
					R_next <= X"ff";
					G_next <= X"a1";
					B_next <= X"cb";
				when X"4d" =>
					R_next <= X"ff";
					G_next <= X"b2";
					B_next <= X"dc";
				when X"4e" =>
					R_next <= X"ff";
					G_next <= X"c3";
					B_next <= X"ed";
				when X"4f" =>
					R_next <= X"ff";
					G_next <= X"d4";
					B_next <= X"fe";
				when X"50" =>
					R_next <= X"4c";
					G_next <= X"00";
					B_next <= X"47";
				when X"51" =>
					R_next <= X"5d";
					G_next <= X"00";
					B_next <= X"58";
				when X"52" =>
					R_next <= X"6e";
					G_next <= X"00";
					B_next <= X"69";
				when X"53" =>
					R_next <= X"7f";
					G_next <= X"00";
					B_next <= X"7a";
				when X"54" =>
					R_next <= X"90";
					G_next <= X"10";
					B_next <= X"8b";
				when X"55" =>
					R_next <= X"a1";
					G_next <= X"21";
					B_next <= X"9c";
				when X"56" =>
					R_next <= X"b2";
					G_next <= X"32";
					B_next <= X"ad";
				when X"57" =>
					R_next <= X"c3";
					G_next <= X"43";
					B_next <= X"be";
				when X"58" =>
					R_next <= X"d4";
					G_next <= X"54";
					B_next <= X"cf";
				when X"59" =>
					R_next <= X"e5";
					G_next <= X"65";
					B_next <= X"e0";
				when X"5a" =>
					R_next <= X"f6";
					G_next <= X"76";
					B_next <= X"f1";
				when X"5b" =>
					R_next <= X"ff";
					G_next <= X"87";
					B_next <= X"ff";
				when X"5c" =>
					R_next <= X"ff";
					G_next <= X"98";
					B_next <= X"ff";
				when X"5d" =>
					R_next <= X"ff";
					G_next <= X"a9";
					B_next <= X"ff";
				when X"5e" =>
					R_next <= X"ff";
					G_next <= X"ba";
					B_next <= X"ff";
				when X"5f" =>
					R_next <= X"ff";
					G_next <= X"cb";
					B_next <= X"ff";
				when X"60" =>
					R_next <= X"30";
					G_next <= X"00";
					B_next <= X"7e";
				when X"61" =>
					R_next <= X"41";
					G_next <= X"00";
					B_next <= X"8f";
				when X"62" =>
					R_next <= X"52";
					G_next <= X"00";
					B_next <= X"a0";
				when X"63" =>
					R_next <= X"63";
					G_next <= X"02";
					B_next <= X"b1";
				when X"64" =>
					R_next <= X"74";
					G_next <= X"13";
					B_next <= X"c2";
				when X"65" =>
					R_next <= X"85";
					G_next <= X"24";
					B_next <= X"d3";
				when X"66" =>
					R_next <= X"96";
					G_next <= X"35";
					B_next <= X"e4";
				when X"67" =>
					R_next <= X"a7";
					G_next <= X"46";
					B_next <= X"f5";
				when X"68" =>
					R_next <= X"b8";
					G_next <= X"57";
					B_next <= X"ff";
				when X"69" =>
					R_next <= X"c9";
					G_next <= X"68";
					B_next <= X"ff";
				when X"6a" =>
					R_next <= X"da";
					G_next <= X"79";
					B_next <= X"ff";
				when X"6b" =>
					R_next <= X"eb";
					G_next <= X"8a";
					B_next <= X"ff";
				when X"6c" =>
					R_next <= X"fc";
					G_next <= X"9b";
					B_next <= X"ff";
				when X"6d" =>
					R_next <= X"ff";
					G_next <= X"ac";
					B_next <= X"ff";
				when X"6e" =>
					R_next <= X"ff";
					G_next <= X"bd";
					B_next <= X"ff";
				when X"6f" =>
					R_next <= X"ff";
					G_next <= X"ce";
					B_next <= X"ff";
				when X"70" =>
					R_next <= X"0a";
					G_next <= X"00";
					B_next <= X"97";
				when X"71" =>
					R_next <= X"1b";
					G_next <= X"00";
					B_next <= X"a8";
				when X"72" =>
					R_next <= X"2c";
					G_next <= X"00";
					B_next <= X"b9";
				when X"73" =>
					R_next <= X"3d";
					G_next <= X"11";
					B_next <= X"ca";
				when X"74" =>
					R_next <= X"4e";
					G_next <= X"22";
					B_next <= X"db";
				when X"75" =>
					R_next <= X"5f";
					G_next <= X"33";
					B_next <= X"ec";
				when X"76" =>
					R_next <= X"70";
					G_next <= X"44";
					B_next <= X"fd";
				when X"77" =>
					R_next <= X"81";
					G_next <= X"55";
					B_next <= X"ff";
				when X"78" =>
					R_next <= X"92";
					G_next <= X"66";
					B_next <= X"ff";
				when X"79" =>
					R_next <= X"a3";
					G_next <= X"77";
					B_next <= X"ff";
				when X"7a" =>
					R_next <= X"b4";
					G_next <= X"88";
					B_next <= X"ff";
				when X"7b" =>
					R_next <= X"c5";
					G_next <= X"99";
					B_next <= X"ff";
				when X"7c" =>
					R_next <= X"d6";
					G_next <= X"aa";
					B_next <= X"ff";
				when X"7d" =>
					R_next <= X"e7";
					G_next <= X"bb";
					B_next <= X"ff";
				when X"7e" =>
					R_next <= X"f8";
					G_next <= X"cc";
					B_next <= X"ff";
				when X"7f" =>
					R_next <= X"ff";
					G_next <= X"dd";
					B_next <= X"ff";
				when X"80" =>
					R_next <= X"00";
					G_next <= X"00";
					B_next <= X"8e";
				when X"81" =>
					R_next <= X"00";
					G_next <= X"05";
					B_next <= X"9f";
				when X"82" =>
					R_next <= X"03";
					G_next <= X"16";
					B_next <= X"b0";
				when X"83" =>
					R_next <= X"14";
					G_next <= X"27";
					B_next <= X"c1";
				when X"84" =>
					R_next <= X"25";
					G_next <= X"38";
					B_next <= X"d2";
				when X"85" =>
					R_next <= X"36";
					G_next <= X"49";
					B_next <= X"e3";
				when X"86" =>
					R_next <= X"47";
					G_next <= X"5a";
					B_next <= X"f4";
				when X"87" =>
					R_next <= X"58";
					G_next <= X"6b";
					B_next <= X"ff";
				when X"88" =>
					R_next <= X"69";
					G_next <= X"7c";
					B_next <= X"ff";
				when X"89" =>
					R_next <= X"7a";
					G_next <= X"8d";
					B_next <= X"ff";
				when X"8a" =>
					R_next <= X"8b";
					G_next <= X"9e";
					B_next <= X"ff";
				when X"8b" =>
					R_next <= X"9c";
					G_next <= X"af";
					B_next <= X"ff";
				when X"8c" =>
					R_next <= X"ad";
					G_next <= X"c0";
					B_next <= X"ff";
				when X"8d" =>
					R_next <= X"be";
					G_next <= X"d1";
					B_next <= X"ff";
				when X"8e" =>
					R_next <= X"cf";
					G_next <= X"e2";
					B_next <= X"ff";
				when X"8f" =>
					R_next <= X"e0";
					G_next <= X"f3";
					B_next <= X"ff";
				when X"90" =>
					R_next <= X"00";
					G_next <= X"0e";
					B_next <= X"64";
				when X"91" =>
					R_next <= X"00";
					G_next <= X"1f";
					B_next <= X"75";
				when X"92" =>
					R_next <= X"00";
					G_next <= X"30";
					B_next <= X"86";
				when X"93" =>
					R_next <= X"00";
					G_next <= X"41";
					B_next <= X"97";
				when X"94" =>
					R_next <= X"03";
					G_next <= X"52";
					B_next <= X"a8";
				when X"95" =>
					R_next <= X"14";
					G_next <= X"63";
					B_next <= X"b9";
				when X"96" =>
					R_next <= X"25";
					G_next <= X"74";
					B_next <= X"ca";
				when X"97" =>
					R_next <= X"36";
					G_next <= X"85";
					B_next <= X"db";
				when X"98" =>
					R_next <= X"47";
					G_next <= X"96";
					B_next <= X"ec";
				when X"99" =>
					R_next <= X"58";
					G_next <= X"a7";
					B_next <= X"fd";
				when X"9a" =>
					R_next <= X"69";
					G_next <= X"b8";
					B_next <= X"ff";
				when X"9b" =>
					R_next <= X"7a";
					G_next <= X"c9";
					B_next <= X"ff";
				when X"9c" =>
					R_next <= X"8b";
					G_next <= X"da";
					B_next <= X"ff";
				when X"9d" =>
					R_next <= X"9c";
					G_next <= X"eb";
					B_next <= X"ff";
				when X"9e" =>
					R_next <= X"ad";
					G_next <= X"fc";
					B_next <= X"ff";
				when X"9f" =>
					R_next <= X"be";
					G_next <= X"ff";
					B_next <= X"ff";
				when X"a0" =>
					R_next <= X"00";
					G_next <= X"24";
					B_next <= X"22";
				when X"a1" =>
					R_next <= X"00";
					G_next <= X"35";
					B_next <= X"33";
				when X"a2" =>
					R_next <= X"00";
					G_next <= X"46";
					B_next <= X"44";
				when X"a3" =>
					R_next <= X"00";
					G_next <= X"57";
					B_next <= X"55";
				when X"a4" =>
					R_next <= X"00";
					G_next <= X"68";
					B_next <= X"66";
				when X"a5" =>
					R_next <= X"02";
					G_next <= X"79";
					B_next <= X"77";
				when X"a6" =>
					R_next <= X"13";
					G_next <= X"8a";
					B_next <= X"88";
				when X"a7" =>
					R_next <= X"24";
					G_next <= X"9b";
					B_next <= X"99";
				when X"a8" =>
					R_next <= X"35";
					G_next <= X"ac";
					B_next <= X"aa";
				when X"a9" =>
					R_next <= X"46";
					G_next <= X"bd";
					B_next <= X"bb";
				when X"aa" =>
					R_next <= X"57";
					G_next <= X"ce";
					B_next <= X"cc";
				when X"ab" =>
					R_next <= X"68";
					G_next <= X"df";
					B_next <= X"dd";
				when X"ac" =>
					R_next <= X"79";
					G_next <= X"f0";
					B_next <= X"ee";
				when X"ad" =>
					R_next <= X"8a";
					G_next <= X"ff";
					B_next <= X"ff";
				when X"ae" =>
					R_next <= X"9b";
					G_next <= X"ff";
					B_next <= X"ff";
				when X"af" =>
					R_next <= X"ac";
					G_next <= X"ff";
					B_next <= X"ff";
				when X"b0" =>
					R_next <= X"00";
					G_next <= X"32";
					B_next <= X"00";
				when X"b1" =>
					R_next <= X"00";
					G_next <= X"43";
					B_next <= X"00";
				when X"b2" =>
					R_next <= X"00";
					G_next <= X"54";
					B_next <= X"00";
				when X"b3" =>
					R_next <= X"00";
					G_next <= X"65";
					B_next <= X"0c";
				when X"b4" =>
					R_next <= X"00";
					G_next <= X"76";
					B_next <= X"1d";
				when X"b5" =>
					R_next <= X"02";
					G_next <= X"87";
					B_next <= X"2e";
				when X"b6" =>
					R_next <= X"13";
					G_next <= X"98";
					B_next <= X"3f";
				when X"b7" =>
					R_next <= X"24";
					G_next <= X"a9";
					B_next <= X"50";
				when X"b8" =>
					R_next <= X"35";
					G_next <= X"ba";
					B_next <= X"61";
				when X"b9" =>
					R_next <= X"46";
					G_next <= X"cb";
					B_next <= X"72";
				when X"ba" =>
					R_next <= X"57";
					G_next <= X"dc";
					B_next <= X"83";
				when X"bb" =>
					R_next <= X"68";
					G_next <= X"ed";
					B_next <= X"94";
				when X"bc" =>
					R_next <= X"79";
					G_next <= X"fe";
					B_next <= X"a5";
				when X"bd" =>
					R_next <= X"8a";
					G_next <= X"ff";
					B_next <= X"b6";
				when X"be" =>
					R_next <= X"9b";
					G_next <= X"ff";
					B_next <= X"c7";
				when X"bf" =>
					R_next <= X"ac";
					G_next <= X"ff";
					B_next <= X"d8";
				when X"c0" =>
					R_next <= X"00";
					G_next <= X"34";
					B_next <= X"00";
				when X"c1" =>
					R_next <= X"00";
					G_next <= X"45";
					B_next <= X"00";
				when X"c2" =>
					R_next <= X"00";
					G_next <= X"56";
					B_next <= X"00";
				when X"c3" =>
					R_next <= X"00";
					G_next <= X"67";
					B_next <= X"00";
				when X"c4" =>
					R_next <= X"05";
					G_next <= X"78";
					B_next <= X"00";
				when X"c5" =>
					R_next <= X"16";
					G_next <= X"89";
					B_next <= X"00";
				when X"c6" =>
					R_next <= X"27";
					G_next <= X"9a";
					B_next <= X"00";
				when X"c7" =>
					R_next <= X"38";
					G_next <= X"ab";
					B_next <= X"0f";
				when X"c8" =>
					R_next <= X"49";
					G_next <= X"bc";
					B_next <= X"20";
				when X"c9" =>
					R_next <= X"5a";
					G_next <= X"cd";
					B_next <= X"31";
				when X"ca" =>
					R_next <= X"6b";
					G_next <= X"de";
					B_next <= X"42";
				when X"cb" =>
					R_next <= X"7c";
					G_next <= X"ef";
					B_next <= X"53";
				when X"cc" =>
					R_next <= X"8d";
					G_next <= X"ff";
					B_next <= X"64";
				when X"cd" =>
					R_next <= X"9e";
					G_next <= X"ff";
					B_next <= X"75";
				when X"ce" =>
					R_next <= X"af";
					G_next <= X"ff";
					B_next <= X"86";
				when X"cf" =>
					R_next <= X"c0";
					G_next <= X"ff";
					B_next <= X"97";
				when X"d0" =>
					R_next <= X"00";
					G_next <= X"2a";
					B_next <= X"00";
				when X"d1" =>
					R_next <= X"00";
					G_next <= X"3b";
					B_next <= X"00";
				when X"d2" =>
					R_next <= X"06";
					G_next <= X"4c";
					B_next <= X"00";
				when X"d3" =>
					R_next <= X"17";
					G_next <= X"5d";
					B_next <= X"00";
				when X"d4" =>
					R_next <= X"28";
					G_next <= X"6e";
					B_next <= X"00";
				when X"d5" =>
					R_next <= X"39";
					G_next <= X"7f";
					B_next <= X"00";
				when X"d6" =>
					R_next <= X"4a";
					G_next <= X"90";
					B_next <= X"00";
				when X"d7" =>
					R_next <= X"5b";
					G_next <= X"a1";
					B_next <= X"00";
				when X"d8" =>
					R_next <= X"6c";
					G_next <= X"b2";
					B_next <= X"00";
				when X"d9" =>
					R_next <= X"7d";
					G_next <= X"c3";
					B_next <= X"09";
				when X"da" =>
					R_next <= X"8e";
					G_next <= X"d4";
					B_next <= X"1a";
				when X"db" =>
					R_next <= X"9f";
					G_next <= X"e5";
					B_next <= X"2b";
				when X"dc" =>
					R_next <= X"b0";
					G_next <= X"f6";
					B_next <= X"3c";
				when X"dd" =>
					R_next <= X"c1";
					G_next <= X"ff";
					B_next <= X"4d";
				when X"de" =>
					R_next <= X"d2";
					G_next <= X"ff";
					B_next <= X"5e";
				when X"df" =>
					R_next <= X"e3";
					G_next <= X"ff";
					B_next <= X"6f";
				when X"e0" =>
					R_next <= X"0d";
					G_next <= X"17";
					B_next <= X"00";
				when X"e1" =>
					R_next <= X"1e";
					G_next <= X"28";
					B_next <= X"00";
				when X"e2" =>
					R_next <= X"2f";
					G_next <= X"39";
					B_next <= X"00";
				when X"e3" =>
					R_next <= X"40";
					G_next <= X"4a";
					B_next <= X"00";
				when X"e4" =>
					R_next <= X"51";
					G_next <= X"5b";
					B_next <= X"00";
				when X"e5" =>
					R_next <= X"62";
					G_next <= X"6c";
					B_next <= X"00";
				when X"e6" =>
					R_next <= X"73";
					G_next <= X"7d";
					B_next <= X"00";
				when X"e7" =>
					R_next <= X"84";
					G_next <= X"8e";
					B_next <= X"00";
				when X"e8" =>
					R_next <= X"95";
					G_next <= X"9f";
					B_next <= X"00";
				when X"e9" =>
					R_next <= X"a6";
					G_next <= X"b0";
					B_next <= X"02";
				when X"ea" =>
					R_next <= X"b7";
					G_next <= X"c1";
					B_next <= X"13";
				when X"eb" =>
					R_next <= X"c8";
					G_next <= X"d2";
					B_next <= X"24";
				when X"ec" =>
					R_next <= X"d9";
					G_next <= X"e3";
					B_next <= X"35";
				when X"ed" =>
					R_next <= X"ea";
					G_next <= X"f4";
					B_next <= X"46";
				when X"ee" =>
					R_next <= X"fb";
					G_next <= X"ff";
					B_next <= X"57";
				when X"ef" =>
					R_next <= X"ff";
					G_next <= X"ff";
					B_next <= X"68";
				when X"f0" =>
					R_next <= X"33";
					G_next <= X"00";
					B_next <= X"00";
				when X"f1" =>
					R_next <= X"44";
					G_next <= X"0f";
					B_next <= X"00";
				when X"f2" =>
					R_next <= X"55";
					G_next <= X"20";
					B_next <= X"00";
				when X"f3" =>
					R_next <= X"66";
					G_next <= X"31";
					B_next <= X"00";
				when X"f4" =>
					R_next <= X"77";
					G_next <= X"42";
					B_next <= X"00";
				when X"f5" =>
					R_next <= X"88";
					G_next <= X"53";
					B_next <= X"00";
				when X"f6" =>
					R_next <= X"99";
					G_next <= X"64";
					B_next <= X"00";
				when X"f7" =>
					R_next <= X"aa";
					G_next <= X"75";
					B_next <= X"00";
				when X"f8" =>
					R_next <= X"bb";
					G_next <= X"86";
					B_next <= X"0e";
				when X"f9" =>
					R_next <= X"cc";
					G_next <= X"97";
					B_next <= X"1f";
				when X"fa" =>
					R_next <= X"dd";
					G_next <= X"a8";
					B_next <= X"30";
				when X"fb" =>
					R_next <= X"ee";
					G_next <= X"b9";
					B_next <= X"41";
				when X"fc" =>
					R_next <= X"ff";
					G_next <= X"ca";
					B_next <= X"52";
				when X"fd" =>
					R_next <= X"ff";
					G_next <= X"db";
					B_next <= X"63";
				when X"fe" =>
					R_next <= X"ff";
					G_next <= X"ec";
					B_next <= X"74";
				when X"ff" =>
					R_next <= X"ff";
					G_next <= X"fd";
					B_next <= X"85";
				when others =>
					--nop
			end case;
		end if;
		end process;
end vhdl;
