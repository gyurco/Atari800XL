
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81ce",
X"bc738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81d5",
X"d40c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757581c8",
X"eb2d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7581c6ff",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80ddf304",
X"fd3d0d75",
X"705254ae",
X"a03f83c0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"c0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83c0",
X"8008732e",
X"a13883c0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183c0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83c2d008",
X"248a38b4",
X"f53fff0b",
X"83c2d00c",
X"800b83c0",
X"800c04ff",
X"3d0d7352",
X"83c0ac08",
X"722e8d38",
X"d93f7151",
X"96993f71",
X"83c0ac0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"558154bc",
X"15088191",
X"387451cf",
X"3f795880",
X"7a2580f7",
X"3883c380",
X"0870892a",
X"5783ff06",
X"78848072",
X"31565657",
X"73782583",
X"38735575",
X"83c2d008",
X"2e8438ff",
X"893f83c2",
X"d0088025",
X"a6387589",
X"2b5198dc",
X"3f83c380",
X"088f3dfc",
X"11555c54",
X"8152f81b",
X"5196c63f",
X"761483c3",
X"800c7583",
X"c2d00c74",
X"53765278",
X"51b3a63f",
X"83c08008",
X"83c38008",
X"1683c380",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8b3861",
X"7a710c54",
X"75547580",
X"2e833881",
X"547383c0",
X"800c8e3d",
X"0d04fc3d",
X"0dfe9b3f",
X"7651feaf",
X"3f863dfc",
X"05537852",
X"775195e9",
X"3f797571",
X"0c5483c0",
X"80085483",
X"c0800880",
X"2e833881",
X"547383c0",
X"800c863d",
X"0d04fe3d",
X"0d7583c2",
X"d0085353",
X"80722489",
X"3871732e",
X"8438fdd6",
X"3f7451fd",
X"ea3f7251",
X"97ae3f83",
X"c0800852",
X"83c08008",
X"802e8338",
X"81527183",
X"c0800c84",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"c0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"c0800c51",
X"823d0d04",
X"80c40b83",
X"c0800c04",
X"fd3d0d75",
X"77715470",
X"535553a9",
X"f83f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfceb3f",
X"735193ab",
X"3f7383c0",
X"ac0c83c0",
X"80085383",
X"c0800880",
X"2e833881",
X"537283c0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcbf3f",
X"72802ea5",
X"38bc1308",
X"527351a9",
X"823f83c0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"c0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83c0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83c2d0",
X"0c7483c0",
X"b00c7583",
X"c2cc0caf",
X"da3f83c0",
X"800881ff",
X"06528153",
X"71993883",
X"c2e8518e",
X"943f83c0",
X"80085283",
X"c0800880",
X"2e833872",
X"52715372",
X"83c0800c",
X"843d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"51a6f33f",
X"83c08008",
X"557483c0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"c0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283c2cc",
X"085181b5",
X"bc3f83c0",
X"800857f9",
X"e13f7952",
X"83c2d451",
X"95b73f83",
X"c0800854",
X"805383c0",
X"8008732e",
X"09810682",
X"833883c0",
X"b0080b0b",
X"81d3dc53",
X"705256a6",
X"b03f0b0b",
X"81d3dc52",
X"80c01651",
X"a6a33f75",
X"bc170c73",
X"82c0170c",
X"810b82c4",
X"170c810b",
X"82c8170c",
X"7382cc17",
X"0cff1782",
X"d0175557",
X"81913983",
X"c0bc3370",
X"822a7081",
X"06515455",
X"72818038",
X"74812a81",
X"06587780",
X"f6387484",
X"2a810682",
X"c4150c83",
X"c0bc3381",
X"0682c815",
X"0c795273",
X"51a5ca3f",
X"7351a5e1",
X"3f83c080",
X"081453af",
X"73708105",
X"553472bc",
X"150c83c0",
X"bd527251",
X"a5ab3f83",
X"c0b40882",
X"c0150c83",
X"c0ca5280",
X"c01451a5",
X"983f7880",
X"2e8d3873",
X"51782d83",
X"c0800880",
X"2e993877",
X"82cc150c",
X"75802e86",
X"387382cc",
X"170c7382",
X"d015ff19",
X"59555676",
X"802e9b38",
X"83c0b452",
X"83c2d451",
X"94ad3f83",
X"c080088a",
X"3883c0bd",
X"335372fe",
X"d2387880",
X"2e893883",
X"c0b00851",
X"fcb83f83",
X"c0b00853",
X"7283c080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb53f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f690",
X"3f83c080",
X"08745387",
X"3d705355",
X"55f6b03f",
X"f7903f73",
X"51d33f63",
X"53745283",
X"c0800851",
X"fab83f92",
X"3d0d0471",
X"83c0800c",
X"0480c012",
X"83c0800c",
X"04803d0d",
X"7282c011",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"c0800c51",
X"823d0d04",
X"f93d0d79",
X"83c09008",
X"57578177",
X"27819638",
X"76881708",
X"27818e38",
X"75335574",
X"822e8938",
X"74832eb3",
X"3880fe39",
X"74547610",
X"83fe0653",
X"76882a8c",
X"17080552",
X"893dfc05",
X"51aa883f",
X"83c08008",
X"80df3802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d13984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"51a9d83f",
X"83c08008",
X"b038029f",
X"05330284",
X"059e0533",
X"71982b71",
X"902b0702",
X"8c059d05",
X"3370882b",
X"72078d3d",
X"337180ff",
X"fffe8006",
X"07515253",
X"57585683",
X"39815574",
X"83c0800c",
X"893d0d04",
X"fb3d0d83",
X"c09008fe",
X"19881208",
X"fe055556",
X"54805674",
X"73278d38",
X"82143375",
X"71299416",
X"08055753",
X"7583c080",
X"0c873d0d",
X"04fc3d0d",
X"7652800b",
X"83c09008",
X"70335152",
X"5370832e",
X"09810691",
X"38951233",
X"94133371",
X"982b7190",
X"2b075555",
X"519b1233",
X"9a133371",
X"882b0774",
X"0783c080",
X"0c55863d",
X"0d04fc3d",
X"0d7683c0",
X"90085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"fed63f83",
X"c0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183c080",
X"0c863d0d",
X"04fa3d0d",
X"7883c090",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fcb13f",
X"81527183",
X"c0800827",
X"a8388352",
X"83c08008",
X"88170827",
X"9c3883c0",
X"80088c16",
X"0c83c080",
X"0851fdbc",
X"3f83c080",
X"0890160c",
X"73752380",
X"527183c0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585e5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"9f269138",
X"7a51fdd2",
X"3f83c080",
X"0856807d",
X"34838139",
X"933d841c",
X"08705859",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"3880705a",
X"5c887f08",
X"5f5a7b81",
X"1d7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535e57",
X"557480e7",
X"3876ae2e",
X"09810683",
X"38815578",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675bb",
X"3888598b",
X"5affab39",
X"76982b55",
X"74802587",
X"3881cdcc",
X"173357ff",
X"9f175574",
X"99268938",
X"e0177081",
X"ff065855",
X"78811a70",
X"81ff0672",
X"1b535b57",
X"55767534",
X"fef8397b",
X"1e7f0c80",
X"5576a026",
X"83388155",
X"748b1934",
X"7a51fc82",
X"3f83c080",
X"0880f538",
X"a0547a22",
X"70852b83",
X"e0065455",
X"901b0852",
X"7c51a493",
X"3f83c080",
X"085783c0",
X"80088181",
X"387c3355",
X"74802e80",
X"f4388b1d",
X"3370832a",
X"70810651",
X"565674b4",
X"388b7d84",
X"1d0883c0",
X"8008595b",
X"5b58ff18",
X"5877ff2e",
X"9a387970",
X"81055b33",
X"79708105",
X"5b337171",
X"31525656",
X"75802ee2",
X"38863975",
X"802e9638",
X"7a51fbe5",
X"3fff8639",
X"83c08008",
X"5683c080",
X"08b63883",
X"39765684",
X"1b088b11",
X"33515574",
X"a7388b1d",
X"3370842a",
X"70810651",
X"56567489",
X"38835694",
X"39815690",
X"397c51fa",
X"943f83c0",
X"8008881c",
X"0cfd8139",
X"7583c080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"51a2d83f",
X"835683c0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"51a2ac3f",
X"83c08008",
X"98388117",
X"33773371",
X"882b0783",
X"c0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"7651a283",
X"3f83c080",
X"08983881",
X"17337733",
X"71882b07",
X"83c08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583c080",
X"0c8a3d0d",
X"04eb3d0d",
X"675a800b",
X"83c0900c",
X"a1a53f83",
X"c0800881",
X"06558256",
X"7483ef38",
X"7475538f",
X"3d705357",
X"59feca3f",
X"83c08008",
X"81ff0657",
X"76812e09",
X"810680d4",
X"38905483",
X"be537452",
X"7551a197",
X"3f83c080",
X"0880c938",
X"8f3d3355",
X"74802e80",
X"c93802bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"33710770",
X"587b575e",
X"525e5759",
X"57fdee3f",
X"83c08008",
X"81ff0657",
X"76832e09",
X"81068638",
X"815682f2",
X"3976802e",
X"86388656",
X"82e839a4",
X"548d5378",
X"527551a0",
X"ae3f8156",
X"83c08008",
X"82d43802",
X"be053302",
X"8405bd05",
X"3371882b",
X"07595d77",
X"ab380280",
X"ce053302",
X"840580cd",
X"05337198",
X"2b71902b",
X"07973d33",
X"70882b72",
X"07029405",
X"80cb0533",
X"71075452",
X"5e575956",
X"02b70533",
X"78712902",
X"8805b605",
X"33028c05",
X"b5053371",
X"882b0770",
X"1d707f8c",
X"050c5f59",
X"57595d8e",
X"3d33821b",
X"3402b905",
X"33903d33",
X"71882b07",
X"5a5c7884",
X"1b2302bb",
X"05330284",
X"05ba0533",
X"71882b07",
X"565c74ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"07515253",
X"575e5c74",
X"76317831",
X"79842a90",
X"3d335471",
X"71315356",
X"5681a6a1",
X"3f83c080",
X"08820570",
X"881c0c83",
X"c08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83c0900c",
X"80567583",
X"c0800c97",
X"3d0d04e9",
X"3d0d83c0",
X"90085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e53f83c0",
X"80085483",
X"c0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f489",
X"3f83c080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383c080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83c09008",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0e93f",
X"83c08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"833f83c0",
X"80085583",
X"c0800880",
X"2eff8938",
X"83c08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"519ad43f",
X"83c08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83c0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83c09008",
X"55568555",
X"73802e81",
X"e3388114",
X"33810653",
X"84557280",
X"2e81d538",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b9388214",
X"3370892b",
X"56537680",
X"2eb73874",
X"52ff1651",
X"81a1a23f",
X"83c08008",
X"ff187654",
X"70535853",
X"81a1923f",
X"83c08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed63f83",
X"c0800853",
X"810b83c0",
X"8008278b",
X"38881408",
X"83c08008",
X"26883880",
X"0b811534",
X"b03983c0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc53f",
X"83c08008",
X"8c3883c0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683c0",
X"800805a8",
X"150c8055",
X"7483c080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83c09008",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1cf3f",
X"83c08008",
X"5583c080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef5",
X"3f83c080",
X"0888170c",
X"7551efa6",
X"3f83c080",
X"08557483",
X"c0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683c0",
X"9008802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f53f83c0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"96dd3f83",
X"c0800841",
X"83c08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"eddf3f83",
X"c0800841",
X"83c08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"8dff3f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f03f83c0",
X"80088332",
X"70307072",
X"079f2c83",
X"c0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"8c8b3f75",
X"83c0800c",
X"9e3d0d04",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"7751e0d2",
X"3f83c080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3381d5dc",
X"0b81d5dc",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"527751e0",
X"813f83c0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583c0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"558b923f",
X"83c08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"8114518a",
X"aa3f83c0",
X"80083070",
X"83c08008",
X"07802583",
X"c0800c53",
X"863d0d04",
X"fc3d0d76",
X"705255e6",
X"ee3f83c0",
X"80085481",
X"5383c080",
X"0880c138",
X"7451e6b1",
X"3f83c080",
X"0881d3ec",
X"5383c080",
X"085253ff",
X"913f83c0",
X"8008a138",
X"81d3f052",
X"7251ff82",
X"3f83c080",
X"08923881",
X"d3f45272",
X"51fef33f",
X"83c08008",
X"802e8338",
X"81547353",
X"7283c080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"e68d3f81",
X"5383c080",
X"08983873",
X"51e5d63f",
X"83c39808",
X"5283c080",
X"0851feba",
X"3f83c080",
X"08537283",
X"c0800c85",
X"3d0d04df",
X"3d0da43d",
X"0870525e",
X"dbfb3f83",
X"c0800833",
X"953d5654",
X"73963881",
X"d6f85274",
X"51898a3f",
X"9a397d52",
X"7851defc",
X"3f84cd39",
X"7d51dbe1",
X"3f83c080",
X"08527451",
X"db913f80",
X"43804280",
X"41804083",
X"c3a00852",
X"943d7052",
X"5de1e43f",
X"83c08008",
X"59800b83",
X"c0800855",
X"5b83c080",
X"087b2e94",
X"38811b74",
X"525be4e6",
X"3f83c080",
X"085483c0",
X"8008ee38",
X"805aff5f",
X"7909709f",
X"2c7b065b",
X"547a7a24",
X"8438ff1b",
X"5af61a70",
X"09709f2c",
X"72067bff",
X"125a5a52",
X"55558075",
X"25953876",
X"51e4ab3f",
X"83c08008",
X"76ff1858",
X"55577380",
X"24ed3874",
X"7f2e8638",
X"a0cf3f74",
X"5f78ff1b",
X"70585d58",
X"807a2595",
X"387751e4",
X"813f83c0",
X"800876ff",
X"18585558",
X"738024ed",
X"38800b83",
X"c7d00c80",
X"0b83c884",
X"0c81d3f8",
X"518d8d3f",
X"81800b83",
X"c8840c81",
X"d480518c",
X"ff3fa80b",
X"83c7d00c",
X"76802e80",
X"e43883c7",
X"d0087779",
X"32703070",
X"72078025",
X"70872b83",
X"c8840c51",
X"56785356",
X"56e3b83f",
X"83c08008",
X"802e8838",
X"81d48851",
X"8cc63f76",
X"51e2fa3f",
X"83c08008",
X"5281d59c",
X"518cb53f",
X"7651e382",
X"3f83c080",
X"0883c7d0",
X"08555775",
X"74258638",
X"a81656f7",
X"397583c7",
X"d00c86f0",
X"7624ff98",
X"3887980b",
X"83c7d00c",
X"77802eb1",
X"387751e2",
X"b83f83c0",
X"80087852",
X"55e2d83f",
X"81d49054",
X"83c08008",
X"8d388739",
X"80763481",
X"ce3981d4",
X"8c547453",
X"735281d3",
X"e0518bd4",
X"3f805481",
X"d3e8518b",
X"cb3f8114",
X"5473a82e",
X"098106ef",
X"38868da0",
X"519cc33f",
X"8052903d",
X"705257b1",
X"a53f8352",
X"7651b19e",
X"3f62818f",
X"3861802e",
X"80fb387b",
X"5473ff2e",
X"96387880",
X"2e818938",
X"7851e1de",
X"3f83c080",
X"08ff1555",
X"59e73978",
X"802e80f4",
X"387851e1",
X"da3f83c0",
X"8008802e",
X"fc903878",
X"51e1a23f",
X"83c08008",
X"5281d3dc",
X"5183df3f",
X"83c08008",
X"a3387c51",
X"85973f83",
X"c0800855",
X"74ff1656",
X"54807425",
X"ae38741d",
X"70335556",
X"73af2efe",
X"cf38e939",
X"7851e0e3",
X"3f83c080",
X"08527c51",
X"84cf3f8f",
X"397f8829",
X"6010057a",
X"0561055a",
X"fc923962",
X"802efbd3",
X"38805276",
X"51afff3f",
X"a33d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"842a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"a80b9088",
X"b834b80b",
X"9088b834",
X"7083c080",
X"0c823d0d",
X"04803d0d",
X"9088b833",
X"7081ff06",
X"70852a81",
X"32708106",
X"51515151",
X"70802e8d",
X"38980b90",
X"88b834b8",
X"0b9088b8",
X"347083c0",
X"800c823d",
X"0d04930b",
X"9088bc34",
X"ff0b9088",
X"a83404ff",
X"3d0d028f",
X"05335280",
X"0b9088bc",
X"348a519a",
X"8d3fdf3f",
X"80f80b90",
X"88a03480",
X"0b908888",
X"34fa1252",
X"71908880",
X"34800b90",
X"88983471",
X"90889034",
X"9088b852",
X"807234b8",
X"7234833d",
X"0d04803d",
X"0d028b05",
X"33517090",
X"88b434fe",
X"bf3f83c0",
X"8008802e",
X"f638823d",
X"0d04803d",
X"0d8439a7",
X"a63ffed9",
X"3f83c080",
X"08802ef3",
X"389088b4",
X"337081ff",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0da30b90",
X"88bc34ff",
X"0b9088a8",
X"349088b8",
X"51a87134",
X"b8713482",
X"3d0d0480",
X"3d0d9088",
X"bc337098",
X"2b708025",
X"83c0800c",
X"5151823d",
X"0d04803d",
X"0d9088b8",
X"337081ff",
X"0670832a",
X"81327081",
X"06515151",
X"5170802e",
X"e838b00b",
X"9088b834",
X"b80b9088",
X"b834823d",
X"0d04803d",
X"0d9080ac",
X"08810683",
X"c0800c82",
X"3d0d04fd",
X"3d0d7577",
X"54548073",
X"25943873",
X"70810555",
X"335281d4",
X"94518788",
X"3fff1353",
X"e939853d",
X"0d04fd3d",
X"0d757753",
X"54733351",
X"70893871",
X"33517080",
X"2ea13873",
X"33723352",
X"53727127",
X"8538ff51",
X"94397073",
X"27853881",
X"518b3981",
X"14811353",
X"54d33980",
X"517083c0",
X"800c853d",
X"0d04fd3d",
X"0d757754",
X"54723370",
X"81ff0652",
X"5270802e",
X"a3387181",
X"ff068114",
X"ffbf1253",
X"54527099",
X"268938a0",
X"127081ff",
X"06535171",
X"74708105",
X"5634d239",
X"80743485",
X"3d0d04ff",
X"bd3d0d80",
X"c63d0852",
X"a53d7052",
X"54ffb33f",
X"80c73d08",
X"52853d70",
X"5253ffa6",
X"3f725273",
X"51fedf3f",
X"80c53d0d",
X"04fe3d0d",
X"74765353",
X"71708105",
X"53335170",
X"73708105",
X"553470f0",
X"38843d0d",
X"04fe3d0d",
X"74528072",
X"33525370",
X"732e8d38",
X"81128114",
X"71335354",
X"5270f538",
X"7283c080",
X"0c843d0d",
X"04f63d0d",
X"7c7e6062",
X"5a5d5b56",
X"80598155",
X"8539747a",
X"29557452",
X"7551818d",
X"fc3f83c0",
X"80087a27",
X"ed387480",
X"2e80e038",
X"74527551",
X"818de63f",
X"83c08008",
X"75537652",
X"54818e8c",
X"3f83c080",
X"087a5375",
X"5256818d",
X"cc3f83c0",
X"80087930",
X"707b079f",
X"2a707780",
X"24075151",
X"54557287",
X"3883c080",
X"08c23876",
X"8118b016",
X"55585889",
X"74258b38",
X"b714537a",
X"853880d7",
X"14537278",
X"34811959",
X"ff9c3980",
X"77348c3d",
X"0d04f73d",
X"0d7b7d7f",
X"62029005",
X"bb053357",
X"59565a5a",
X"b0587283",
X"38a05875",
X"70708105",
X"52337159",
X"54559039",
X"8074258e",
X"38ff1477",
X"70810559",
X"33545472",
X"ef3873ff",
X"15555380",
X"73258938",
X"77527951",
X"782def39",
X"75337557",
X"5372802e",
X"90387252",
X"7951782d",
X"75708105",
X"573353ed",
X"398b3d0d",
X"04ee3d0d",
X"64666969",
X"70708105",
X"52335b4a",
X"5c5e5e76",
X"802e82f9",
X"3876a52e",
X"09810682",
X"e0388070",
X"41677070",
X"81055233",
X"714a5957",
X"5f76b02e",
X"0981068c",
X"38757081",
X"05573376",
X"4857815f",
X"d0175675",
X"892680da",
X"3876675c",
X"59805c93",
X"39778a24",
X"80c3387b",
X"8a29187b",
X"7081055d",
X"335a5cd0",
X"197081ff",
X"06585889",
X"7727a438",
X"ff9f1970",
X"81ff06ff",
X"a91b5a51",
X"56857627",
X"9238ffbf",
X"197081ff",
X"06515675",
X"85268a38",
X"c9195877",
X"8025ffb9",
X"387a477b",
X"407881ff",
X"06577680",
X"e42e80e5",
X"387680e4",
X"24a73876",
X"80d82e81",
X"86387680",
X"d8249038",
X"76802e81",
X"cc3876a5",
X"2e81b638",
X"81b93976",
X"80e32e81",
X"8c3881af",
X"397680f5",
X"2e9b3876",
X"80f5248b",
X"387680f3",
X"2e818138",
X"81993976",
X"80f82e80",
X"ca38818f",
X"39913d70",
X"55578053",
X"8a527984",
X"1b710853",
X"5b56fbfd",
X"3f7655ab",
X"3979841b",
X"7108943d",
X"705b5b52",
X"5b567580",
X"258c3875",
X"3056ad78",
X"340280c1",
X"05577654",
X"80538a52",
X"7551fbd1",
X"3f77557e",
X"54b83991",
X"3d705577",
X"80d83270",
X"30708025",
X"56515856",
X"90527984",
X"1b710853",
X"5b57fbad",
X"3f7555db",
X"3979841b",
X"83123354",
X"5b569839",
X"79841b71",
X"08575b56",
X"80547f53",
X"7c527d51",
X"fc9c3f87",
X"3976527d",
X"517c2d66",
X"70335881",
X"0547fd83",
X"39943d0d",
X"047283c0",
X"940c7183",
X"c0980c04",
X"fb3d0d88",
X"3d707084",
X"05520857",
X"54755383",
X"c0940852",
X"83c09808",
X"51fcc63f",
X"873d0d04",
X"ff3d0d73",
X"70085351",
X"02930533",
X"72347008",
X"8105710c",
X"833d0d04",
X"fc3d0d87",
X"3d881155",
X"7854bdb8",
X"5351fc99",
X"3f805287",
X"3d51d13f",
X"863d0d04",
X"fc3d0d76",
X"557483c3",
X"ac082eaf",
X"38805374",
X"5187c13f",
X"83c08008",
X"81ff06ff",
X"147081ff",
X"06723070",
X"9f2a5152",
X"55535472",
X"802e8438",
X"71dd3873",
X"fe387483",
X"c3ac0c86",
X"3d0d04ff",
X"3d0dff0b",
X"83c3ac0c",
X"84a53f81",
X"5187853f",
X"83c08008",
X"81ff0652",
X"71ee3881",
X"d33f7183",
X"c0800c83",
X"3d0d04fc",
X"3d0d7602",
X"8405a205",
X"22028805",
X"a605227a",
X"54555555",
X"ff823f72",
X"802ea038",
X"83c3c014",
X"33757081",
X"05573481",
X"147083ff",
X"ff06ff15",
X"7083ffff",
X"06565255",
X"52dd3980",
X"0b83c080",
X"0c863d0d",
X"04fc3d0d",
X"76787a11",
X"56535580",
X"5371742e",
X"93387215",
X"51703383",
X"c3c01334",
X"81128114",
X"5452ea39",
X"800b83c0",
X"800c863d",
X"0d04fd3d",
X"0d905483",
X"c3ac0851",
X"86f43f83",
X"c0800881",
X"ff06ff15",
X"71307130",
X"7073079f",
X"2a729f2a",
X"06525552",
X"555372db",
X"38853d0d",
X"04803d0d",
X"83c3b808",
X"1083c3b0",
X"08079080",
X"a80c823d",
X"0d04800b",
X"83c3b80c",
X"e43f0481",
X"0b83c3b8",
X"0cdb3f04",
X"ed3f0471",
X"83c3b40c",
X"04803d0d",
X"8051f43f",
X"810b83c3",
X"b80c810b",
X"83c3b00c",
X"ffbb3f82",
X"3d0d0480",
X"3d0d7230",
X"70740780",
X"2583c3b0",
X"0c51ffa5",
X"3f823d0d",
X"04803d0d",
X"028b0533",
X"9080a40c",
X"9080a808",
X"70810651",
X"5170f538",
X"9080a408",
X"7081ff06",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"81ff51d1",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"823d0d04",
X"803d0d73",
X"902b7307",
X"9080b40c",
X"823d0d04",
X"04fb3d0d",
X"78028405",
X"9f053370",
X"982b5557",
X"55728025",
X"9b387580",
X"ff065680",
X"5280f751",
X"e03f83c0",
X"800881ff",
X"06547381",
X"2680ff38",
X"8051fee7",
X"3fffa23f",
X"8151fedf",
X"3fff9a3f",
X"7551feed",
X"3f74982a",
X"51fee63f",
X"74902a70",
X"81ff0652",
X"53feda3f",
X"74882a70",
X"81ff0652",
X"53fece3f",
X"7481ff06",
X"51fec63f",
X"81557580",
X"c02e0981",
X"06863881",
X"95558d39",
X"7580c82e",
X"09810684",
X"38818755",
X"7451fea5",
X"3f8a55fe",
X"c83f83c0",
X"800881ff",
X"0670982b",
X"54547280",
X"258c38ff",
X"157081ff",
X"06565374",
X"e2387383",
X"c0800c87",
X"3d0d04fa",
X"3d0dfdc5",
X"3f8051fd",
X"da3f8a54",
X"fe933fff",
X"147081ff",
X"06555373",
X"f3387374",
X"535580c0",
X"51fea63f",
X"83c08008",
X"81ff0654",
X"73812e09",
X"8106829f",
X"3883aa52",
X"80c851fe",
X"8c3f83c0",
X"800881ff",
X"06537281",
X"2e098106",
X"81a83874",
X"54873d74",
X"115456fd",
X"c83f83c0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e5",
X"38029a05",
X"33537281",
X"2e098106",
X"81d93802",
X"9b053353",
X"80ce9054",
X"7281aa2e",
X"8d3881c7",
X"3980e451",
X"8ab43fff",
X"14547380",
X"2e81b838",
X"820a5281",
X"e951fda5",
X"3f83c080",
X"0881ff06",
X"5372de38",
X"725280fa",
X"51fd923f",
X"83c08008",
X"81ff0653",
X"72819038",
X"72547316",
X"53fcd63f",
X"83c08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e83887",
X"3d337086",
X"2a708106",
X"5154548c",
X"557280e3",
X"38845580",
X"de397452",
X"81e951fc",
X"cc3f83c0",
X"800881ff",
X"06538255",
X"81e95681",
X"73278638",
X"735580c1",
X"5680ce90",
X"548a3980",
X"e45189a6",
X"3fff1454",
X"73802ea9",
X"38805275",
X"51fc9a3f",
X"83c08008",
X"81ff0653",
X"72e13884",
X"805280d0",
X"51fc863f",
X"83c08008",
X"81ff0653",
X"72802e83",
X"38805574",
X"83c3bc34",
X"8051fb87",
X"3ffbc23f",
X"883d0d04",
X"fb3d0d77",
X"54800b83",
X"c3bc3370",
X"832a7081",
X"06515557",
X"5572752e",
X"09810685",
X"3873892b",
X"54735280",
X"d151fbbd",
X"3f83c080",
X"0881ff06",
X"5372bd38",
X"82b8c054",
X"fb833f83",
X"c0800881",
X"ff065372",
X"81ff2e09",
X"81068938",
X"ff145473",
X"e7389f39",
X"7281fe2e",
X"09810696",
X"3883c7c0",
X"5283c3c0",
X"51faed3f",
X"fad33ffa",
X"d03f8339",
X"81558051",
X"fa893ffa",
X"c43f7481",
X"ff0683c0",
X"800c873d",
X"0d04fb3d",
X"0d7783c3",
X"c0565481",
X"51f9ec3f",
X"83c3bc33",
X"70832a70",
X"81065154",
X"56728538",
X"73892b54",
X"735280d8",
X"51fab63f",
X"83c08008",
X"81ff0653",
X"7280e438",
X"81ff51f9",
X"d43f81fe",
X"51f9ce3f",
X"84805374",
X"70810556",
X"3351f9c1",
X"3fff1370",
X"83ffff06",
X"515372eb",
X"387251f9",
X"b03f7251",
X"f9ab3ff9",
X"d03f83c0",
X"80089f06",
X"53a78854",
X"72852e8c",
X"38993980",
X"e45186de",
X"3fff1454",
X"f9b33f83",
X"c0800881",
X"ff2e8438",
X"73e93880",
X"51f8e43f",
X"f99f3f80",
X"0b83c080",
X"0c873d0d",
X"047183c7",
X"c40c8880",
X"800b83c7",
X"c00c8480",
X"800b83c7",
X"c80c04f0",
X"3d0d8380",
X"805683c7",
X"c4081683",
X"c7c00817",
X"56547433",
X"743483c7",
X"c8081654",
X"80743481",
X"16567583",
X"80a02e09",
X"8106db38",
X"83d08056",
X"83c7c408",
X"1683c7c0",
X"08175654",
X"74337434",
X"83c7c808",
X"16548074",
X"34811656",
X"7583d090",
X"2e098106",
X"db3883a8",
X"805683c7",
X"c4081683",
X"c7c00817",
X"56547433",
X"743483c7",
X"c8081654",
X"80743481",
X"16567583",
X"a8902e09",
X"8106db38",
X"805683c7",
X"c4081683",
X"c7c80817",
X"55557333",
X"75348116",
X"56758180",
X"802e0981",
X"06e43887",
X"843f893d",
X"58a25381",
X"cfcc5277",
X"518183f0",
X"3f80578c",
X"805683c7",
X"c8081677",
X"19555573",
X"33753481",
X"16811858",
X"5676a22e",
X"098106e6",
X"38860b87",
X"a8833480",
X"0b87a882",
X"34800b87",
X"809a34af",
X"0b878096",
X"34bf0b87",
X"80973480",
X"0b878098",
X"349f0b87",
X"80993480",
X"0b87809b",
X"34f80b87",
X"a8893476",
X"87a88034",
X"820b87d0",
X"8f34820b",
X"87a88134",
X"840b8780",
X"9f34ff0b",
X"87d08b34",
X"923d0d04",
X"fe3d0d80",
X"5383c7c8",
X"081383c7",
X"c4081452",
X"52703372",
X"34811353",
X"72818080",
X"2e098106",
X"e4388380",
X"805383c7",
X"c8081383",
X"c7c40814",
X"52527033",
X"72348113",
X"53728380",
X"a02e0981",
X"06e43883",
X"d0805383",
X"c7c80813",
X"83c7c408",
X"14525270",
X"33723481",
X"13537283",
X"d0902e09",
X"8106e438",
X"83a88053",
X"83c7c808",
X"1383c7c4",
X"08145252",
X"70337234",
X"81135372",
X"83a8902e",
X"098106e4",
X"38843d0d",
X"04803d0d",
X"90809008",
X"810683c0",
X"800c823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087081",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fd0676",
X"1007720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870822c",
X"bf0683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe830676",
X"822b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087088",
X"2c870683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f1ff06",
X"76882b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"912cbf06",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fc87",
X"ffff0676",
X"912b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087099",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70ffbf0a",
X"0676992b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90808008",
X"70882c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"0870892c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708a",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8b2c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708c2cbf",
X"0683c080",
X"0c51823d",
X"0d04fe3d",
X"0d7481e6",
X"29872a90",
X"80a00c84",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70810554",
X"34ff1151",
X"f039843d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"8405540c",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"81808053",
X"80528880",
X"0a51ffb3",
X"3fa08053",
X"80528280",
X"0a51c73f",
X"843d0d04",
X"803d0d81",
X"51fcab3f",
X"72802e90",
X"388051fd",
X"ff3fce3f",
X"81d6d033",
X"51fdf53f",
X"8151fcbc",
X"3f8051fc",
X"b73f8051",
X"fc883f82",
X"3d0d04fd",
X"3d0d7552",
X"805480ff",
X"72258838",
X"810bff80",
X"135354ff",
X"bf125170",
X"99268638",
X"e01252b0",
X"39ff9f12",
X"51997127",
X"a738d012",
X"e0135451",
X"70892685",
X"38725298",
X"39728f26",
X"85387252",
X"8f3971ba",
X"2e098106",
X"85389a52",
X"83398052",
X"73802e85",
X"38818012",
X"527181ff",
X"0683c080",
X"0c853d0d",
X"04803d0d",
X"84d8c051",
X"80717081",
X"05533470",
X"84e0c02e",
X"098106f0",
X"38823d0d",
X"04fe3d0d",
X"02970533",
X"51fef43f",
X"83c08008",
X"81ff0683",
X"c7d00854",
X"52807324",
X"9b3883c8",
X"80081372",
X"83c88408",
X"07535371",
X"733483c7",
X"d0088105",
X"83c7d00c",
X"843d0d04",
X"fa3d0d82",
X"800a1b55",
X"8057883d",
X"fc055479",
X"53745278",
X"51ffbb92",
X"3f883d0d",
X"04fe3d0d",
X"83c7e808",
X"527451c1",
X"f63f83c0",
X"80088c38",
X"76537552",
X"83c7e808",
X"51c63f84",
X"3d0d04fe",
X"3d0d83c7",
X"e8085375",
X"527451ff",
X"bcb43f83",
X"c080088d",
X"38775376",
X"5283c7e8",
X"0851ffa0",
X"3f843d0d",
X"04fd3d0d",
X"83c7e808",
X"51ffbba7",
X"3f83c080",
X"0890802e",
X"098106ad",
X"38805483",
X"c1808053",
X"83c08008",
X"5283c7e8",
X"0851fef0",
X"3f87c180",
X"80143387",
X"c1908015",
X"34811454",
X"7390802e",
X"098106e9",
X"38853d0d",
X"0481d49c",
X"0b83c080",
X"0c04fc3d",
X"0d765473",
X"902e80ff",
X"38739024",
X"8e387384",
X"2e983873",
X"862ea638",
X"82b93973",
X"932e8195",
X"3873942e",
X"81cf3882",
X"aa398180",
X"80538280",
X"805283c7",
X"e40851fe",
X"8f3f82b5",
X"39805481",
X"80805380",
X"c0805283",
X"c7e40851",
X"fdfa3f82",
X"80805380",
X"c0805283",
X"c7e40851",
X"fdea3f84",
X"81808014",
X"338481c0",
X"80153484",
X"82808014",
X"338482c0",
X"80153481",
X"14547380",
X"c0802e09",
X"8106dc38",
X"81eb3982",
X"80805381",
X"80805283",
X"c7e40851",
X"fdb23f80",
X"54848280",
X"80143384",
X"81808015",
X"34811454",
X"73818080",
X"2e098106",
X"e83881bd",
X"39818080",
X"5380c080",
X"5283c7e4",
X"0851fd84",
X"3f805584",
X"81808015",
X"54733384",
X"81c08016",
X"34733384",
X"82808016",
X"34733384",
X"82c08016",
X"34811555",
X"7480c080",
X"2e098106",
X"d63880fd",
X"39818080",
X"53a08052",
X"83c7e408",
X"51fcc53f",
X"80558481",
X"80801554",
X"73338481",
X"a0801634",
X"73338481",
X"c0801634",
X"73338481",
X"e0801634",
X"73338482",
X"80801634",
X"73338482",
X"a0801634",
X"73338482",
X"c0801634",
X"73338482",
X"e0801634",
X"81155574",
X"a0802e09",
X"8106ffb6",
X"389f39fb",
X"9c3f800b",
X"83c7d00c",
X"800b83c8",
X"840c81d4",
X"a051e7fc",
X"3f81b78d",
X"c051f8fe",
X"3f863d0d",
X"04fc3d0d",
X"76705255",
X"ffbec83f",
X"83c08008",
X"54815383",
X"c0800880",
X"c2387451",
X"ffbe8a3f",
X"83c08008",
X"81d4bc53",
X"83c08008",
X"5253d6ea",
X"3f83c080",
X"08a13881",
X"d4c05272",
X"51d6db3f",
X"83c08008",
X"923881d4",
X"c4527251",
X"d6cc3f83",
X"c0800880",
X"2e833881",
X"54735372",
X"83c0800c",
X"863d0d04",
X"f13d0d80",
X"d5a90b83",
X"c3a00c83",
X"c7e40851",
X"d7f93f83",
X"c7e40851",
X"ffb3f63f",
X"ff0b81d4",
X"c05383c0",
X"80085256",
X"d68c3f83",
X"c0800880",
X"2e9f3880",
X"58913ddc",
X"11555590",
X"53f01552",
X"83c7e408",
X"51ffb5d2",
X"3f02b705",
X"335681a5",
X"3983c7e4",
X"0851ffb6",
X"ae3f83c0",
X"80085783",
X"c0800882",
X"80802e09",
X"81068338",
X"845683c0",
X"80088180",
X"802e0981",
X"0680e138",
X"805c805b",
X"805a8059",
X"f9933f80",
X"0b83c7d0",
X"0c800b83",
X"c8840c81",
X"d4c851e5",
X"f33f80d0",
X"0b83c7d0",
X"0c81d4d8",
X"51e5e53f",
X"80f80b83",
X"c7d00c81",
X"d4ec51e5",
X"d73f7580",
X"25a23880",
X"52893d70",
X"52558bbe",
X"3f835274",
X"518bb73f",
X"78557480",
X"25833890",
X"56807525",
X"dd388656",
X"7680c080",
X"2e098106",
X"85389356",
X"8c3976a0",
X"802e0981",
X"06833894",
X"567551fa",
X"ad3f913d",
X"0d04f73d",
X"0d805a80",
X"59805880",
X"57807056",
X"56f88a3f",
X"800b83c7",
X"d00c800b",
X"83c8840c",
X"81d58051",
X"e4ea3f81",
X"800b83c8",
X"840c81d5",
X"8451e4dc",
X"3f80d00b",
X"83c7d00c",
X"74307076",
X"07802570",
X"872b83c8",
X"840c5153",
X"f3ac3f83",
X"c0800852",
X"81d58c51",
X"e4b63f80",
X"f80b83c7",
X"d00c7481",
X"32703070",
X"72078025",
X"70872b83",
X"c8840c51",
X"5454f9a9",
X"3f83c080",
X"085281d5",
X"9851e48c",
X"3f81a00b",
X"83c7d00c",
X"74823270",
X"30707207",
X"80257087",
X"2b83c884",
X"0c515483",
X"c7e80852",
X"54ffb0ed",
X"3f83c080",
X"085281d5",
X"a051e3dc",
X"3f81c80b",
X"83c7d00c",
X"74833270",
X"30707207",
X"80257087",
X"2b83c884",
X"0c515483",
X"c7e40852",
X"54ffb0bd",
X"3f81d5a8",
X"5383c080",
X"08802e8f",
X"3883c7e4",
X"0851ffb0",
X"a83f83c0",
X"80085372",
X"5281d5b0",
X"51e3953f",
X"81f00b83",
X"c7d00c74",
X"84327030",
X"70720780",
X"2570872b",
X"83c8840c",
X"515581d5",
X"b85253e2",
X"f33f868d",
X"a051f3f6",
X"3f805287",
X"3d705253",
X"88d83f83",
X"52725188",
X"d13f7953",
X"7281c138",
X"77155574",
X"80258538",
X"72559039",
X"84752585",
X"38845587",
X"39748426",
X"81a03874",
X"842981cf",
X"f0055372",
X"0804f196",
X"3f83c080",
X"08775553",
X"73812e09",
X"81068938",
X"83c08008",
X"10539039",
X"73ff2e09",
X"81068838",
X"83c08008",
X"812c5390",
X"73258538",
X"90538839",
X"72802483",
X"38815372",
X"51f0f03f",
X"80d439f1",
X"823f83c0",
X"80081753",
X"72802585",
X"38805388",
X"39877325",
X"83388753",
X"7251f0fc",
X"3fb43976",
X"86387880",
X"2eac3883",
X"c39c0883",
X"c3980cad",
X"e50b83c3",
X"a00c83c7",
X"e80851d2",
X"ae3ff5f5",
X"3f903978",
X"802e8b38",
X"fa963f81",
X"538c3978",
X"87387580",
X"2efc9638",
X"80537283",
X"c0800c8b",
X"3d0d04ff",
X"3d0d83c7",
X"f05180e2",
X"eb3ff19d",
X"3f83c080",
X"08802e86",
X"38805180",
X"da39f1a2",
X"3f83c080",
X"0880ce38",
X"f1c23f83",
X"c0800880",
X"2eaa3881",
X"51eeff3f",
X"ebb93f80",
X"0b83c7d0",
X"0cfbbb3f",
X"83c08008",
X"52ff0b83",
X"c7d00ced",
X"cb3f71a1",
X"387151ee",
X"dd3f9f39",
X"f0f93f83",
X"c0800880",
X"2e943881",
X"51eecb3f",
X"eb853ff9",
X"8f3feda8",
X"3f8151f2",
X"8b3f833d",
X"0d04fe3d",
X"0d805283",
X"c7f05180",
X"d2aa3f82",
X"80805380",
X"52818180",
X"8051f18f",
X"3f80c080",
X"53805284",
X"81808051",
X"f1a03f90",
X"80805286",
X"84808051",
X"ffb0fd3f",
X"83c08008",
X"a43881d6",
X"e051ffb5",
X"c03f83c7",
X"e8085381",
X"d5c05283",
X"c0800851",
X"ffb09f3f",
X"83c08008",
X"8438f3f9",
X"3f8151f1",
X"a33ffe9f",
X"3ffc3983",
X"c08c0802",
X"83c08c0c",
X"fb3d0d02",
X"81d5cc0b",
X"83c39c0c",
X"81d4c40b",
X"83c3940c",
X"81d4c00b",
X"83c3a80c",
X"81d5d00b",
X"83c3a40c",
X"83c08c08",
X"fc050c80",
X"0b83c7d4",
X"0b83c08c",
X"08f8050c",
X"83c08c08",
X"f4050cff",
X"aef63f83",
X"c0800886",
X"05fc0683",
X"c08c08f0",
X"050c0283",
X"c08c08f0",
X"0508310d",
X"833d7083",
X"c08c08f8",
X"05087084",
X"0583c08c",
X"08f8050c",
X"0c51ffab",
X"be3f83c0",
X"8c08f405",
X"08810583",
X"c08c08f4",
X"050c83c0",
X"8c08f405",
X"08872e09",
X"8106ffab",
X"38869480",
X"8051e8d1",
X"3fff0b83",
X"c7d00c80",
X"0b83c884",
X"0c84d8c0",
X"0b83c880",
X"0c8151ec",
X"913f8151",
X"ecb63f80",
X"51ecb13f",
X"8151ecd7",
X"3f8251ec",
X"ff3f8051",
X"eda73f80",
X"51edd13f",
X"80d0c152",
X"8051ddb5",
X"3ffdaf3f",
X"83c08c08",
X"fc05080d",
X"800b83c0",
X"800c873d",
X"0d83c08c",
X"0c04fa3d",
X"0d785580",
X"750c800b",
X"84160c80",
X"0b88160c",
X"83c7f051",
X"80def93f",
X"edff3f83",
X"c0800887",
X"d0883370",
X"81ff0651",
X"535671a7",
X"3887d080",
X"3383c894",
X"3487d081",
X"3383c890",
X"3487d082",
X"3383c888",
X"3487d083",
X"3383c88c",
X"34ff0b87",
X"d08b3487",
X"d0893387",
X"d08f3370",
X"822a7081",
X"06703070",
X"72077009",
X"709f2c77",
X"069e0657",
X"51515651",
X"51545480",
X"74980653",
X"5371882e",
X"09810683",
X"38815371",
X"98327030",
X"70802575",
X"71318419",
X"0c515152",
X"80748606",
X"53537182",
X"2e098106",
X"83388153",
X"71863270",
X"30708025",
X"75713178",
X"0c515152",
X"83c89433",
X"5281aa72",
X"27843881",
X"750c83c8",
X"94335271",
X"bb268438",
X"ff750c83",
X"c8903352",
X"81aa7227",
X"8638810b",
X"84160c83",
X"c8903352",
X"71bb2686",
X"38ff0b84",
X"160c83c8",
X"88335281",
X"aa722784",
X"3881750c",
X"83c88833",
X"5271bb26",
X"8438ff75",
X"0c83c88c",
X"335281aa",
X"72278638",
X"810b8416",
X"0c83c88c",
X"335271bb",
X"268638ff",
X"0b84160c",
X"80577394",
X"2eaa3887",
X"80903387",
X"80913387",
X"80923370",
X"81ff0672",
X"74060687",
X"80933371",
X"06810651",
X"52545454",
X"72772e09",
X"81068338",
X"81577688",
X"160c7580",
X"2eb03875",
X"812a7081",
X"06778106",
X"3184170c",
X"5275832a",
X"76822a71",
X"81067181",
X"0631770c",
X"53537584",
X"2a810688",
X"160c7585",
X"2a81068c",
X"160c883d",
X"0d04fe3d",
X"0d747654",
X"527151fc",
X"d93f7281",
X"2ea23881",
X"73268d38",
X"72822ea8",
X"3872832e",
X"9c38e639",
X"7108e238",
X"841208dd",
X"38881208",
X"d838a539",
X"88120881",
X"2e9e3891",
X"39881208",
X"812e9538",
X"71089138",
X"8412088c",
X"388c1208",
X"812e0981",
X"06ffb238",
X"843d0d04",
X"fb3d0d78",
X"0284059f",
X"05335556",
X"800b81d1",
X"f0565381",
X"732b7406",
X"5271802e",
X"83388152",
X"74708205",
X"56227073",
X"902b0790",
X"809c0c51",
X"81135372",
X"882e0981",
X"06d93880",
X"5383c89c",
X"13335170",
X"81ff2eb2",
X"38701081",
X"d0900570",
X"22555180",
X"73177033",
X"701081d0",
X"90057022",
X"51515152",
X"5273712e",
X"91388112",
X"5271862e",
X"098106f1",
X"38739080",
X"9c0c8113",
X"5372862e",
X"098106ff",
X"b8388053",
X"72167033",
X"51517081",
X"ff2e9438",
X"701081d0",
X"90057022",
X"70848080",
X"0790809c",
X"0c515181",
X"13537286",
X"2e098106",
X"d7388053",
X"72165170",
X"3383c89c",
X"14348113",
X"5372862e",
X"098106ec",
X"38873d0d",
X"0404ff3d",
X"0d740284",
X"058f0533",
X"52527088",
X"38719080",
X"940c8e39",
X"70812e09",
X"81068638",
X"71908098",
X"0c833d0d",
X"04fb3d0d",
X"029f0533",
X"79982b70",
X"982c7c98",
X"2b70982c",
X"83c8b815",
X"70337098",
X"2b70982c",
X"51585c5a",
X"51555154",
X"5470732e",
X"09810694",
X"3883c898",
X"14337098",
X"2b70982c",
X"51525670",
X"722eb138",
X"72753471",
X"83c89815",
X"3483c899",
X"3383c8b9",
X"3371982b",
X"71902b07",
X"83c89833",
X"70882b72",
X"0783c8b8",
X"33710790",
X"80b80c52",
X"59535452",
X"873d0d04",
X"fe3d0d74",
X"81113371",
X"3371882b",
X"0783c080",
X"0c535184",
X"3d0d0483",
X"c8a43383",
X"c0800c04",
X"f53d0d02",
X"bb053302",
X"8405bf05",
X"33028805",
X"80c30533",
X"028c0580",
X"c6052266",
X"5c5a5e5c",
X"567a557b",
X"548953a1",
X"527d5180",
X"d2fb3f83",
X"c0800881",
X"ff0683c0",
X"800c8d3d",
X"0d0483c0",
X"8c080283",
X"c08c0cf5",
X"3d0d83c0",
X"8c088805",
X"0883c08c",
X"088f0533",
X"83c08c08",
X"92052202",
X"8c057390",
X"0583c08c",
X"08e8050c",
X"83c08c08",
X"f8050c83",
X"c08c08f0",
X"050c83c0",
X"8c08ec05",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08f005",
X"0883c08c",
X"08e0050c",
X"83c08c08",
X"fc050c83",
X"c08c08f0",
X"05088927",
X"8a38890b",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"05088605",
X"87fffc06",
X"83c08c08",
X"e0050c02",
X"83c08c08",
X"e0050831",
X"0d853d70",
X"5583c08c",
X"08ec0508",
X"5483c08c",
X"08f00508",
X"5383c08c",
X"08f40508",
X"5283c08c",
X"08e4050c",
X"80dcd43f",
X"83c08008",
X"81ff0683",
X"c08c08e4",
X"050883c0",
X"8c08ec05",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"e0050880",
X"2e8c3883",
X"c08c08f8",
X"05080d89",
X"c83983c0",
X"8c08f005",
X"08802e89",
X"a63883c0",
X"8c08ec05",
X"08810533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508842e",
X"a938840b",
X"83c08c08",
X"e0050825",
X"88c73883",
X"c08c08e0",
X"0508852e",
X"859b3883",
X"c08c08e0",
X"0508a12e",
X"87ad3888",
X"ac39800b",
X"83c08c08",
X"ec050885",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08fc050c",
X"83c08c08",
X"e0050883",
X"2e098106",
X"88833883",
X"c08c08e8",
X"05088105",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e0050881",
X"2687e638",
X"810b83c0",
X"8c08e005",
X"0880d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08fc",
X"050c83c0",
X"8c08ec05",
X"08820533",
X"83c08c08",
X"e0050887",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088b",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"e005088c",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088d",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"e005088e",
X"052383c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088a",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"70940508",
X"fcffff06",
X"7194050c",
X"83c08c08",
X"e0050c83",
X"c08c08ec",
X"05088605",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"f4050c83",
X"c08c08e0",
X"050883c0",
X"8c08fc05",
X"082e0981",
X"06b63883",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c83",
X"c08c08fc",
X"050883c0",
X"8c08e005",
X"088b0534",
X"83c08c08",
X"ec050887",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"812e8f38",
X"83c08c08",
X"e0050882",
X"2eb73884",
X"8c3983c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c820b",
X"83c08c08",
X"e005088a",
X"053483d9",
X"3983c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08fc0508",
X"83c08c08",
X"e005088a",
X"053483a1",
X"3983c08c",
X"08fc0508",
X"802e8395",
X"3883c08c",
X"08ec0508",
X"83053383",
X"0683c08c",
X"08e0050c",
X"83c08c08",
X"e0050883",
X"2e098106",
X"82f33883",
X"c08c08ec",
X"05088205",
X"3370982b",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c83c0",
X"8c08e005",
X"08802582",
X"cc3883c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c83c0",
X"8c08ec05",
X"08860533",
X"83c08c08",
X"e0050880",
X"d6053483",
X"c08c08e0",
X"05088405",
X"83c08c08",
X"ec050882",
X"05338f06",
X"83c08c08",
X"e4050c83",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0883c08c",
X"08e00508",
X"3483c08c",
X"08ec0508",
X"84053383",
X"c08c08e0",
X"05088105",
X"34800b83",
X"c08c08e0",
X"05088205",
X"3483c08c",
X"08e00508",
X"08ff83ff",
X"06828007",
X"83c08c08",
X"e005080c",
X"83c08c08",
X"e8050881",
X"05338105",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"050883c0",
X"8c08e805",
X"08810534",
X"81833983",
X"c08c08fc",
X"0508802e",
X"80f73883",
X"c08c08ec",
X"05088605",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e00508a2",
X"2e098106",
X"80d73883",
X"c08c08ec",
X"05088805",
X"3383c08c",
X"08ec0508",
X"87053371",
X"82802905",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c5283c0",
X"8c08e405",
X"0c83c08c",
X"08f4050c",
X"83c08c08",
X"e4050883",
X"c08c08e0",
X"05088805",
X"2383c08c",
X"08ec0508",
X"3383c08c",
X"08f00508",
X"71317083",
X"ffff0683",
X"c08c08f0",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08ec0508",
X"0583c08c",
X"08ec050c",
X"f6d03983",
X"c08c08f8",
X"05080d83",
X"c08c08f0",
X"050883c0",
X"8c08e005",
X"0c83c08c",
X"08f80508",
X"0d83c08c",
X"08e00508",
X"83c0800c",
X"8d3d0d83",
X"c08c0c04",
X"83c08c08",
X"0283c08c",
X"0ce63d0d",
X"83c08c08",
X"88050802",
X"840583c0",
X"8c08e805",
X"0c83c08c",
X"08d4050c",
X"800b83c8",
X"c03483c0",
X"8c08d405",
X"08900583",
X"c08c08c0",
X"050c800b",
X"83c08c08",
X"c0050834",
X"800b83c0",
X"8c08c005",
X"08810534",
X"800b83c0",
X"8c08c405",
X"0c83c08c",
X"08c40508",
X"80d82983",
X"c08c08c0",
X"05080583",
X"c08c08ff",
X"b4050c80",
X"0b83c08c",
X"08ffb405",
X"0880d805",
X"0c83c08c",
X"08ffb405",
X"08840583",
X"c08c08ff",
X"b4050c83",
X"c08c08c4",
X"050883c0",
X"8c08ffb4",
X"05083488",
X"0b83c08c",
X"08ffb405",
X"08810534",
X"800b83c0",
X"8c08ffb4",
X"05088205",
X"3483c08c",
X"08ffb405",
X"0808ffa1",
X"ff06a080",
X"0783c08c",
X"08ffb405",
X"080c83c0",
X"8c08c405",
X"08810570",
X"81ff0683",
X"c08c08c4",
X"050c83c0",
X"8c08ffb4",
X"050c810b",
X"83c08c08",
X"c4050827",
X"fedb3883",
X"c08c08ec",
X"05705483",
X"c08c08c8",
X"050c9252",
X"83c08c08",
X"d4050851",
X"80cffb3f",
X"83c08008",
X"81ff0670",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"8eb43883",
X"c08c08f4",
X"0551f18c",
X"3f83c080",
X"0883ffff",
X"0683c08c",
X"08f60552",
X"83c08c08",
X"e4050cf0",
X"f33f83c0",
X"800883ff",
X"ff0683c0",
X"8c08fd05",
X"3383c08c",
X"08ffb805",
X"0883c08c",
X"08c4050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"dc050c83",
X"c08c08c4",
X"050883c0",
X"8c08ffbc",
X"05082780",
X"fe3883c0",
X"8c08c805",
X"085483c0",
X"8c08c405",
X"08538952",
X"83c08c08",
X"d4050851",
X"80cf803f",
X"83c08008",
X"81ff0683",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b8050880",
X"f23883c0",
X"8c08ee05",
X"51eff13f",
X"83c08008",
X"83ffff06",
X"5383c08c",
X"08c40508",
X"5283c08c",
X"08d40508",
X"51f0b33f",
X"83c08c08",
X"c4050881",
X"057081ff",
X"0683c08c",
X"08c4050c",
X"83c08c08",
X"ffb4050c",
X"fef13983",
X"c08c08c0",
X"05088105",
X"3383c08c",
X"08ffb405",
X"0c81db0b",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb40508",
X"802e8caa",
X"38943983",
X"c08c08ff",
X"b8050883",
X"c08c08ff",
X"bc050c8c",
X"953983c0",
X"8c08f105",
X"335283c0",
X"8c08d405",
X"085180cd",
X"fe3f800b",
X"83c08c08",
X"c0050881",
X"053383c0",
X"8c08ffb4",
X"050c83c0",
X"8c08c405",
X"0c83c08c",
X"08c40508",
X"83c08c08",
X"ffb40508",
X"278ab038",
X"83c08c08",
X"c4050880",
X"d8297083",
X"c08c08c0",
X"05080570",
X"88057083",
X"053383c0",
X"8c08cc05",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"d8050c83",
X"c08c08cc",
X"050887f0",
X"3883c08c",
X"08c80508",
X"22028405",
X"71860587",
X"fffc0683",
X"c08c08ff",
X"b4050c83",
X"c08c08e0",
X"050c83c0",
X"8c08ffb8",
X"050c0283",
X"c08c08ff",
X"b4050831",
X"0d893d70",
X"5983c08c",
X"08ffb805",
X"085883c0",
X"8c08ffbc",
X"05088705",
X"335783c0",
X"8c08ffb4",
X"050ca255",
X"83c08c08",
X"cc050854",
X"86538181",
X"5283c08c",
X"08d40508",
X"5180c0cd",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"d0050c83",
X"c08c08d0",
X"050881c1",
X"3883c08c",
X"08ffbc05",
X"08960553",
X"83c08c08",
X"ffb80508",
X"5283c08c",
X"08ffb405",
X"0851a480",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb40508",
X"802e8185",
X"3883c08c",
X"08ffbc05",
X"08940583",
X"c08c08ff",
X"bc050896",
X"05337086",
X"2a83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08cc050c",
X"83c08c08",
X"ffb40508",
X"832e0981",
X"0680c638",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"c8050882",
X"053483c8",
X"a4337081",
X"0583c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb405",
X"0883c8a4",
X"3483c08c",
X"08ffb805",
X"0883c08c",
X"08cc0508",
X"3483c08c",
X"08e00508",
X"0d83c08c",
X"08d00508",
X"81ff0683",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b80508fb",
X"fe3883c0",
X"8c08d805",
X"0883c08c",
X"08c00508",
X"05880570",
X"82053351",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb40508",
X"832e0981",
X"0680e338",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb40508",
X"81057081",
X"ff065183",
X"c08c08ff",
X"b4050c81",
X"0b83c08c",
X"08ffb405",
X"0827dd38",
X"800b83c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb4",
X"05088105",
X"7081ff06",
X"5183c08c",
X"08ffb405",
X"0c970b83",
X"c08c08ff",
X"b4050827",
X"dd3883c0",
X"8c08e405",
X"0880f932",
X"70307080",
X"25515183",
X"c08c08ff",
X"b4050c83",
X"c08c08dc",
X"0508912e",
X"09810680",
X"f93883c0",
X"8c08ffb4",
X"0508802e",
X"80ec3883",
X"c08c08c4",
X"050880e2",
X"38850b83",
X"c08c08c0",
X"0508a605",
X"34a00b83",
X"c08c08c0",
X"0508a705",
X"34850b83",
X"c08c08c0",
X"0508a805",
X"3480c00b",
X"83c08c08",
X"c00508a9",
X"0534860b",
X"83c08c08",
X"c00508aa",
X"0534900b",
X"83c08c08",
X"c00508ab",
X"0534860b",
X"83c08c08",
X"c00508ac",
X"0534a00b",
X"83c08c08",
X"c00508ad",
X"053483c0",
X"8c08e405",
X"0889d832",
X"70307080",
X"25515183",
X"c08c08ff",
X"b4050c83",
X"c08c08dc",
X"050883ed",
X"ec2e0981",
X"0680f638",
X"817083c0",
X"8c08ffb4",
X"05080683",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b4050880",
X"2e80ce38",
X"83c08c08",
X"c4050880",
X"c438840b",
X"83c08c08",
X"c00508aa",
X"053480c0",
X"0b83c08c",
X"08c00508",
X"ab053484",
X"0b83c08c",
X"08c00508",
X"ac053490",
X"0b83c08c",
X"08c00508",
X"ad053483",
X"c08c08ff",
X"b8050883",
X"c08c08c0",
X"05088c05",
X"3483c08c",
X"08e40508",
X"80f93270",
X"30708025",
X"515183c0",
X"8c08ffb4",
X"050c83c0",
X"8c08dc05",
X"08862e09",
X"810680c3",
X"38817083",
X"c08c08ff",
X"b4050806",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb40508",
X"802e9c38",
X"83c08c08",
X"c4050893",
X"3883c08c",
X"08ffb805",
X"0883c08c",
X"08c00508",
X"8d053483",
X"c08c08e4",
X"0508b4b4",
X"32703070",
X"80255151",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"dc050890",
X"892e0981",
X"06a23883",
X"c08c08ff",
X"b4050880",
X"2e963883",
X"c08c08c4",
X"05088d38",
X"820b83c0",
X"8c08c005",
X"088d0534",
X"83c08c08",
X"c4050880",
X"d82983c0",
X"8c08c005",
X"08057084",
X"05708305",
X"3383c08c",
X"08ffb405",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"ffbc050c",
X"80588057",
X"83c08c08",
X"ffb40508",
X"56805580",
X"548a53a1",
X"5283c08c",
X"08d40508",
X"51b8fe3f",
X"83c08008",
X"81ff0670",
X"30709f2a",
X"5183c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"08a02e8c",
X"3883c08c",
X"08ffb405",
X"08f5f838",
X"83c08c08",
X"ffbc0508",
X"8b053383",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b4050880",
X"2eb33883",
X"c08c08c8",
X"05088305",
X"3383c08c",
X"08ffb405",
X"0c805880",
X"5783c08c",
X"08ffb405",
X"08568055",
X"80548b53",
X"a15283c0",
X"8c08d405",
X"0851b7f9",
X"3f83c08c",
X"08c40508",
X"81057081",
X"ff0683c0",
X"8c08c005",
X"08810533",
X"5283c08c",
X"08c4050c",
X"83c08c08",
X"ffb4050c",
X"f5bf3980",
X"0b83c08c",
X"08c4050c",
X"83c08c08",
X"c4050880",
X"d82983c0",
X"8c08d405",
X"0805709a",
X"053383c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb4",
X"0508822e",
X"098106a9",
X"3883c8c0",
X"56815580",
X"5483c08c",
X"08ffb405",
X"085383c0",
X"8c08ffb8",
X"05089705",
X"335283c0",
X"8c08d405",
X"0851e3c0",
X"3f83c08c",
X"08c40508",
X"81057081",
X"ff0683c0",
X"8c08c405",
X"0c83c08c",
X"08ffb405",
X"0c810b83",
X"c08c08c4",
X"050827fe",
X"fb38810b",
X"83c08c08",
X"c0050834",
X"800b83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08e805",
X"080d83c0",
X"8c08ffbc",
X"050883c0",
X"800c9c3d",
X"0d83c08c",
X"0c04f43d",
X"0d901f59",
X"800b811a",
X"33555b7a",
X"742781ad",
X"387a80d8",
X"29198a11",
X"33555573",
X"832e0981",
X"06818838",
X"94153357",
X"80527651",
X"e0f83f80",
X"53805276",
X"51e1963f",
X"aaed3f83",
X"c080085c",
X"80587781",
X"c4291c87",
X"11335555",
X"73802e80",
X"c0387408",
X"81d0842e",
X"098106b5",
X"3880755b",
X"567580d8",
X"291a9a11",
X"33555573",
X"832e0981",
X"069238a4",
X"15703355",
X"55767427",
X"8738ff14",
X"54737534",
X"81167081",
X"ff065754",
X"817627d1",
X"38811870",
X"81ff0659",
X"548f7827",
X"ffa43883",
X"c8a433ff",
X"05547383",
X"c8a43481",
X"1b7081ff",
X"06811b33",
X"5f5c547c",
X"7b26fed5",
X"38800b83",
X"c0800c8e",
X"3d0d0483",
X"c08c0802",
X"83c08c0c",
X"e63d0d83",
X"c08c0888",
X"05080284",
X"05719005",
X"70337083",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08c8",
X"050c83c0",
X"8c08dc05",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"ffa40508",
X"802e9696",
X"38800b83",
X"c08c08c8",
X"05088105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08d0050c",
X"83c08c08",
X"d0050883",
X"c08c08ff",
X"a4050825",
X"95de3883",
X"c08c08d0",
X"050880d8",
X"2983c08c",
X"08c80508",
X"05840570",
X"86053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"a4050880",
X"2e94ea38",
X"a8933f83",
X"c08c08ff",
X"bc050880",
X"d4050883",
X"c0800826",
X"94d33802",
X"83c08c08",
X"ffbc0508",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08d8",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08fc05",
X"2383c08c",
X"08ffa405",
X"08860583",
X"fc0683c0",
X"8c08ffa4",
X"050c0283",
X"c08c08ff",
X"a4050831",
X"0d853d70",
X"5583c08c",
X"08fc0554",
X"83c08c08",
X"ffbc0508",
X"5383c08c",
X"08e00508",
X"5283c08c",
X"08c4050c",
X"afeb3f83",
X"c0800881",
X"ff0683c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508939c",
X"3883c08c",
X"08ffbc05",
X"08870533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e80d5",
X"3883c08c",
X"08ffbc05",
X"08860533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"822e0981",
X"06b33883",
X"c08c08fc",
X"052283c0",
X"8c08ffa4",
X"050c870b",
X"83c08c08",
X"ffa40508",
X"27973883",
X"c08c08c4",
X"05088205",
X"5283c08c",
X"08c40508",
X"3351dacc",
X"3f83c08c",
X"08ffbc05",
X"08860533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"832e0981",
X"06928538",
X"83c08c08",
X"ffbc0508",
X"92057082",
X"053383c0",
X"8c08fc05",
X"2283c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08c0050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffa80508",
X"2691c538",
X"800b83c0",
X"8c08e405",
X"0c800b83",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"b0050810",
X"83c08c08",
X"05f80583",
X"c08c08ff",
X"b0050884",
X"2983c08c",
X"08ffb005",
X"08100583",
X"c08c08c0",
X"05080570",
X"84057033",
X"83c08c08",
X"c4050805",
X"703383c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffb8",
X"05082383",
X"c08c08ff",
X"a8050881",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508902e",
X"098106be",
X"3883c08c",
X"08ffa805",
X"083383c0",
X"8c08c405",
X"08058105",
X"70337082",
X"802983c0",
X"8c08ffb4",
X"05080551",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffb805",
X"082383c0",
X"8c08ffac",
X"05088605",
X"2283c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa805",
X"08a23883",
X"c08c08ff",
X"ac050888",
X"052283c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"050881ff",
X"2e80e538",
X"83c08c08",
X"ffb80508",
X"227083c0",
X"8c08ffa8",
X"05083170",
X"82802971",
X"3183c08c",
X"08ffac05",
X"08880522",
X"7083c08c",
X"08ffa805",
X"08317073",
X"355383c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c5183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"b8050823",
X"83c08c08",
X"ffb00508",
X"81057081",
X"ff0683c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa4",
X"050c810b",
X"83c08c08",
X"ffb00508",
X"27fce038",
X"83c08c08",
X"f8052283",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a40508bf",
X"26913883",
X"c08c08e4",
X"05088207",
X"83c08c08",
X"e4050c81",
X"c00b83c0",
X"8c08ffa4",
X"05082791",
X"3883c08c",
X"08e40508",
X"810783c0",
X"8c08e405",
X"0c83c08c",
X"08fa0522",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"bf269138",
X"83c08c08",
X"e4050888",
X"0783c08c",
X"08e4050c",
X"81c00b83",
X"c08c08ff",
X"a4050827",
X"913883c0",
X"8c08e405",
X"08840783",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffb00508",
X"1083c08c",
X"08c00508",
X"05709005",
X"703383c0",
X"8c08c405",
X"08057033",
X"72810533",
X"70720651",
X"535183c0",
X"8c08ffa8",
X"050c5183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e9b3890",
X"0b83c08c",
X"08ffb005",
X"082b83c0",
X"8c08e405",
X"080783c0",
X"8c08e405",
X"0c83c08c",
X"08ffb005",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a4050c97",
X"0b83c08c",
X"08ffb005",
X"0827fef4",
X"3883c08c",
X"08ffbc05",
X"08900533",
X"83c08c08",
X"e4050883",
X"c08c08ff",
X"a4050c83",
X"c08c08c0",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffbc",
X"05088c05",
X"082e85e0",
X"3883c08c",
X"08ffa405",
X"0883c08c",
X"08ffbc05",
X"088c050c",
X"83c08c08",
X"ffbc0508",
X"89053383",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a8050880",
X"2e859a38",
X"83c08c08",
X"e40583c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffa4",
X"05088f06",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"b0050c83",
X"c08c08d4",
X"050c83c0",
X"8c08ffa8",
X"0508822e",
X"09810681",
X"c238800b",
X"83c08c08",
X"ffa40508",
X"862a7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffa8",
X"05082e8c",
X"3881c00b",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffb00508",
X"872a7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"943883c0",
X"8c08ffa8",
X"05088190",
X"3283c08c",
X"08ffa805",
X"0c83c08c",
X"08ffb005",
X"08842a70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e943883",
X"c08c08ff",
X"a8050880",
X"d03283c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffb0",
X"050883c0",
X"8c08ffa8",
X"05083283",
X"c08c08ff",
X"b0050c80",
X"0b83c08c",
X"08f0050c",
X"800b83c0",
X"8c08f405",
X"23800b81",
X"d2803383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"b805082e",
X"82d33883",
X"c08c08f0",
X"0581d280",
X"0b83c08c",
X"08ffac05",
X"0c83c08c",
X"08cc050c",
X"83c08c08",
X"ffac0508",
X"3383c08c",
X"08ffac05",
X"08810533",
X"81722b81",
X"722b0770",
X"83c08c08",
X"ffb00508",
X"065283c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffa8",
X"05082e09",
X"810681be",
X"3883c08c",
X"08ffb805",
X"08852680",
X"f63883c0",
X"8c08ffac",
X"05088205",
X"337081ff",
X"0683c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"08802e80",
X"ca3883c0",
X"8c08ffb8",
X"050883c0",
X"8c08ffb8",
X"05088105",
X"7081ff06",
X"83c08c08",
X"cc050873",
X"055383c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffa4",
X"05083483",
X"c08c08ff",
X"ac050883",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"9d38810b",
X"83c08c08",
X"ffa40508",
X"2b83c08c",
X"08d40508",
X"080783c0",
X"8c08d405",
X"080c83c0",
X"8c08ffac",
X"05088405",
X"703383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa4",
X"0508fdc8",
X"3883c08c",
X"08f00552",
X"8051ce88",
X"3f83c08c",
X"08e40508",
X"5283c08c",
X"08c00508",
X"51cfc33f",
X"83c08c08",
X"fb053370",
X"81800a29",
X"810a0570",
X"982c5583",
X"c08c08ff",
X"a4050c83",
X"c08c08f9",
X"05337081",
X"800a2981",
X"0a057098",
X"2c5583c0",
X"8c08ffa4",
X"050c83c0",
X"8c08c005",
X"085383c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa8",
X"050ccf99",
X"3f83c08c",
X"08ffbc05",
X"08880533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e84e0",
X"3883c08c",
X"08ffbc05",
X"08900533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"812684c0",
X"38807081",
X"d2b80b81",
X"d2b80b81",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffb4",
X"05082e81",
X"ae3883c0",
X"8c08ffac",
X"05088429",
X"83c08c08",
X"ffa80508",
X"05703383",
X"c08c08c4",
X"05080570",
X"33728105",
X"33707206",
X"51535183",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2eaa3881",
X"0b83c08c",
X"08ffac05",
X"082b83c0",
X"8c08ffb4",
X"05080770",
X"83ffff06",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffac0508",
X"81057081",
X"ff0681d2",
X"b8718429",
X"71057081",
X"05335153",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"fed43883",
X"c08c08ff",
X"bc05088a",
X"052283c0",
X"8c08c005",
X"0c83c08c",
X"08ffb405",
X"0883c08c",
X"08c00508",
X"2e82ad38",
X"800b83c0",
X"8c08e805",
X"0c800b83",
X"c08c08ec",
X"05238070",
X"83c08c08",
X"e80583c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffb0",
X"050c81af",
X"3983c08c",
X"08ffb405",
X"0883c08c",
X"08ffac05",
X"082c7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"80e73883",
X"c08c08ff",
X"b0050883",
X"c08c08ff",
X"b0050881",
X"057081ff",
X"0683c08c",
X"08ffb805",
X"08730583",
X"c08c08ff",
X"bc050890",
X"053383c0",
X"8c08ffac",
X"05088429",
X"05535383",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a8050881",
X"d2ba0533",
X"83c08c08",
X"ffa40508",
X"3483c08c",
X"08ffac05",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a4050c8f",
X"0b83c08c",
X"08ffac05",
X"082783c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb0",
X"05088526",
X"8c3883c0",
X"8c08ffa4",
X"0508fea9",
X"3883c08c",
X"08e80552",
X"8051c8b8",
X"3f83c08c",
X"08ffb405",
X"0883c08c",
X"08ffbc05",
X"088a0523",
X"83c08c08",
X"ffbc0508",
X"80d20533",
X"83c08c08",
X"ffbc0508",
X"80d40508",
X"0583c08c",
X"08ffbc05",
X"0880d405",
X"0c83c08c",
X"08d80508",
X"0d83c08c",
X"08d00508",
X"81800a29",
X"81800a05",
X"70982c83",
X"c08c08c8",
X"05088105",
X"3383c08c",
X"08ffa805",
X"0c5183c0",
X"8c08d005",
X"0c83c08c",
X"08ffa805",
X"0883c08c",
X"08d00508",
X"24eaa438",
X"800b83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08dc05",
X"080d83c0",
X"8c08ffa8",
X"050883c0",
X"800c9c3d",
X"0d83c08c",
X"0c04f33d",
X"0d02bf05",
X"33028405",
X"80c30533",
X"83c8c033",
X"5a5b5979",
X"802e8d38",
X"78780657",
X"76802e8e",
X"38818939",
X"78780657",
X"76802e80",
X"ff3883c8",
X"c033707a",
X"07585879",
X"88387809",
X"70790651",
X"577683c8",
X"c0349297",
X"3f83c080",
X"085e805c",
X"8f5d7d1c",
X"87113358",
X"5876802e",
X"80c13877",
X"0881d084",
X"2e098106",
X"b638805b",
X"815a7d1c",
X"701c9a11",
X"33595959",
X"76822e09",
X"81069438",
X"83c8c056",
X"81558054",
X"76539718",
X"33527851",
X"c98a3fff",
X"1a80d81c",
X"5c5a7980",
X"25d038ff",
X"1d81c41d",
X"5d5d7c80",
X"25ffa738",
X"8f3d0d04",
X"e93d0d69",
X"6c028805",
X"80ea0522",
X"5c5a5b80",
X"7071415e",
X"58ff7879",
X"7a7b7c7d",
X"464c4a45",
X"405d4362",
X"993d3462",
X"02840580",
X"dd053477",
X"792280ff",
X"ff065445",
X"72792379",
X"782e8887",
X"387a7081",
X"055c3370",
X"842a718c",
X"0670822a",
X"5a565683",
X"06ff1b70",
X"83ffff06",
X"5c545680",
X"5475742e",
X"91387a70",
X"81055c33",
X"ff1b7083",
X"ffff065c",
X"54548176",
X"279b3873",
X"81ff067b",
X"7081055d",
X"33557482",
X"802905ff",
X"1b7083ff",
X"ff065c54",
X"54827627",
X"aa387383",
X"ffff067b",
X"7081055d",
X"3370902b",
X"72077d70",
X"81055f33",
X"70982b72",
X"07fe1f70",
X"83ffff06",
X"40525252",
X"5254547e",
X"802e80c4",
X"387686f7",
X"38748a2e",
X"09810694",
X"38811f70",
X"81ff0681",
X"1e7081ff",
X"065f5240",
X"5386dc39",
X"748c2e09",
X"810686d3",
X"38ff1f70",
X"81ff06ff",
X"1e7081ff",
X"065f5240",
X"537b6325",
X"86bd38ff",
X"4386b839",
X"76812e83",
X"bb387681",
X"24893876",
X"802e8d38",
X"86a53976",
X"822e84a6",
X"38869c39",
X"f8155372",
X"84268495",
X"38728429",
X"81d2f805",
X"53720804",
X"64802e80",
X"cd387822",
X"83808006",
X"53728380",
X"802e0981",
X"06bc3880",
X"56756427",
X"a438751e",
X"7083ffff",
X"0677101b",
X"90117283",
X"2a585157",
X"51537375",
X"34728706",
X"81712b51",
X"53728116",
X"34811670",
X"81ff0657",
X"53977627",
X"cc387f84",
X"0740800b",
X"993d4356",
X"61167033",
X"70982b70",
X"982c5151",
X"51538073",
X"2480fb38",
X"6073291e",
X"7083ffff",
X"067a2283",
X"80800652",
X"58537283",
X"80802e09",
X"810680de",
X"38608832",
X"70307072",
X"07802563",
X"90327030",
X"70720780",
X"25730753",
X"54585155",
X"5373802e",
X"bd387687",
X"065372b6",
X"38758429",
X"76100579",
X"11841179",
X"832a5757",
X"51537375",
X"34608116",
X"34658614",
X"23668814",
X"23758738",
X"7f810740",
X"8d397581",
X"2e098106",
X"85387f82",
X"07408116",
X"7081ff06",
X"57538176",
X"27fee538",
X"6361291e",
X"7083ffff",
X"065f5380",
X"704642ff",
X"02840580",
X"dd0534ff",
X"0b993d34",
X"83f53981",
X"1c7081ff",
X"065d5380",
X"4273812e",
X"0981068e",
X"38778180",
X"0a298180",
X"0a055880",
X"d3397380",
X"2e893873",
X"822e0981",
X"068d387c",
X"81800a29",
X"81800a05",
X"5da43981",
X"5f83b839",
X"ff1c7081",
X"ff065d53",
X"7b632583",
X"38ff437c",
X"802e9238",
X"7c81800a",
X"2981ff0a",
X"055d7c98",
X"2c5d8393",
X"3977802e",
X"92387781",
X"800a2981",
X"ff0a0558",
X"77982c58",
X"82fd3977",
X"53839e39",
X"74892680",
X"f4387484",
X"2981d38c",
X"05537208",
X"0473872e",
X"82e13873",
X"852e82db",
X"3873882e",
X"82d53873",
X"8c2e82cf",
X"3873892e",
X"09810686",
X"38814582",
X"c2397381",
X"2e098106",
X"82b93862",
X"802582b3",
X"387b982b",
X"70982c51",
X"4382a839",
X"7383ffff",
X"0646829f",
X"397383ff",
X"ff064782",
X"96397381",
X"ff064182",
X"8e397381",
X"1a348287",
X"397381ff",
X"064481ff",
X"397e5382",
X"a0397481",
X"2e81e338",
X"74812489",
X"3874802e",
X"8d3881e7",
X"3974822e",
X"81d83881",
X"de397456",
X"7b833881",
X"56745373",
X"862e0981",
X"06973875",
X"81065372",
X"802e8e38",
X"782282ff",
X"ff06fe80",
X"800753b6",
X"397b8338",
X"81537382",
X"2e098106",
X"97387281",
X"06537280",
X"2e8e3878",
X"2281ffff",
X"06818080",
X"07539339",
X"7b9638fc",
X"14537281",
X"268e3878",
X"22ff8080",
X"07537279",
X"2380e539",
X"80557381",
X"2e098106",
X"83387355",
X"77537780",
X"2e893874",
X"81065372",
X"80ca3872",
X"d0155455",
X"72812683",
X"38815577",
X"802eb938",
X"74810653",
X"72802eb0",
X"38782283",
X"80800653",
X"72838080",
X"2e098106",
X"9f3873b0",
X"2e098106",
X"87386199",
X"3d349139",
X"73b12e09",
X"81068938",
X"61028405",
X"80dd0534",
X"61810553",
X"8c396174",
X"31810553",
X"84396114",
X"537283ff",
X"ff064279",
X"f7fb387d",
X"832a5372",
X"821a3478",
X"22838080",
X"06537283",
X"80802e09",
X"81068838",
X"81537f87",
X"2e833880",
X"537283c0",
X"800c993d",
X"0d04fd3d",
X"0d758311",
X"33821233",
X"71982b71",
X"902b0781",
X"14337088",
X"2b720775",
X"33710783",
X"c0800c52",
X"53545654",
X"52853d0d",
X"04f63d0d",
X"02b70533",
X"028405bb",
X"05330288",
X"05bf0533",
X"5b5b5b80",
X"58805778",
X"882b7a07",
X"5680557a",
X"548153a3",
X"527c5192",
X"cc3f83c0",
X"800881ff",
X"0683c080",
X"0c8c3d0d",
X"04f63d0d",
X"02b70533",
X"028405bb",
X"05330288",
X"05bf0533",
X"5b5b5b80",
X"58805778",
X"882b7a07",
X"5680557a",
X"548353a3",
X"527c5192",
X"903f83c0",
X"800881ff",
X"0683c080",
X"0c8c3d0d",
X"04f73d0d",
X"02b30533",
X"028405b6",
X"0522605a",
X"58568055",
X"80548053",
X"81a3527b",
X"5191e23f",
X"83c08008",
X"81ff0683",
X"c0800c8b",
X"3d0d04ee",
X"3d0d6490",
X"115c5c80",
X"7b34800b",
X"841c0c80",
X"0b881c34",
X"810b891c",
X"34880b8a",
X"1c34800b",
X"8b1c3488",
X"1b08c106",
X"8107881c",
X"0c8f3d70",
X"545d8852",
X"7b519c92",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"81a93890",
X"3d335e81",
X"db5a7d89",
X"2e098106",
X"8199387c",
X"5392527b",
X"519beb3f",
X"83c08008",
X"81ff0670",
X"5b597881",
X"82387c58",
X"88577856",
X"a9557854",
X"865381a0",
X"527b5190",
X"d03f83c0",
X"800881ff",
X"06705b59",
X"7880e038",
X"02ba0533",
X"7b347c54",
X"78537d52",
X"7b519bd3",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"80c13802",
X"bd053352",
X"7b519beb",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"aa38817b",
X"335a5a79",
X"79269938",
X"80547953",
X"88527b51",
X"fdbb3f81",
X"1a7081ff",
X"067c3352",
X"5b59e439",
X"810b881c",
X"34805a79",
X"83c0800c",
X"943d0d04",
X"800b83c0",
X"800c04f9",
X"3d0d7902",
X"8405ab05",
X"338e3d70",
X"54585858",
X"ffbbf53f",
X"8a3d8a05",
X"51ffbbec",
X"3f7551fc",
X"8d3f83c0",
X"80088486",
X"812ebe38",
X"83c08008",
X"84868126",
X"993883c0",
X"80088482",
X"802e80e6",
X"3883c080",
X"08848281",
X"2e9f3881",
X"b43983c0",
X"800880c0",
X"82832e80",
X"f43883c0",
X"800880c0",
X"86832e80",
X"e8388199",
X"3983c09c",
X"33558056",
X"74762e09",
X"8106818b",
X"38745476",
X"53915277",
X"51fbd63f",
X"74547653",
X"90527751",
X"fbcb3f74",
X"54765384",
X"527751fb",
X"fc3f810b",
X"83c09c34",
X"81b15680",
X"de398054",
X"76539152",
X"7751fba9",
X"3f805476",
X"53905277",
X"51fb9e3f",
X"800b83c0",
X"9c347652",
X"87183351",
X"97963fb5",
X"39805476",
X"53945277",
X"51fb823f",
X"80547653",
X"90527751",
X"faf73f75",
X"51ffbaa0",
X"3f83c080",
X"08892a81",
X"06537652",
X"87183351",
X"90cd3f80",
X"0b83c09c",
X"34805675",
X"83c0800c",
X"893d0d04",
X"f23d0d60",
X"90115a58",
X"800b881a",
X"33715956",
X"5674762e",
X"82a53882",
X"ac3f8419",
X"0883c080",
X"08268295",
X"3878335a",
X"810b8e3d",
X"23903df8",
X"1155f405",
X"53991852",
X"77518ae5",
X"3f83c080",
X"0881ff06",
X"70575574",
X"772e0981",
X"0681d938",
X"86397456",
X"81d23981",
X"5682578e",
X"3d337706",
X"5574802e",
X"bb38800b",
X"8d3d3490",
X"3df00554",
X"84537552",
X"7751facd",
X"3f83c080",
X"0881ff06",
X"55749d38",
X"7b537552",
X"7751fce7",
X"3f83c080",
X"0881ff06",
X"557481b1",
X"2e818b38",
X"74ffb338",
X"761081fc",
X"06811770",
X"81ff0658",
X"56578776",
X"27ffa838",
X"8156757a",
X"2680eb38",
X"800b8d3d",
X"348c3d70",
X"55578453",
X"75527751",
X"f9f73f83",
X"c0800881",
X"ff065574",
X"80c13876",
X"51ffb89c",
X"3f83c080",
X"08828706",
X"55748281",
X"2e098106",
X"aa3802ae",
X"05338107",
X"55740284",
X"05ae0534",
X"7b537552",
X"7751fbeb",
X"3f83c080",
X"0881ff06",
X"557481b1",
X"2e903874",
X"feb83881",
X"167081ff",
X"065755ff",
X"91398056",
X"7581ff06",
X"56973f83",
X"c080088f",
X"d005841a",
X"0c755776",
X"83c0800c",
X"903d0d04",
X"049080a0",
X"0883c080",
X"0c04ff3d",
X"0d7387e8",
X"2951ff9e",
X"f13f833d",
X"0d040483",
X"c8c40b83",
X"c0800c04",
X"fd3d0d75",
X"77545480",
X"0b83c8a4",
X"34728a38",
X"9090800b",
X"84150c90",
X"3972812e",
X"09810688",
X"38909880",
X"0b84150c",
X"84140883",
X"c8bc0c80",
X"0b88150c",
X"800b8c15",
X"0c83c8bc",
X"0853820b",
X"87801434",
X"8151ff9e",
X"3f83c8bc",
X"0853800b",
X"88143483",
X"c8bc0853",
X"810b8780",
X"143483c8",
X"bc085380",
X"0b8c1434",
X"83c8bc08",
X"53800ba4",
X"14349174",
X"34800b83",
X"c0a03480",
X"0b83c0a4",
X"34800b83",
X"c0a83480",
X"547381c4",
X"2983c8c8",
X"0553800b",
X"83143481",
X"147081ff",
X"0655538f",
X"7427e638",
X"853d0d04",
X"fe3d0d74",
X"76821133",
X"70bf0681",
X"712bff05",
X"56515152",
X"53907127",
X"8338ff52",
X"76517171",
X"2383c8bc",
X"08518713",
X"33901234",
X"800b83c0",
X"a434800b",
X"83c0a834",
X"8813338a",
X"14335252",
X"71802eaa",
X"387081ff",
X"06518452",
X"70833870",
X"527183c0",
X"a4348a13",
X"33703070",
X"8025842b",
X"70880751",
X"51525370",
X"83c0a834",
X"90397081",
X"ff065170",
X"83389852",
X"7183c0a8",
X"34800b83",
X"c0800c84",
X"3d0d04f1",
X"3d0d6165",
X"68028c05",
X"80cb0533",
X"02900580",
X"ce052202",
X"940580d6",
X"05224240",
X"415a4040",
X"fd8b3f83",
X"c08008a7",
X"88055b80",
X"70715b5b",
X"52839439",
X"83c8bc08",
X"517d9412",
X"3483c0a4",
X"33810755",
X"80705456",
X"7f862680",
X"ea387f84",
X"2981d3c0",
X"0583c8bc",
X"08535170",
X"0804800b",
X"841334a1",
X"39773370",
X"30708025",
X"83713151",
X"51525370",
X"8413348d",
X"39810b84",
X"1334b839",
X"830b8413",
X"34817054",
X"56ad3981",
X"0b841334",
X"a2397733",
X"70307080",
X"25837131",
X"51515253",
X"70841334",
X"80783352",
X"52708338",
X"81527178",
X"34815374",
X"88075583",
X"c0a83383",
X"c8bc0852",
X"57810b81",
X"d0123483",
X"c8bc0851",
X"810b8190",
X"12347e80",
X"2eae3872",
X"802ea938",
X"7eff1e52",
X"547083ff",
X"ff065372",
X"83ffff2e",
X"97387370",
X"81055533",
X"83c8bc08",
X"53517081",
X"c01334ff",
X"1351de39",
X"83c8bc08",
X"a8113353",
X"51768812",
X"3483c8bc",
X"08517471",
X"3481ff52",
X"913983c8",
X"bc08a011",
X"33708106",
X"51525370",
X"8f38fafd",
X"3f7a83c0",
X"800826e6",
X"38818839",
X"810ba014",
X"3483c8bc",
X"08a81133",
X"80ff0670",
X"78075253",
X"5170802e",
X"80ed3871",
X"862a7081",
X"06515170",
X"802e9138",
X"80783352",
X"53708338",
X"81537278",
X"3480e039",
X"71842a70",
X"81065151",
X"70802e9b",
X"38811970",
X"83ffff06",
X"7d30709f",
X"2a51525a",
X"51787c2e",
X"098106af",
X"38a43971",
X"832a7081",
X"06515170",
X"802e9338",
X"811a7081",
X"ff065b51",
X"79832e09",
X"81069038",
X"8a3971a3",
X"06517080",
X"2e853871",
X"519239f9",
X"e43f7a83",
X"c0800826",
X"fce23871",
X"81bf0651",
X"7083c080",
X"0c913d0d",
X"04f63d0d",
X"02b30533",
X"028405b7",
X"05330288",
X"05ba0522",
X"59595980",
X"0b8c3d34",
X"8c3dfc05",
X"56805580",
X"54765377",
X"527851fb",
X"f23f83c0",
X"800881ff",
X"0683c080",
X"0c8c3d0d",
X"04f33d0d",
X"7f626402",
X"8c0580c2",
X"05227222",
X"81153342",
X"5f415e59",
X"59807823",
X"7d537833",
X"528151ff",
X"a03f83c0",
X"800881ff",
X"06567580",
X"2e863875",
X"5481ad39",
X"83c8bc08",
X"a8113382",
X"1b337086",
X"2a708106",
X"73982b53",
X"51575c56",
X"57798025",
X"83388156",
X"73762e87",
X"3881f054",
X"81823981",
X"8c173370",
X"81ff0679",
X"227d7131",
X"902b7090",
X"2c700970",
X"9f2c7206",
X"70525253",
X"51535757",
X"54757424",
X"83387555",
X"74848080",
X"29fc8080",
X"0570902c",
X"515574ff",
X"2e943883",
X"c8bc0881",
X"80113351",
X"54737c70",
X"81055e34",
X"db397722",
X"76055473",
X"78237909",
X"709f2a70",
X"8106821c",
X"3381bf06",
X"71862b07",
X"51515154",
X"73821a34",
X"7c76268a",
X"38772254",
X"7a7426fe",
X"bb388054",
X"7383c080",
X"0c8f3d0d",
X"04f93d0d",
X"7a57800b",
X"893d2389",
X"3dfc0553",
X"76527951",
X"f8da3f83",
X"c0800881",
X"ff067057",
X"55749638",
X"7c547b53",
X"883d2252",
X"7651fde5",
X"3f83c080",
X"0881ff06",
X"567583c0",
X"800c893d",
X"0d04f03d",
X"0d626602",
X"880580ce",
X"0522415d",
X"5e800284",
X"0580d205",
X"227f8105",
X"33ff115a",
X"5d5a5d81",
X"da5876bf",
X"2680e938",
X"78802e80",
X"e1387a58",
X"787b2783",
X"38785882",
X"1e337087",
X"2a585a76",
X"923d3492",
X"3dfc0556",
X"77557b54",
X"7e537d33",
X"528251f8",
X"de3f83c0",
X"800881ff",
X"065d800b",
X"923d3358",
X"5a76802e",
X"8338815a",
X"821e3380",
X"ff067a87",
X"2b075776",
X"821f347c",
X"91387878",
X"317083ff",
X"ff06791e",
X"5e5a57ff",
X"9b397c58",
X"7783c080",
X"0c923d0d",
X"04f83d0d",
X"7b028405",
X"b2052258",
X"58800b8a",
X"3d238a3d",
X"fc055377",
X"527a51f6",
X"f73f83c0",
X"800881ff",
X"06705755",
X"7496387d",
X"54765389",
X"3d225277",
X"51feaf3f",
X"83c08008",
X"81ff0656",
X"7583c080",
X"0c8a3d0d",
X"04ec3d0d",
X"666e0288",
X"0580df05",
X"33028c05",
X"80e30533",
X"02900580",
X"e7053302",
X"940580eb",
X"05330298",
X"0580ee05",
X"22414341",
X"5f5c4057",
X"0280f205",
X"22963d23",
X"963df005",
X"53841770",
X"53775259",
X"f6863f83",
X"c0800881",
X"ff065877",
X"81e53877",
X"7a818006",
X"58408077",
X"25833881",
X"4079943d",
X"347b0284",
X"0580c905",
X"347c0284",
X"0580ca05",
X"347d0284",
X"0580cb05",
X"347a953d",
X"347a882a",
X"57760284",
X"0580cd05",
X"34953d22",
X"57760284",
X"0580ce05",
X"3476882a",
X"57760284",
X"0580cf05",
X"3477923d",
X"34963dec",
X"11575788",
X"55f41754",
X"923d2253",
X"77527751",
X"f6953f83",
X"c0800881",
X"ff065877",
X"80ed387e",
X"802e80cb",
X"38923d22",
X"79085858",
X"7f802e9c",
X"38768180",
X"8007790c",
X"7e54963d",
X"fc055377",
X"83ffff06",
X"527851f9",
X"fc3f9939",
X"76828080",
X"07790c7e",
X"54953d22",
X"537783ff",
X"ff065278",
X"51fc8f3f",
X"83c08008",
X"81ff0658",
X"779d3892",
X"3d225380",
X"527f3070",
X"80258471",
X"31535157",
X"f9873f83",
X"c0800881",
X"ff065877",
X"83c0800c",
X"963d0d04",
X"f63d0d7c",
X"028405b7",
X"05335b5b",
X"80588057",
X"80568055",
X"79548553",
X"80527a51",
X"fda33f83",
X"c0800881",
X"ff065978",
X"85387987",
X"1c347883",
X"c0800c8c",
X"3d0d04f9",
X"3d0d02a7",
X"05330284",
X"05ab0533",
X"028805af",
X"05335859",
X"57800b83",
X"c8cb3354",
X"5472742e",
X"9f388114",
X"7081ff06",
X"5553738f",
X"2681b638",
X"7381c429",
X"83c8c805",
X"83113351",
X"5372e338",
X"7381c429",
X"83c8c405",
X"55800b87",
X"16347688",
X"1634758a",
X"16347789",
X"16348075",
X"0c83c8bc",
X"088c160c",
X"800b8416",
X"34880b85",
X"1634800b",
X"86163484",
X"1508ffa1",
X"ff06a080",
X"0784160c",
X"81147081",
X"ff065353",
X"7451febc",
X"3f83c080",
X"0881ff06",
X"70555372",
X"80cd388a",
X"39730875",
X"0c725480",
X"c2397281",
X"d6d45556",
X"81d6d408",
X"802eb238",
X"75842914",
X"70087653",
X"70085154",
X"54722d83",
X"c0800881",
X"ff065372",
X"802ece38",
X"81167081",
X"ff0681d6",
X"d4718429",
X"11535657",
X"537208d0",
X"38805473",
X"83c0800c",
X"893d0d04",
X"f93d0d79",
X"57800b84",
X"180883c8",
X"bc0c58f0",
X"883f8817",
X"0883c080",
X"082783ed",
X"38effa3f",
X"83c08008",
X"81058818",
X"0c83c8bc",
X"08b81133",
X"7081ff06",
X"51515473",
X"812ea438",
X"73812488",
X"3873782e",
X"8a38b839",
X"73822e95",
X"38b13976",
X"3381f006",
X"5473902e",
X"a6389177",
X"34a13973",
X"58763381",
X"f0065473",
X"902e0981",
X"069138ef",
X"a83f83c0",
X"800881c8",
X"058c180c",
X"a0773480",
X"567581c4",
X"2983c8cb",
X"11335555",
X"73802eaa",
X"3883c8c4",
X"15700856",
X"5474802e",
X"9d388815",
X"08802e96",
X"388c1408",
X"83c8bc08",
X"2e098106",
X"89387351",
X"88150854",
X"732d8116",
X"7081ff06",
X"57548f76",
X"27ffba38",
X"76335473",
X"b02e8199",
X"3873b024",
X"8f387391",
X"2eab3873",
X"a02e80f5",
X"3882a639",
X"7380d02e",
X"81e43873",
X"80d0248b",
X"387380c0",
X"2e819938",
X"828f3973",
X"81802e81",
X"fb388285",
X"39805675",
X"81c42983",
X"c8c81183",
X"11335659",
X"5573802e",
X"a83883c8",
X"c4157008",
X"56547480",
X"2e9b388c",
X"140883c8",
X"bc082e09",
X"81068e38",
X"73518415",
X"0854732d",
X"800b8319",
X"34811670",
X"81ff0657",
X"548f7627",
X"ffb93892",
X"773481b5",
X"39edc23f",
X"8c170883",
X"c0800827",
X"81a738b0",
X"773481a1",
X"3983c8bc",
X"0854800b",
X"8c153483",
X"c8bc0854",
X"840b8815",
X"3480c077",
X"34ed963f",
X"83c08008",
X"b2058c18",
X"0c80fa39",
X"ed873f8c",
X"170883c0",
X"80082780",
X"ec3883c8",
X"bc085481",
X"0b8c1534",
X"83c8bc08",
X"54800b88",
X"153483c8",
X"bc085488",
X"0ba01534",
X"ecdb3f83",
X"c0800894",
X"058c180c",
X"80d07734",
X"bc3983c8",
X"bc08a011",
X"3370832a",
X"70810651",
X"51555573",
X"802ea638",
X"880ba016",
X"34ecae3f",
X"8c170883",
X"c0800827",
X"9438ff80",
X"77348e39",
X"77538052",
X"8051fa8b",
X"3fff9077",
X"3483c8bc",
X"08a01133",
X"70832a70",
X"81065151",
X"55557380",
X"2e863888",
X"0ba01634",
X"893d0d04",
X"f43d0d02",
X"bb053302",
X"8405bf05",
X"335d5d80",
X"0b83c8c8",
X"0b83c8c4",
X"0b8c1172",
X"71881475",
X"5c5a5b5f",
X"5c595b58",
X"83153353",
X"72802e81",
X"88387333",
X"537c732e",
X"09810680",
X"fc388114",
X"33537b73",
X"2e098106",
X"80ef3875",
X"0883c8bc",
X"082e0981",
X"0680e238",
X"80567581",
X"c42983c8",
X"cc117033",
X"831e335b",
X"57555374",
X"782e0981",
X"06973883",
X"c8d01308",
X"79082e09",
X"81068a38",
X"81143352",
X"7451fef8",
X"3f811670",
X"81ff0657",
X"538f7627",
X"c5388077",
X"08545472",
X"742e9138",
X"76518413",
X"0853722d",
X"83c08008",
X"81ff0654",
X"800b831b",
X"347353a9",
X"39811881",
X"c41681c4",
X"1681c419",
X"81c41f81",
X"c41e81c4",
X"1d6081c4",
X"05415d5e",
X"5f595656",
X"588f7825",
X"feca3880",
X"537283c0",
X"800c8e3d",
X"0d04f83d",
X"0d02ae05",
X"227d5957",
X"80568155",
X"80548653",
X"8180527a",
X"51f4ee3f",
X"83c08008",
X"81ff0683",
X"c0800c8a",
X"3d0d04f7",
X"3d0d02b2",
X"05220284",
X"05b70533",
X"605a5b57",
X"80568255",
X"79548653",
X"8180527b",
X"51f4be3f",
X"83c08008",
X"81ff0683",
X"c0800c8b",
X"3d0d04f8",
X"3d0d02af",
X"05335980",
X"58805780",
X"56805578",
X"54895380",
X"527a51f4",
X"943f83c0",
X"800881ff",
X"0683c080",
X"0c8a3d0d",
X"0483c08c",
X"080283c0",
X"8c0cfd3d",
X"0d805383",
X"c08c088c",
X"05085283",
X"c08c0888",
X"05085183",
X"d43f83c0",
X"80087083",
X"c0800c54",
X"853d0d83",
X"c08c0c04",
X"83c08c08",
X"0283c08c",
X"0cfd3d0d",
X"815383c0",
X"8c088c05",
X"085283c0",
X"8c088805",
X"085183a1",
X"3f83c080",
X"087083c0",
X"800c5485",
X"3d0d83c0",
X"8c0c0483",
X"c08c0802",
X"83c08c0c",
X"f93d0d80",
X"0b83c08c",
X"08fc050c",
X"83c08c08",
X"88050880",
X"25b93883",
X"c08c0888",
X"05083083",
X"c08c0888",
X"050c800b",
X"83c08c08",
X"f4050c83",
X"c08c08fc",
X"05088a38",
X"810b83c0",
X"8c08f405",
X"0c83c08c",
X"08f40508",
X"83c08c08",
X"fc050c83",
X"c08c088c",
X"05088025",
X"b93883c0",
X"8c088c05",
X"083083c0",
X"8c088c05",
X"0c800b83",
X"c08c08f0",
X"050c83c0",
X"8c08fc05",
X"088a3881",
X"0b83c08c",
X"08f0050c",
X"83c08c08",
X"f0050883",
X"c08c08fc",
X"050c8053",
X"83c08c08",
X"8c050852",
X"83c08c08",
X"88050851",
X"81df3f83",
X"c0800870",
X"83c08c08",
X"f8050c54",
X"83c08c08",
X"fc050880",
X"2e903883",
X"c08c08f8",
X"05083083",
X"c08c08f8",
X"050c83c0",
X"8c08f805",
X"087083c0",
X"800c5489",
X"3d0d83c0",
X"8c0c0483",
X"c08c0802",
X"83c08c0c",
X"fb3d0d80",
X"0b83c08c",
X"08fc050c",
X"83c08c08",
X"88050880",
X"25993883",
X"c08c0888",
X"05083083",
X"c08c0888",
X"050c810b",
X"83c08c08",
X"fc050c83",
X"c08c088c",
X"05088025",
X"903883c0",
X"8c088c05",
X"083083c0",
X"8c088c05",
X"0c815383",
X"c08c088c",
X"05085283",
X"c08c0888",
X"050851bd",
X"3f83c080",
X"087083c0",
X"8c08f805",
X"0c5483c0",
X"8c08fc05",
X"08802e90",
X"3883c08c",
X"08f80508",
X"3083c08c",
X"08f8050c",
X"83c08c08",
X"f8050870",
X"83c0800c",
X"54873d0d",
X"83c08c0c",
X"0483c08c",
X"080283c0",
X"8c0cfd3d",
X"0d810b83",
X"c08c08fc",
X"050c800b",
X"83c08c08",
X"f8050c83",
X"c08c088c",
X"050883c0",
X"8c088805",
X"0827b938",
X"83c08c08",
X"fc050880",
X"2eae3880",
X"0b83c08c",
X"088c0508",
X"24a23883",
X"c08c088c",
X"05081083",
X"c08c088c",
X"050c83c0",
X"8c08fc05",
X"081083c0",
X"8c08fc05",
X"0cffb839",
X"83c08c08",
X"fc050880",
X"2e80e138",
X"83c08c08",
X"8c050883",
X"c08c0888",
X"050826ad",
X"3883c08c",
X"08880508",
X"83c08c08",
X"8c050831",
X"83c08c08",
X"88050c83",
X"c08c08f8",
X"050883c0",
X"8c08fc05",
X"080783c0",
X"8c08f805",
X"0c83c08c",
X"08fc0508",
X"812a83c0",
X"8c08fc05",
X"0c83c08c",
X"088c0508",
X"812a83c0",
X"8c088c05",
X"0cff9539",
X"83c08c08",
X"90050880",
X"2e933883",
X"c08c0888",
X"05087083",
X"c08c08f4",
X"050c5191",
X"3983c08c",
X"08f80508",
X"7083c08c",
X"08f4050c",
X"5183c08c",
X"08f40508",
X"83c0800c",
X"853d0d83",
X"c08c0c04",
X"83c08c08",
X"0283c08c",
X"0cff3d0d",
X"800b83c0",
X"8c08fc05",
X"0c83c08c",
X"08880508",
X"8106ff11",
X"70097083",
X"c08c088c",
X"05080683",
X"c08c08fc",
X"05081183",
X"c08c08fc",
X"050c83c0",
X"8c088805",
X"08812a83",
X"c08c0888",
X"050c83c0",
X"8c088c05",
X"081083c0",
X"8c088c05",
X"0c515151",
X"5183c08c",
X"08880508",
X"802e8438",
X"ffab3983",
X"c08c08fc",
X"05087083",
X"c0800c51",
X"833d0d83",
X"c08c0c04",
X"fc3d0d76",
X"70797b55",
X"5555558f",
X"72278c38",
X"72750783",
X"06517080",
X"2ea938ff",
X"125271ff",
X"2e983872",
X"70810554",
X"33747081",
X"055634ff",
X"125271ff",
X"2e098106",
X"ea387483",
X"c0800c86",
X"3d0d0474",
X"51727084",
X"05540871",
X"70840553",
X"0c727084",
X"05540871",
X"70840553",
X"0c727084",
X"05540871",
X"70840553",
X"0c727084",
X"05540871",
X"70840553",
X"0cf01252",
X"718f26c9",
X"38837227",
X"95387270",
X"84055408",
X"71708405",
X"530cfc12",
X"52718326",
X"ed387054",
X"ff813900",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00002d6a",
X"00002dab",
X"00002dcb",
X"00002def",
X"00002dfb",
X"00003980",
X"0000420e",
X"000042d7",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3a00",
X"0c0c3b00",
X"0a0a0005",
X"0b0b0005",
X"07070005",
X"04044500",
X"05054400",
X"0e0f2900",
X"06060004",
X"08080004",
X"09090004",
X"080f4300",
X"090f4200",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"00005044",
X"0000534b",
X"00005157",
X"0000534b",
X"00005194",
X"000051e5",
X"00005224",
X"0000522d",
X"0000534b",
X"0000534b",
X"0000534b",
X"0000534b",
X"00005236",
X"0000523e",
X"00005245",
X"0000544b",
X"00005544",
X"00005658",
X"0000594e",
X"00005969",
X"00005955",
X"00005969",
X"00005970",
X"0000597b",
X"00005982",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"31364b00",
X"556e6b6e",
X"6f776e20",
X"74797065",
X"206f6620",
X"63617274",
X"72696467",
X"65210000",
X"41353200",
X"43415200",
X"42494e00",
X"31366b20",
X"63617274",
X"20747970",
X"65000000",
X"4c656674",
X"20666f72",
X"206f6e65",
X"20636869",
X"70000000",
X"52696768",
X"7420666f",
X"72207477",
X"6f206368",
X"69700000",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a257300",
X"45786974",
X"00000000",
X"35323030",
X"2e726f6d",
X"00000000",
X"524f4d00",
X"4d454d00",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"00000000",
X"000069b4",
X"00006804",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"35323030",
X"00000000",
X"2f617461",
X"72353230",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
