
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81e2",
X"98738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81ea",
X"a40c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757581dc",
X"c52d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7581dad9",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80e4b904",
X"fd3d0d75",
X"705254ae",
X"c33f83c0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"c0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83c0",
X"8008732e",
X"a13883c0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183c0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83c2d808",
X"248a38b5",
X"983fff0b",
X"83c2d80c",
X"800b83c0",
X"800c04ff",
X"3d0d7352",
X"83c0b408",
X"722e9b38",
X"d93f8183",
X"0b9088a0",
X"0c715196",
X"c93f8193",
X"0b9088a0",
X"0c7183c0",
X"b40c833d",
X"0d04f43d",
X"0d7e6062",
X"5c5a5580",
X"568154bc",
X"1508762e",
X"09810681",
X"92387451",
X"ffb93f79",
X"58757a25",
X"80f73883",
X"c3880870",
X"892a5783",
X"ff067884",
X"80723156",
X"56577378",
X"25833873",
X"557583c2",
X"d8082e84",
X"38fef33f",
X"83c2d808",
X"8025a638",
X"75892b51",
X"98fd3f83",
X"c388088f",
X"3dfc1155",
X"5c548152",
X"f81b5196",
X"e73f7614",
X"83c3880c",
X"7583c2d8",
X"0c745376",
X"527851b3",
X"b33f83c0",
X"800883c3",
X"88081683",
X"c3880c78",
X"7631761b",
X"5b595677",
X"8024ff8b",
X"38617a71",
X"0c547554",
X"75802e83",
X"38815473",
X"83c0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"853f7651",
X"fe993f86",
X"3dfc0553",
X"78527751",
X"968a3f79",
X"75710c54",
X"83c08008",
X"5483c080",
X"08802e83",
X"38815473",
X"83c0800c",
X"863d0d04",
X"fe3d0d75",
X"83c2d808",
X"53538072",
X"24953871",
X"732e9038",
X"80c30b90",
X"88a00c71",
X"9088a40c",
X"fdb43f80",
X"d30b9088",
X"a00c7451",
X"fdc13f80",
X"e30b9088",
X"a00c7251",
X"97b53f80",
X"f30b9088",
X"a00c83c0",
X"80085283",
X"c0800880",
X"2e833881",
X"527183c0",
X"800c843d",
X"0d04803d",
X"0d7280c0",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"3d0d72bc",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"c40b83c0",
X"800c04fd",
X"3d0d7577",
X"71547053",
X"5553a9e4",
X"3f82c813",
X"08bc150c",
X"82c01308",
X"80c0150c",
X"fcb43f73",
X"5193ab3f",
X"7383c0b4",
X"0c83c080",
X"085383c0",
X"8008802e",
X"83388153",
X"7283c080",
X"0c853d0d",
X"04fd3d0d",
X"75775553",
X"fc883f72",
X"802ea538",
X"bc130852",
X"7351a8ee",
X"3f83c080",
X"088f3877",
X"527251ff",
X"9a3f83c0",
X"8008538a",
X"3982cc13",
X"0853d839",
X"81537283",
X"c0800c85",
X"3d0d04fe",
X"3d0dff0b",
X"83c2d80c",
X"7483c0b8",
X"0c7583c2",
X"d40cafc6",
X"3f83c080",
X"0881ff06",
X"52815371",
X"993883c2",
X"f0518e94",
X"3f83c080",
X"085283c0",
X"8008802e",
X"83387252",
X"71537283",
X"c0800c84",
X"3d0d04fa",
X"3d0d787a",
X"82c41208",
X"82c41208",
X"70722459",
X"56565757",
X"73732e09",
X"81069138",
X"80c01652",
X"80c01751",
X"a6df3f83",
X"c0800855",
X"7483c080",
X"0c883d0d",
X"04f63d0d",
X"7c5b807b",
X"715c5457",
X"7a772e8c",
X"38811a82",
X"cc140854",
X"5a72f638",
X"805980d9",
X"397a5481",
X"5780707b",
X"7b315a57",
X"55ff1853",
X"74732580",
X"c13882cc",
X"14085273",
X"51ff8c3f",
X"800b83c0",
X"800825a1",
X"3882cc14",
X"0882cc11",
X"0882cc16",
X"0c7482cc",
X"120c5375",
X"802e8638",
X"7282cc17",
X"0c725480",
X"577382cc",
X"15088117",
X"575556ff",
X"b8398119",
X"59800bff",
X"1b545478",
X"73258338",
X"81547681",
X"32707506",
X"515372ff",
X"90388c3d",
X"0d04f73d",
X"0d7b7d5a",
X"5a82d052",
X"83c2d408",
X"5181c8df",
X"3f83c080",
X"0857f9aa",
X"3f795283",
X"c2dc5195",
X"b73f83c0",
X"80085480",
X"5383c080",
X"08732e09",
X"81068283",
X"3883c0b8",
X"080b0b81",
X"e7bc5370",
X"5256a69c",
X"3f0b0b81",
X"e7bc5280",
X"c01651a6",
X"8f3f75bc",
X"170c7382",
X"c0170c81",
X"0b82c417",
X"0c810b82",
X"c8170c73",
X"82cc170c",
X"ff1782d0",
X"17555781",
X"913983c0",
X"c4337082",
X"2a708106",
X"51545572",
X"81803874",
X"812a8106",
X"587780f6",
X"3874842a",
X"810682c4",
X"150c83c0",
X"c4338106",
X"82c8150c",
X"79527351",
X"a5b63f73",
X"51a5cd3f",
X"83c08008",
X"1453af73",
X"70810555",
X"3472bc15",
X"0c83c0c5",
X"527251a5",
X"973f83c0",
X"bc0882c0",
X"150c83c0",
X"d25280c0",
X"1451a584",
X"3f78802e",
X"8d387351",
X"782d83c0",
X"8008802e",
X"99387782",
X"cc150c75",
X"802e8638",
X"7382cc17",
X"0c7382d0",
X"15ff1959",
X"55567680",
X"2e9b3883",
X"c0bc5283",
X"c2dc5194",
X"ad3f83c0",
X"80088a38",
X"83c0c533",
X"5372fed2",
X"3878802e",
X"893883c0",
X"b80851fc",
X"b83f83c0",
X"b8085372",
X"83c0800c",
X"8b3d0d04",
X"ff3d0d80",
X"527351fd",
X"b53f833d",
X"0d04f03d",
X"0d627052",
X"54f5d93f",
X"83c08008",
X"7453873d",
X"70535555",
X"f5f93ff6",
X"d93f7351",
X"d33f6353",
X"745283c0",
X"800851fa",
X"b83f923d",
X"0d047183",
X"c0800c04",
X"80c01283",
X"c0800c04",
X"803d0d72",
X"82c01108",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"7282cc11",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d7282c4",
X"110883c0",
X"800c5182",
X"3d0d04f9",
X"3d0d7983",
X"c0900857",
X"57817727",
X"81963876",
X"88170827",
X"818e3875",
X"33557482",
X"2e893874",
X"832eb338",
X"80fe3974",
X"54761083",
X"fe065376",
X"882a8c17",
X"08055289",
X"3dfc0551",
X"a9f43f83",
X"c0800880",
X"df38029d",
X"0533893d",
X"3371882b",
X"07565680",
X"d1398454",
X"76822b83",
X"fc065376",
X"872a8c17",
X"08055289",
X"3dfc0551",
X"a9c43f83",
X"c08008b0",
X"38029f05",
X"33028405",
X"9e053371",
X"982b7190",
X"2b07028c",
X"059d0533",
X"70882b72",
X"078d3d33",
X"7180ffff",
X"fe800607",
X"51525357",
X"58568339",
X"81557483",
X"c0800c89",
X"3d0d04fb",
X"3d0d83c0",
X"9008fe19",
X"881208fe",
X"05555654",
X"80567473",
X"278d3882",
X"14337571",
X"29941608",
X"05575375",
X"83c0800c",
X"873d0d04",
X"fc3d0d76",
X"52800b83",
X"c0900870",
X"33515253",
X"70832e09",
X"81069138",
X"95123394",
X"13337198",
X"2b71902b",
X"07555551",
X"9b12339a",
X"13337188",
X"2b077407",
X"83c0800c",
X"55863d0d",
X"04fc3d0d",
X"7683c090",
X"08555580",
X"75238815",
X"08537281",
X"2e883888",
X"14087326",
X"85388152",
X"b2397290",
X"38733352",
X"71832e09",
X"81068538",
X"90140853",
X"728c160c",
X"72802e8d",
X"387251fe",
X"d63f83c0",
X"80085285",
X"39901408",
X"52719016",
X"0c805271",
X"83c0800c",
X"863d0d04",
X"fa3d0d78",
X"83c09008",
X"71228105",
X"7083ffff",
X"06575457",
X"5573802e",
X"88389015",
X"08537286",
X"38835280",
X"e739738f",
X"06527180",
X"da388113",
X"90160c8c",
X"15085372",
X"9038830b",
X"84172257",
X"52737627",
X"80c638bf",
X"39821633",
X"ff057484",
X"2a065271",
X"b2387251",
X"fcb13f81",
X"527183c0",
X"800827a8",
X"38835283",
X"c0800888",
X"1708279c",
X"3883c080",
X"088c160c",
X"83c08008",
X"51fdbc3f",
X"83c08008",
X"90160c73",
X"75238052",
X"7183c080",
X"0c883d0d",
X"04f23d0d",
X"60626458",
X"5e5b7533",
X"5574a02e",
X"09810688",
X"38811670",
X"4456ef39",
X"62703356",
X"5674af2e",
X"09810684",
X"38811643",
X"800b881c",
X"0c627033",
X"5155749f",
X"2691387a",
X"51fdd23f",
X"83c08008",
X"56807d34",
X"83813993",
X"3d841c08",
X"7058595f",
X"8a55a076",
X"70810558",
X"34ff1555",
X"74ff2e09",
X"8106ef38",
X"80705a5c",
X"887f085f",
X"5a7b811d",
X"7081ff06",
X"60137033",
X"70af3270",
X"30a07327",
X"71802507",
X"5151525b",
X"535e5755",
X"7480e738",
X"76ae2e09",
X"81068338",
X"8155787a",
X"27750755",
X"74802e9f",
X"38798832",
X"703078ae",
X"32703070",
X"73079f2a",
X"53515751",
X"5675bb38",
X"88598b5a",
X"ffab3976",
X"982b5574",
X"80258738",
X"81e1a817",
X"3357ff9f",
X"17557499",
X"268938e0",
X"177081ff",
X"06585578",
X"811a7081",
X"ff06721b",
X"535b5755",
X"767534fe",
X"f8397b1e",
X"7f0c8055",
X"76a02683",
X"38815574",
X"8b19347a",
X"51fc823f",
X"83c08008",
X"80f538a0",
X"547a2270",
X"852b83e0",
X"06545590",
X"1b08527c",
X"51a3ff3f",
X"83c08008",
X"5783c080",
X"08818138",
X"7c335574",
X"802e80f4",
X"388b1d33",
X"70832a70",
X"81065156",
X"5674b438",
X"8b7d841d",
X"0883c080",
X"08595b5b",
X"58ff1858",
X"77ff2e9a",
X"38797081",
X"055b3379",
X"7081055b",
X"33717131",
X"52565675",
X"802ee238",
X"86397580",
X"2e96387a",
X"51fbe53f",
X"ff863983",
X"c0800856",
X"83c08008",
X"b6388339",
X"7656841b",
X"088b1133",
X"515574a7",
X"388b1d33",
X"70842a70",
X"81065156",
X"56748938",
X"83569439",
X"81569039",
X"7c51fa94",
X"3f83c080",
X"08881c0c",
X"fd813975",
X"83c0800c",
X"903d0d04",
X"f83d0d7a",
X"7c595782",
X"5483fe53",
X"77527651",
X"a2c43f83",
X"5683c080",
X"0880ec38",
X"81173377",
X"3371882b",
X"07565682",
X"567482d4",
X"d52e0981",
X"0680d438",
X"7554b653",
X"77527651",
X"a2983f83",
X"c0800898",
X"38811733",
X"77337188",
X"2b0783c0",
X"80085256",
X"56748182",
X"c62eac38",
X"825480d2",
X"53775276",
X"51a1ef3f",
X"83c08008",
X"98388117",
X"33773371",
X"882b0783",
X"c0800852",
X"56567481",
X"82c62e83",
X"38815675",
X"83c0800c",
X"8a3d0d04",
X"eb3d0d67",
X"5a800b83",
X"c0900ca1",
X"913f83c0",
X"80088106",
X"55825674",
X"83ef3874",
X"75538f3d",
X"70535759",
X"feca3f83",
X"c0800881",
X"ff065776",
X"812e0981",
X"0680d438",
X"905483be",
X"53745275",
X"51a1833f",
X"83c08008",
X"80c9388f",
X"3d335574",
X"802e80c9",
X"3802bf05",
X"33028405",
X"be053371",
X"982b7190",
X"2b07028c",
X"05bd0533",
X"70882b72",
X"07953d33",
X"71077058",
X"7b575e52",
X"5e575957",
X"fdee3f83",
X"c0800881",
X"ff065776",
X"832e0981",
X"06863881",
X"5682f239",
X"76802e86",
X"38865682",
X"e839a454",
X"8d537852",
X"7551a09a",
X"3f815683",
X"c0800882",
X"d43802be",
X"05330284",
X"05bd0533",
X"71882b07",
X"595d77ab",
X"380280ce",
X"05330284",
X"0580cd05",
X"3371982b",
X"71902b07",
X"973d3370",
X"882b7207",
X"02940580",
X"cb053371",
X"0754525e",
X"57595602",
X"b7053378",
X"71290288",
X"05b60533",
X"028c05b5",
X"05337188",
X"2b07701d",
X"707f8c05",
X"0c5f5957",
X"595d8e3d",
X"33821b34",
X"02b90533",
X"903d3371",
X"882b075a",
X"5c78841b",
X"2302bb05",
X"33028405",
X"ba053371",
X"882b0756",
X"5c74ab38",
X"0280ca05",
X"33028405",
X"80c90533",
X"71982b71",
X"902b0796",
X"3d337088",
X"2b720702",
X"940580c7",
X"05337107",
X"51525357",
X"5e5c7476",
X"31783179",
X"842a903d",
X"33547171",
X"31535656",
X"81b9c43f",
X"83c08008",
X"82057088",
X"1c0c83c0",
X"8008e08a",
X"05565674",
X"83dffe26",
X"83388257",
X"83fff676",
X"27853883",
X"57893986",
X"5676802e",
X"80db3876",
X"7a347683",
X"2e098106",
X"b0380280",
X"d6053302",
X"840580d5",
X"05337198",
X"2b71902b",
X"07993d33",
X"70882b72",
X"07029405",
X"80d30533",
X"71077f90",
X"050c525e",
X"57585686",
X"39771b90",
X"1b0c841a",
X"228c1b08",
X"1971842a",
X"05941c0c",
X"5d800b81",
X"1b347983",
X"c0900c80",
X"567583c0",
X"800c973d",
X"0d04e93d",
X"0d83c090",
X"08568554",
X"75802e81",
X"8238800b",
X"81173499",
X"3de01146",
X"6a548a3d",
X"705458ec",
X"0551f6e5",
X"3f83c080",
X"085483c0",
X"800880df",
X"38893d33",
X"5473802e",
X"913802ab",
X"05337084",
X"2a810651",
X"5574802e",
X"86388354",
X"80c13976",
X"51f4893f",
X"83c08008",
X"a0170c02",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"9c1c0c52",
X"78981b0c",
X"53565957",
X"810b8117",
X"34745473",
X"83c0800c",
X"993d0d04",
X"f53d0d7d",
X"7f617283",
X"c090085a",
X"5d5d595c",
X"807b0c85",
X"5775802e",
X"81e03881",
X"16338106",
X"55845774",
X"802e81d2",
X"38913974",
X"81173486",
X"39800b81",
X"17348157",
X"81c0399c",
X"16089817",
X"08315574",
X"78278338",
X"74587780",
X"2e81a938",
X"98160870",
X"83ff0656",
X"577480cf",
X"38821633",
X"ff057789",
X"2a067081",
X"ff065a55",
X"78a03876",
X"8738a016",
X"08558d39",
X"a4160851",
X"f0e93f83",
X"c0800855",
X"817527ff",
X"a83874a4",
X"170ca416",
X"0851f283",
X"3f83c080",
X"085583c0",
X"8008802e",
X"ff893883",
X"c0800819",
X"a8170c98",
X"160883ff",
X"06848071",
X"31515577",
X"75278338",
X"77557483",
X"ffff0654",
X"98160883",
X"ff0653a8",
X"16085279",
X"577b8338",
X"7b577651",
X"9ac03f83",
X"c08008fe",
X"d0389816",
X"08159817",
X"0c741a78",
X"76317c08",
X"177d0c59",
X"5afed339",
X"80577683",
X"c0800c8d",
X"3d0d04fa",
X"3d0d7883",
X"c0900855",
X"56855573",
X"802e81e3",
X"38811433",
X"81065384",
X"5572802e",
X"81d5389c",
X"14085372",
X"76278338",
X"72569814",
X"0857800b",
X"98150c75",
X"802e81b9",
X"38821433",
X"70892b56",
X"5376802e",
X"b7387452",
X"ff165181",
X"b4c53f83",
X"c08008ff",
X"18765470",
X"53585381",
X"b4b53f83",
X"c0800873",
X"26963874",
X"30707806",
X"7098170c",
X"777131a4",
X"17085258",
X"51538939",
X"a0140870",
X"a4160c53",
X"747627b9",
X"387251ee",
X"d63f83c0",
X"80085381",
X"0b83c080",
X"08278b38",
X"88140883",
X"c0800826",
X"8838800b",
X"811534b0",
X"3983c080",
X"08a4150c",
X"98140815",
X"98150c75",
X"753156c4",
X"39981408",
X"16709816",
X"0c735256",
X"efc53f83",
X"c080088c",
X"3883c080",
X"08811534",
X"81559439",
X"821433ff",
X"0576892a",
X"0683c080",
X"0805a815",
X"0c805574",
X"83c0800c",
X"883d0d04",
X"ef3d0d63",
X"56855583",
X"c0900880",
X"2e80d238",
X"933df405",
X"84170c64",
X"53883d70",
X"53765257",
X"f1cf3f83",
X"c0800855",
X"83c08008",
X"b438883d",
X"33547380",
X"2ea13802",
X"a7053370",
X"842a7081",
X"06515555",
X"83557380",
X"2e973876",
X"51eef53f",
X"83c08008",
X"88170c75",
X"51efa63f",
X"83c08008",
X"557483c0",
X"800c933d",
X"0d04e43d",
X"0d6ea13d",
X"08405e85",
X"5683c090",
X"08802e84",
X"85389e3d",
X"f405841f",
X"0c7e9838",
X"7d51eef5",
X"3f83c080",
X"085683ee",
X"39814181",
X"f6398341",
X"81f13993",
X"3d7f9605",
X"4159807f",
X"8295055e",
X"56756081",
X"ff053483",
X"41901e08",
X"762e81d3",
X"38a0547d",
X"2270852b",
X"83e00654",
X"58901e08",
X"52785196",
X"c93f83c0",
X"80084183",
X"c08008ff",
X"b8387833",
X"5c7b802e",
X"ffb4388b",
X"193370bf",
X"06718106",
X"52435574",
X"802e80de",
X"387b81bf",
X"0655748f",
X"2480d338",
X"9a193355",
X"7480cb38",
X"f31d7058",
X"5d815675",
X"8b2e0981",
X"0685388e",
X"568b3975",
X"9a2e0981",
X"0683389c",
X"56751970",
X"70810552",
X"33713381",
X"1a821a5f",
X"5b525b55",
X"74863879",
X"77348539",
X"80df7734",
X"777b5757",
X"7aa02e09",
X"8106c038",
X"81567b81",
X"e5327030",
X"709f2a51",
X"51557bae",
X"2e933874",
X"802e8e38",
X"61832a70",
X"81065155",
X"74802e97",
X"387d51ed",
X"df3f83c0",
X"80084183",
X"c0800887",
X"38901e08",
X"feaf3880",
X"60347580",
X"2e88387c",
X"527f518d",
X"eb3f6080",
X"2e863880",
X"0b901f0c",
X"60566083",
X"2e853860",
X"81d03889",
X"1f57901e",
X"08802e81",
X"a8388056",
X"75197033",
X"515574a0",
X"2ea03874",
X"852e0981",
X"06843881",
X"e5557477",
X"70810559",
X"34811670",
X"81ff0657",
X"55877627",
X"d7388819",
X"335574a0",
X"2ea938ae",
X"77708105",
X"59348856",
X"75197033",
X"515574a0",
X"2e953874",
X"77708105",
X"59348116",
X"7081ff06",
X"57558a76",
X"27e2388b",
X"19337f88",
X"05349f19",
X"339e1a33",
X"71982b71",
X"902b079d",
X"1c337088",
X"2b72079c",
X"1e337107",
X"640c5299",
X"1d33981e",
X"3371882b",
X"07535153",
X"57595674",
X"7f840523",
X"97193396",
X"1a337188",
X"2b075656",
X"747f8605",
X"23807734",
X"7d51ebf0",
X"3f83c080",
X"08833270",
X"30707207",
X"9f2c83c0",
X"80080652",
X"5656961f",
X"3355748a",
X"38891f52",
X"961f518b",
X"f73f7583",
X"c0800c9e",
X"3d0d04f4",
X"3d0d7e8f",
X"3dec1156",
X"56589053",
X"f0155277",
X"51e0b13f",
X"83c08008",
X"80d63878",
X"902e0981",
X"0680cd38",
X"02ab0533",
X"81eaac0b",
X"81eaac33",
X"5758568c",
X"3974762e",
X"8a388417",
X"70335657",
X"74f33876",
X"33705755",
X"74802eac",
X"38821722",
X"708a2b90",
X"3dec0556",
X"70555656",
X"96800a52",
X"7751dfe0",
X"3f83c080",
X"08863878",
X"752e8538",
X"80568539",
X"81173356",
X"7583c080",
X"0c8e3d0d",
X"04fc3d0d",
X"76705255",
X"8afe3f83",
X"c0800815",
X"ff055473",
X"752e8e38",
X"73335372",
X"ae2e8638",
X"ff1454ef",
X"39775281",
X"14518a96",
X"3f83c080",
X"08307083",
X"c0800807",
X"802583c0",
X"800c5386",
X"3d0d04fa",
X"3d0d7857",
X"80775256",
X"e6c23f83",
X"c0800883",
X"c0800833",
X"53547176",
X"2e80c738",
X"733383c0",
X"94173356",
X"53749138",
X"765183c3",
X"ac085271",
X"2d83c080",
X"0852ad39",
X"ff9f1352",
X"71992689",
X"38e01370",
X"81ff0654",
X"52747332",
X"70307072",
X"07802578",
X"05811770",
X"33545758",
X"545271ff",
X"bb388052",
X"7183c080",
X"0c883d0d",
X"04fc3d0d",
X"76705255",
X"e6803f83",
X"c0800854",
X"815383c0",
X"800880d0",
X"387451e5",
X"c33f83c0",
X"800881e7",
X"cc5383c0",
X"80085253",
X"fea33f83",
X"c08008b0",
X"3881e7d0",
X"527251fe",
X"943f83c0",
X"8008a138",
X"81e7d452",
X"7251fe85",
X"3f83c080",
X"08923881",
X"e7d85272",
X"51fdf63f",
X"83c08008",
X"802e8338",
X"81547353",
X"7283c080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"e5903f81",
X"5383c080",
X"08983873",
X"51e4d93f",
X"83c3a008",
X"5283c080",
X"0851fdbd",
X"3f83c080",
X"08537283",
X"c0800c85",
X"3d0d04dd",
X"3d0da63d",
X"085f800b",
X"81eba033",
X"555b737b",
X"2e85cc38",
X"86537a52",
X"83c09451",
X"a1cd3f7e",
X"51daae3f",
X"83c08008",
X"33973d56",
X"54737b2e",
X"09810696",
X"3881ebcc",
X"52745187",
X"db3f9a39",
X"7e527851",
X"dde13f85",
X"96397e51",
X"da8f3f83",
X"c0800852",
X"7451d9bf",
X"3f804480",
X"43804280",
X"41adbb52",
X"963d7052",
X"5ee0cb3f",
X"83c08008",
X"59800b83",
X"c0800855",
X"5c83c080",
X"087c2e94",
X"38811c74",
X"525ce3cd",
X"3f83c080",
X"085483c0",
X"8008ee38",
X"805aff40",
X"7909709f",
X"2c7b065b",
X"547b7a24",
X"8438ff1c",
X"5af61a70",
X"09709f2c",
X"72067bff",
X"125a5a52",
X"55558075",
X"25953876",
X"51e3923f",
X"83c08008",
X"76ff1858",
X"55577380",
X"24ed3874",
X"602e8638",
X"a2833f74",
X"4078ff1b",
X"70585e58",
X"807a2595",
X"387751e2",
X"e83f83c0",
X"800876ff",
X"18585558",
X"738024ed",
X"38800b83",
X"c7dc0c81",
X"800b83c8",
X"940c81e7",
X"dc518bdf",
X"3f800b83",
X"c8940c83",
X"c0945281",
X"e7e4518b",
X"ce3fa80b",
X"83c7dc0c",
X"76802e80",
X"e43883c7",
X"dc087779",
X"32703070",
X"72078025",
X"70872b83",
X"c8940c51",
X"56785356",
X"56e29b3f",
X"83c08008",
X"802e8838",
X"81e7f051",
X"8b953f76",
X"51e1dd3f",
X"83c08008",
X"5281e9c4",
X"518b843f",
X"7651e1e5",
X"3f83c080",
X"0883c7dc",
X"08555775",
X"74258638",
X"a81656f7",
X"397583c7",
X"dc0c86f0",
X"7624ff98",
X"3887980b",
X"83c7dc0c",
X"77802ea9",
X"387751e1",
X"9b3f83c0",
X"80087852",
X"55e1bb3f",
X"81e7f854",
X"83c08008",
X"853881e7",
X"f4547453",
X"735281e7",
X"c0518aab",
X"3f805481",
X"e7c8518a",
X"a23f8114",
X"5473a82e",
X"098106ef",
X"38868da0",
X"519dfb3f",
X"8052913d",
X"705257b6",
X"a93f8352",
X"7651b6a2",
X"3f645473",
X"ff2e0981",
X"069738ff",
X"1b700970",
X"9f2c7206",
X"52555b80",
X"0b83c094",
X"1c3481c2",
X"39807425",
X"ab387a85",
X"2e098106",
X"91388653",
X"805283c0",
X"94519dc3",
X"3f805b81",
X"a5397383",
X"c0941c34",
X"811b5b81",
X"99398076",
X"34819339",
X"63818f38",
X"62802e80",
X"fb387c54",
X"73ff2e96",
X"3878802e",
X"81893878",
X"51dffa3f",
X"83c08008",
X"ff155559",
X"e7397880",
X"2e80f438",
X"7851dff6",
X"3f83c080",
X"08802efb",
X"c7387851",
X"dfbe3f83",
X"c0800852",
X"81e7bc51",
X"81e73f83",
X"c08008a3",
X"387d5183",
X"9f3f83c0",
X"80085574",
X"ff165654",
X"807425ae",
X"38741e70",
X"33555673",
X"af2eff8a",
X"38e93978",
X"51deff3f",
X"83c08008",
X"527d5182",
X"d73f8f39",
X"60882961",
X"10057a05",
X"62055afb",
X"c7396380",
X"2efb8a38",
X"80527651",
X"b4b43fa5",
X"3d0d04ff",
X"3d0d028f",
X"05337010",
X"81059088",
X"900c5283",
X"3d0d04ff",
X"3d0d028f",
X"05335290",
X"88840870",
X"892a7081",
X"06515151",
X"70802e86",
X"38aced3f",
X"ea397190",
X"88800c83",
X"3d0d0480",
X"3d0d9088",
X"8c087088",
X"2a708106",
X"51515170",
X"802e8638",
X"acca3fea",
X"39908888",
X"0883c080",
X"0c823d0d",
X"04908894",
X"0883c080",
X"0c04fd3d",
X"0d757754",
X"54807325",
X"94387370",
X"81055533",
X"5281e7fc",
X"5187883f",
X"ff1353e9",
X"39853d0d",
X"04fd3d0d",
X"75775354",
X"73335170",
X"89387133",
X"5170802e",
X"a1387333",
X"72335253",
X"72712785",
X"38ff5194",
X"39707327",
X"85388151",
X"8b398114",
X"81135354",
X"d3398051",
X"7083c080",
X"0c853d0d",
X"04fd3d0d",
X"75775454",
X"72337081",
X"ff065252",
X"70802ea3",
X"387181ff",
X"068114ff",
X"bf125354",
X"52709926",
X"8938a012",
X"7081ff06",
X"53517174",
X"70810556",
X"34d23980",
X"7434853d",
X"0d04ffbd",
X"3d0d80c6",
X"3d0852a5",
X"3d705254",
X"ffb33f80",
X"c73d0852",
X"853d7052",
X"53ffa63f",
X"72527351",
X"fedf3f80",
X"c53d0d04",
X"fe3d0d74",
X"76535371",
X"70810553",
X"33517073",
X"70810555",
X"3470f038",
X"843d0d04",
X"fe3d0d74",
X"52807233",
X"52537073",
X"2e8d3881",
X"12811471",
X"33535452",
X"70f53872",
X"83c0800c",
X"843d0d04",
X"f63d0d7c",
X"7e60625a",
X"5d5b5680",
X"59815585",
X"39747a29",
X"55745275",
X"5181a1b3",
X"3f83c080",
X"087a27ed",
X"3874802e",
X"80e03874",
X"52755181",
X"a19d3f83",
X"c0800875",
X"53765254",
X"81a1c33f",
X"83c08008",
X"7a537552",
X"5681a183",
X"3f83c080",
X"08793070",
X"7b079f2a",
X"70778024",
X"07515154",
X"55728738",
X"83c08008",
X"c2387681",
X"18b01655",
X"58588974",
X"258b38b7",
X"14537a85",
X"3880d714",
X"53727834",
X"811959ff",
X"9c398077",
X"348c3d0d",
X"04f73d0d",
X"7b7d7f62",
X"029005bb",
X"05335759",
X"565a5ab0",
X"58728338",
X"a0587570",
X"70810552",
X"33715954",
X"55903980",
X"74258e38",
X"ff147770",
X"81055933",
X"545472ef",
X"3873ff15",
X"55538073",
X"25893877",
X"52795178",
X"2def3975",
X"33755753",
X"72802e90",
X"38725279",
X"51782d75",
X"70810557",
X"3353ed39",
X"8b3d0d04",
X"ee3d0d64",
X"66696970",
X"70810552",
X"335b4a5c",
X"5e5e7680",
X"2e82f938",
X"76a52e09",
X"810682e0",
X"38807041",
X"67707081",
X"05523371",
X"4a59575f",
X"76b02e09",
X"81068c38",
X"75708105",
X"57337648",
X"57815fd0",
X"17567589",
X"2680da38",
X"76675c59",
X"805c9339",
X"778a2480",
X"c3387b8a",
X"29187b70",
X"81055d33",
X"5a5cd019",
X"7081ff06",
X"58588977",
X"27a438ff",
X"9f197081",
X"ff06ffa9",
X"1b5a5156",
X"85762792",
X"38ffbf19",
X"7081ff06",
X"51567585",
X"268a38c9",
X"19587780",
X"25ffb938",
X"7a477b40",
X"7881ff06",
X"577680e4",
X"2e80e538",
X"7680e424",
X"a7387680",
X"d82e8186",
X"387680d8",
X"24903876",
X"802e81cc",
X"3876a52e",
X"81b63881",
X"b9397680",
X"e32e818c",
X"3881af39",
X"7680f52e",
X"9b387680",
X"f5248b38",
X"7680f32e",
X"81813881",
X"99397680",
X"f82e80ca",
X"38818f39",
X"913d7055",
X"5780538a",
X"5279841b",
X"7108535b",
X"56fbfd3f",
X"7655ab39",
X"79841b71",
X"08943d70",
X"5b5b525b",
X"56758025",
X"8c387530",
X"56ad7834",
X"0280c105",
X"57765480",
X"538a5275",
X"51fbd13f",
X"77557e54",
X"b839913d",
X"70557780",
X"d8327030",
X"70802556",
X"51585690",
X"5279841b",
X"7108535b",
X"57fbad3f",
X"7555db39",
X"79841b83",
X"1233545b",
X"56983979",
X"841b7108",
X"575b5680",
X"547f537c",
X"527d51fc",
X"9c3f8739",
X"76527d51",
X"7c2d6670",
X"33588105",
X"47fd8339",
X"943d0d04",
X"7283c09c",
X"0c7183c0",
X"a00c04fb",
X"3d0d883d",
X"70708405",
X"52085754",
X"755383c0",
X"9c085283",
X"c0a00851",
X"fcc63f87",
X"3d0d04ff",
X"3d0d7370",
X"08535102",
X"93053372",
X"34700881",
X"05710c83",
X"3d0d04fc",
X"3d0d873d",
X"88115578",
X"54bddb53",
X"51fc993f",
X"8052873d",
X"51d13f86",
X"3d0d04fc",
X"3d0d7655",
X"7483c3b8",
X"082eaf38",
X"80537451",
X"87cc3f83",
X"c0800881",
X"ff06ff14",
X"7081ff06",
X"7230709f",
X"2a515255",
X"53547280",
X"2e843871",
X"dd3873fe",
X"387483c3",
X"b80c863d",
X"0d04ff3d",
X"0dff0b83",
X"c3b80c84",
X"b43f8151",
X"87903f83",
X"c0800881",
X"ff065271",
X"ee3881d4",
X"3f7183c0",
X"800c833d",
X"0d04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"823f7280",
X"2ea03883",
X"c3cc1433",
X"75708105",
X"57348114",
X"7083ffff",
X"06ff1570",
X"83ffff06",
X"56525552",
X"dd39800b",
X"83c0800c",
X"863d0d04",
X"fc3d0d76",
X"787a1156",
X"53558053",
X"71742e93",
X"38721551",
X"703383c3",
X"cc133481",
X"12811454",
X"52ea3980",
X"0b83c080",
X"0c863d0d",
X"04fd3d0d",
X"905483c3",
X"b8085186",
X"fd3f83c0",
X"800881ff",
X"06ff1571",
X"30713070",
X"73079f2a",
X"729f2a06",
X"52555255",
X"5372db38",
X"853d0d04",
X"803d0d83",
X"c3c40883",
X"2b83c3c0",
X"08079080",
X"a80c823d",
X"0d04800b",
X"83c3c40c",
X"e33f0481",
X"0b83c3c4",
X"0cda3f04",
X"ed3f0471",
X"83c3bc0c",
X"04803d0d",
X"8051f43f",
X"810b83c3",
X"c40c860b",
X"83c3c00c",
X"ffba3f82",
X"3d0d0484",
X"0b83c3c0",
X"0cffad3f",
X"04860b83",
X"c3c00cff",
X"a33f0483",
X"0b83c3c0",
X"0cff993f",
X"04870b83",
X"c3c00cff",
X"8f3f0480",
X"3d0d028b",
X"05339080",
X"a40c9080",
X"a8087081",
X"06515170",
X"f5389080",
X"a4087081",
X"ff0683c0",
X"800c5182",
X"3d0d0480",
X"3d0d81ff",
X"51d13f83",
X"c0800881",
X"ff0683c0",
X"800c823d",
X"0d04803d",
X"0d73902b",
X"73079080",
X"b40c823d",
X"0d0404fb",
X"3d0d7802",
X"84059f05",
X"3370982b",
X"55575572",
X"80259b38",
X"7580ff06",
X"56805280",
X"f751e03f",
X"83c08008",
X"81ff0654",
X"73812680",
X"fb38fee1",
X"3fffa43f",
X"fed13fff",
X"9e3f7551",
X"fef13f74",
X"982a51fe",
X"ea3f7490",
X"2a7081ff",
X"065253fe",
X"de3f7488",
X"2a7081ff",
X"065253fe",
X"d23f7481",
X"ff0651fe",
X"ca3f8155",
X"7580c02e",
X"09810686",
X"38819555",
X"8d397580",
X"c82e0981",
X"06843881",
X"87557451",
X"fea93f8a",
X"55fecc3f",
X"83c08008",
X"81ff0670",
X"982b5454",
X"7280258c",
X"38ff1570",
X"81ff0656",
X"5374e238",
X"7383c080",
X"0c873d0d",
X"04fa3d0d",
X"fdb73ffd",
X"d83f8a54",
X"fe993fff",
X"147081ff",
X"06555373",
X"f3387374",
X"535580c0",
X"51feac3f",
X"83c08008",
X"81ff0654",
X"73812e09",
X"8106829f",
X"3883aa52",
X"80c851fe",
X"923f83c0",
X"800881ff",
X"06537281",
X"2e098106",
X"81a83874",
X"54873d74",
X"115456fd",
X"ce3f83c0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e5",
X"38029a05",
X"33537281",
X"2e098106",
X"81d93802",
X"9b053353",
X"80ce9054",
X"7281aa2e",
X"8d3881c7",
X"3980e451",
X"8d883fff",
X"14547380",
X"2e81b838",
X"820a5281",
X"e951fdab",
X"3f83c080",
X"0881ff06",
X"5372de38",
X"725280fa",
X"51fd983f",
X"83c08008",
X"81ff0653",
X"72819038",
X"72547316",
X"53fcdc3f",
X"83c08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e83887",
X"3d337086",
X"2a708106",
X"5154548c",
X"557280e3",
X"38845580",
X"de397452",
X"81e951fc",
X"d23f83c0",
X"800881ff",
X"06538255",
X"81e95681",
X"73278638",
X"735580c1",
X"5680ce90",
X"548a3980",
X"e4518bfa",
X"3fff1454",
X"73802ea9",
X"38805275",
X"51fca03f",
X"83c08008",
X"81ff0653",
X"72e13884",
X"805280d0",
X"51fc8c3f",
X"83c08008",
X"81ff0653",
X"72802e83",
X"38805574",
X"83c3c834",
X"fb873ffb",
X"ca3f883d",
X"0d04fb3d",
X"0d775480",
X"0b83c3c8",
X"3370832a",
X"70810651",
X"55575572",
X"752e0981",
X"06853873",
X"892b5473",
X"5280d151",
X"fbc53f83",
X"c0800881",
X"ff065372",
X"bd3882b8",
X"c054fb8b",
X"3f83c080",
X"0881ff06",
X"537281ff",
X"2e098106",
X"8938ff14",
X"5473e738",
X"9f397281",
X"fe2e0981",
X"06963883",
X"c7cc5283",
X"c3cc51fa",
X"f53ffadb",
X"3ffad83f",
X"83398155",
X"fa8b3ffa",
X"ce3f7481",
X"ff0683c0",
X"800c873d",
X"0d04fb3d",
X"0d7783c3",
X"cc5654f9",
X"e63f83c3",
X"c8337083",
X"2a708106",
X"51545672",
X"85387389",
X"2b547352",
X"80d851fa",
X"c23f83c0",
X"800881ff",
X"06537280",
X"e23881ff",
X"51f9e03f",
X"81fe51f9",
X"da3f8480",
X"53747081",
X"05563351",
X"f9cd3fff",
X"137083ff",
X"ff065153",
X"72eb3872",
X"51f9bc3f",
X"7251f9b7",
X"3ff9dc3f",
X"83c08008",
X"9f0653a7",
X"88547285",
X"2e8c3899",
X"3980e451",
X"89b83fff",
X"1454f9bf",
X"3f83c080",
X"0881ff2e",
X"843873e9",
X"38f8ea3f",
X"f9ad3f80",
X"0b83c080",
X"0c873d0d",
X"047183c7",
X"d00c8880",
X"800b83c7",
X"cc0c8480",
X"800b83c7",
X"d40c04f0",
X"3d0d8380",
X"805683c7",
X"d0081683",
X"c7cc0817",
X"56547433",
X"743483c7",
X"d4081654",
X"80743481",
X"16567583",
X"80a02e09",
X"8106db38",
X"83d08056",
X"83c7d008",
X"1683c7cc",
X"08175654",
X"74337434",
X"83c7d408",
X"16548074",
X"34811656",
X"7583d090",
X"2e098106",
X"db3883a8",
X"805683c7",
X"d0081683",
X"c7cc0817",
X"56547433",
X"743483c7",
X"d4081654",
X"80743481",
X"16567583",
X"a8902e09",
X"8106db38",
X"805683c7",
X"d0081683",
X"c7d40817",
X"55557333",
X"75348116",
X"56758180",
X"802e0981",
X"06e43889",
X"e03f893d",
X"58a25381",
X"e3a85277",
X"518197a2",
X"3f80578c",
X"805683c7",
X"d4081677",
X"19555573",
X"33753481",
X"16811858",
X"5676a22e",
X"098106e6",
X"38860b87",
X"a8833480",
X"0b87a882",
X"34800b87",
X"809a34af",
X"0b878096",
X"34bf0b87",
X"80973480",
X"0b878098",
X"349f0b87",
X"80993480",
X"0b87809b",
X"34f80b87",
X"a8893476",
X"87a88034",
X"820b87d0",
X"8f34820b",
X"87a88134",
X"840b8780",
X"9f34ff0b",
X"87d08b34",
X"923d0d04",
X"fe3d0d80",
X"5383c7d4",
X"081383c7",
X"d0081452",
X"52703372",
X"34811353",
X"72818080",
X"2e098106",
X"e4388380",
X"805383c7",
X"d4081383",
X"c7d00814",
X"52527033",
X"72348113",
X"53728380",
X"a02e0981",
X"06e43883",
X"d0805383",
X"c7d40813",
X"83c7d008",
X"14525270",
X"33723481",
X"13537283",
X"d0902e09",
X"8106e438",
X"83a88053",
X"83c7d408",
X"1383c7d0",
X"08145252",
X"70337234",
X"81135372",
X"83a8902e",
X"098106e4",
X"38843d0d",
X"04803d0d",
X"90809008",
X"810683c0",
X"800c823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087081",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fd0676",
X"1007720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870822c",
X"bf0683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe830676",
X"822b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087088",
X"2c870683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f1ff06",
X"76882b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"8b2c8106",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870efff",
X"06768b2b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70912cbf",
X"0683c080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870fc",
X"87ffff06",
X"76912b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"992c8106",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870ffbf",
X"0a067699",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"08709a2c",
X"830683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"cf0a0676",
X"9a2b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"9008709c",
X"2c870683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f10a06",
X"769c2b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80bc0887",
X"0683c080",
X"0c823d0d",
X"04ff3d0d",
X"9080bc70",
X"0870f806",
X"7607720c",
X"5252833d",
X"0d04803d",
X"0d9080bc",
X"0870842c",
X"810683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"bc700870",
X"ef067684",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d9080bc",
X"0870852c",
X"810683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"bc700870",
X"df067685",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d9080bc",
X"0870862c",
X"810683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"bc700870",
X"ffbf0676",
X"862b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"80087088",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"892c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708a2c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708b2c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708c",
X"2cbf0683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"922c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"70932c81",
X"0683c080",
X"0c51823d",
X"0d04fe3d",
X"0d7481e6",
X"29872a90",
X"80a00c84",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70810554",
X"34ff1151",
X"f039843d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"8405540c",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"81808053",
X"80528880",
X"0a51ffb3",
X"3fa08053",
X"80528280",
X"0a51c73f",
X"843d0d04",
X"803d0d81",
X"51f9cf3f",
X"72802e90",
X"388051fb",
X"d03fce3f",
X"81eba433",
X"51fbc63f",
X"8151f9e0",
X"3f8051f9",
X"db3f8051",
X"f9ac3f82",
X"3d0d04fd",
X"3d0d7552",
X"805480ff",
X"72258838",
X"810bff80",
X"135354ff",
X"bf125170",
X"99268638",
X"e01252b0",
X"39ff9f12",
X"51997127",
X"a738d012",
X"e0135451",
X"70892685",
X"38725298",
X"39728f26",
X"85387252",
X"8f3971ba",
X"2e098106",
X"85389a52",
X"83398052",
X"73802e85",
X"38818012",
X"527181ff",
X"0683c080",
X"0c853d0d",
X"04803d0d",
X"8498c051",
X"80717081",
X"05533470",
X"84a0c02e",
X"098106f0",
X"38823d0d",
X"04fe3d0d",
X"02970533",
X"51fef43f",
X"83c08008",
X"81ff0683",
X"c7dc0854",
X"52807324",
X"9b3883c8",
X"90081372",
X"83c89408",
X"07535371",
X"733483c7",
X"dc088105",
X"83c7dc0c",
X"843d0d04",
X"fa3d0d82",
X"800a1b55",
X"8057883d",
X"fc055479",
X"53745278",
X"51ffb8a4",
X"3f883d0d",
X"04fe3d0d",
X"83c7f408",
X"527451ff",
X"bfa83f83",
X"c080088c",
X"38765375",
X"5283c7f4",
X"0851c53f",
X"843d0d04",
X"fe3d0d83",
X"c7f40853",
X"75527451",
X"ffb9e63f",
X"83c08008",
X"8d387753",
X"765283c7",
X"f40851ff",
X"9f3f843d",
X"0d04f73d",
X"0d98ee3f",
X"83c08008",
X"81ff06ff",
X"05577683",
X"38815780",
X"ebcc3f83",
X"c0800883",
X"c0800856",
X"5a871533",
X"5473802e",
X"80df3874",
X"0881e3e4",
X"2e098106",
X"80d33880",
X"0b911633",
X"55597379",
X"2e80c638",
X"74569a16",
X"33547383",
X"2e098106",
X"a438a416",
X"70335558",
X"80527351",
X"96d83f80",
X"53805273",
X"5196f83f",
X"81145476",
X"74258338",
X"80547378",
X"34811980",
X"d8179117",
X"33565759",
X"78742e09",
X"8106ffbe",
X"3881c415",
X"8ca01b55",
X"5574742e",
X"098106ff",
X"88388b3d",
X"0d04f63d",
X"0d80eabe",
X"3f83c080",
X"087d83c0",
X"80085859",
X"5b7783c7",
X"dc0c8716",
X"33557480",
X"2e81a738",
X"75085473",
X"81e7942e",
X"09810693",
X"38901633",
X"53871633",
X"5281e884",
X"51e6f83f",
X"81883973",
X"81e3e42e",
X"09810680",
X"fd387452",
X"81e89851",
X"e6e13f80",
X"70911833",
X"565b5973",
X"792e80e6",
X"38a41657",
X"f6173355",
X"79802e91",
X"38ff1554",
X"73822689",
X"38a81870",
X"83c7dc0c",
X"5874812e",
X"09810687",
X"3881e8a0",
X"518d3974",
X"822e0981",
X"068a3881",
X"e8a851e6",
X"9a3f9539",
X"74832e09",
X"81068f38",
X"76338105",
X"5281e8b4",
X"51e6843f",
X"815a8119",
X"80d81891",
X"18335658",
X"5978742e",
X"098106ff",
X"9f38a818",
X"81c4178c",
X"a01d5657",
X"5875742e",
X"098106fe",
X"b8388c3d",
X"0d04fd3d",
X"0d83c7f4",
X"0851ffb5",
X"d93f83c0",
X"80089080",
X"2e098106",
X"ad388054",
X"83c18080",
X"5383c080",
X"085283c7",
X"f40851fb",
X"ef3f87c1",
X"80801433",
X"87c19080",
X"15348114",
X"54739080",
X"2e098106",
X"e938853d",
X"0d0481e8",
X"c40b83c0",
X"800c04fc",
X"3d0d7654",
X"73902e80",
X"ff387390",
X"248e3873",
X"842e9838",
X"73862ea6",
X"3882b939",
X"73932e81",
X"95387394",
X"2e81cf38",
X"82aa3981",
X"80805382",
X"80805283",
X"c7f00851",
X"fb8e3f82",
X"b5398054",
X"81808053",
X"80c08052",
X"83c7f008",
X"51faf93f",
X"82808053",
X"80c08052",
X"83c7f008",
X"51fae93f",
X"84818080",
X"14338481",
X"c0801534",
X"84828080",
X"14338482",
X"c0801534",
X"81145473",
X"80c0802e",
X"098106dc",
X"3881eb39",
X"82808053",
X"81808052",
X"83c7f008",
X"51fab13f",
X"80548482",
X"80801433",
X"84818080",
X"15348114",
X"54738180",
X"802e0981",
X"06e83881",
X"bd398180",
X"805380c0",
X"805283c7",
X"f00851fa",
X"833f8055",
X"84818080",
X"15547333",
X"8481c080",
X"16347333",
X"84828080",
X"16347333",
X"8482c080",
X"16348115",
X"557480c0",
X"802e0981",
X"06d63880",
X"fd398180",
X"8053a080",
X"5283c7f0",
X"0851f9c4",
X"3f805584",
X"81808015",
X"54733384",
X"81a08016",
X"34733384",
X"81c08016",
X"34733384",
X"81e08016",
X"34733384",
X"82808016",
X"34733384",
X"82a08016",
X"34733384",
X"82c08016",
X"34733384",
X"82e08016",
X"34811555",
X"74a0802e",
X"098106ff",
X"b6389f39",
X"f89b3f80",
X"0b83c7dc",
X"0c800b83",
X"c8940c81",
X"e8c851e2",
X"9a3f81b7",
X"8dc051f5",
X"fd3f863d",
X"0d04fc3d",
X"0d767052",
X"55ffb8fa",
X"3f83c080",
X"08548153",
X"83c08008",
X"80c23874",
X"51ffb8bc",
X"3f83c080",
X"0881e8e4",
X"5383c080",
X"085253d1",
X"9c3f83c0",
X"8008a138",
X"81e8e852",
X"7251d18d",
X"3f83c080",
X"08923881",
X"e8ec5272",
X"51d0fe3f",
X"83c08008",
X"802e8338",
X"81547353",
X"7283c080",
X"0c863d0d",
X"04f03d0d",
X"80dbae0b",
X"83c3ac0c",
X"83c7f008",
X"51d3a83f",
X"83c7f008",
X"51ffadf1",
X"3fff0b81",
X"e8e85383",
X"c0800852",
X"56d0be3f",
X"83c08008",
X"802e9f38",
X"8058923d",
X"d8115555",
X"9053f015",
X"5283c7f0",
X"0851ffaf",
X"e33f02bb",
X"05335681",
X"a53983c7",
X"f00851ff",
X"b0e03f83",
X"c0800857",
X"83c08008",
X"8280802e",
X"09810683",
X"38845683",
X"c0800881",
X"80802e09",
X"810680e1",
X"38805c80",
X"5b805a80",
X"59f6923f",
X"800b83c7",
X"dc0c800b",
X"83c8940c",
X"81e8f051",
X"e0913f80",
X"d00b83c7",
X"dc0c81e9",
X"8051e083",
X"3f80f80b",
X"83c7dc0c",
X"81e99451",
X"dff53f75",
X"8025a238",
X"8052893d",
X"7052558c",
X"893f8352",
X"74518c82",
X"3f785574",
X"80258338",
X"90568075",
X"25dd3886",
X"567680c0",
X"802e0981",
X"06853893",
X"568c3976",
X"a0802e09",
X"81068338",
X"94567551",
X"faad3f92",
X"3d0d04f6",
X"3d0d805a",
X"80598058",
X"80578070",
X"5656f589",
X"3f800b83",
X"c7dc0c80",
X"0b83c894",
X"0c81e9a8",
X"51df883f",
X"81800b83",
X"c8940c81",
X"e9ac51de",
X"fa3f80d0",
X"0b83c7dc",
X"0c743070",
X"76078025",
X"70872b83",
X"c8940c51",
X"53edcf3f",
X"83c08008",
X"5281e9b4",
X"51ded43f",
X"80f80b83",
X"c7dc0c74",
X"81327030",
X"70720780",
X"2570872b",
X"83c8940c",
X"515454f9",
X"a93f83c0",
X"80085281",
X"e9c051de",
X"aa3f81a0",
X"0b83c7dc",
X"0c748232",
X"70307072",
X"07802570",
X"872b83c8",
X"940c5154",
X"83c7f408",
X"5254ffaa",
X"e83f83c0",
X"80085281",
X"e9c851dd",
X"fa3f81c8",
X"0b83c7dc",
X"0c748332",
X"70307072",
X"07802570",
X"872b83c8",
X"940c5154",
X"83c7f008",
X"5254ffaa",
X"b83f81e9",
X"d05383c0",
X"8008802e",
X"8f3883c7",
X"f00851ff",
X"aaa33f83",
X"c0800853",
X"725281e9",
X"d851ddb3",
X"3f81f00b",
X"83c7dc0c",
X"74843270",
X"30707207",
X"80257087",
X"2b83c894",
X"0c515481",
X"e9e05254",
X"dd913f82",
X"c00b83c7",
X"dc0c7485",
X"32703070",
X"72078025",
X"70872b83",
X"c8940c51",
X"5481e9f8",
X"5254dcef",
X"3f800b83",
X"c8940c83",
X"9051f5ae",
X"3f868da0",
X"51f0c73f",
X"8052873d",
X"70525388",
X"f53f8352",
X"725188ee",
X"3f795372",
X"81cb3877",
X"15557480",
X"25853872",
X"55903985",
X"75258538",
X"85558739",
X"74852681",
X"aa387484",
X"2981e3cc",
X"05537208",
X"04eb8b3f",
X"83c08008",
X"77555373",
X"812e0981",
X"06893883",
X"c0800810",
X"53903973",
X"ff2e0981",
X"06883883",
X"c0800881",
X"2c539073",
X"25853890",
X"53883972",
X"80248338",
X"81537251",
X"eae53f80",
X"de39eaf7",
X"3f83c080",
X"08175372",
X"80258538",
X"80538839",
X"87732583",
X"38875372",
X"51eaf13f",
X"be397686",
X"3878802e",
X"b63883c3",
X"a40883c3",
X"a00caf99",
X"0b83c3ac",
X"0c83c7f4",
X"0851cdaf",
X"3ff5c73f",
X"9a397880",
X"2e9538f9",
X"e83f8153",
X"96397880",
X"2e8938f2",
X"b13f8439",
X"78873875",
X"802efbde",
X"38805372",
X"83c0800c",
X"8c3d0d04",
X"ff3d0d83",
X"c8805180",
X"edc33fed",
X"ba3f83c0",
X"8008802e",
X"86388051",
X"80da39ed",
X"bf3f83c0",
X"800880ce",
X"38edca3f",
X"83c08008",
X"802eaa38",
X"8151e8ea",
X"3fe5a43f",
X"800b83c7",
X"dc0cfb83",
X"3f83c080",
X"0852ff0b",
X"83c7dc0c",
X"e7b63f71",
X"a1387151",
X"e8c83f9f",
X"39edab3f",
X"83c08008",
X"802e9438",
X"8151e8b6",
X"3fe4f03f",
X"f8d73fe7",
X"933f8151",
X"eed23f83",
X"3d0d04fe",
X"3d0d8052",
X"83c88051",
X"80dd803f",
X"82808053",
X"80528181",
X"808051ed",
X"d63f80c0",
X"80538052",
X"84818080",
X"51ede73f",
X"90808052",
X"86848080",
X"51ffaaf7",
X"3f83c080",
X"08ad3883",
X"c7fc0851",
X"80f3a33f",
X"81ebb451",
X"ffafb13f",
X"83c7f408",
X"5381ea80",
X"5283c080",
X"0851ffaa",
X"903f83c0",
X"80088438",
X"f3b83f81",
X"51ede13f",
X"fe963ffc",
X"3983c08c",
X"080283c0",
X"8c0cfb3d",
X"0d0281ea",
X"8c0b83c3",
X"a40c81e8",
X"ec0b83c3",
X"9c0c81e8",
X"e80b83c3",
X"b40c81ea",
X"900b83c3",
X"b00c83c0",
X"8c08fc05",
X"0c800b83",
X"c7e00b83",
X"c08c08f8",
X"050c83c0",
X"8c08f405",
X"0cffa8e7",
X"3f83c080",
X"088605fc",
X"0683c08c",
X"08f0050c",
X"0283c08c",
X"08f00508",
X"310d833d",
X"7083c08c",
X"08f80508",
X"70840583",
X"c08c08f8",
X"050c0c51",
X"ffa4f83f",
X"83c08c08",
X"f4050881",
X"0583c08c",
X"08f4050c",
X"83c08c08",
X"f4050888",
X"2e098106",
X"ffab3886",
X"94808051",
X"e2b33fff",
X"0b83c7dc",
X"0c800b83",
X"c8940c84",
X"98c00b83",
X"c8900c81",
X"51e5f33f",
X"8151e698",
X"3f8051e6",
X"933f8151",
X"e6b93f82",
X"51e6e13f",
X"8051e7b6",
X"3f8051e7",
X"e03f80d3",
X"c5528051",
X"d7923ffd",
X"a63f83c0",
X"8c08fc05",
X"080d800b",
X"83c0800c",
X"873d0d83",
X"c08c0c04",
X"fa3d0d78",
X"5580750c",
X"800b8416",
X"0c800b88",
X"160c800b",
X"8c160c80",
X"0b90160c",
X"83c88051",
X"80e9be3f",
X"ea893f83",
X"c0800887",
X"d0883370",
X"81ff0651",
X"535671a7",
X"3887d080",
X"3383c8a8",
X"3487d081",
X"3383c8a0",
X"3487d082",
X"3383c898",
X"3487d083",
X"3383c89c",
X"34ff0b87",
X"d08b3487",
X"d0893387",
X"d08f3370",
X"822a7081",
X"06703070",
X"72077009",
X"709f2c77",
X"069e0657",
X"51515651",
X"51545480",
X"74980653",
X"5371882e",
X"09810683",
X"38815371",
X"98327030",
X"70802575",
X"71318419",
X"0c515152",
X"80748606",
X"53537182",
X"2e098106",
X"83388153",
X"71863270",
X"30708025",
X"75713178",
X"0c515152",
X"83c8a833",
X"5281aa72",
X"27843881",
X"750c83c8",
X"a8335271",
X"bb268438",
X"ff750c83",
X"c8a03352",
X"81aa7227",
X"8638810b",
X"84160c83",
X"c8a03352",
X"71bb2686",
X"38ff0b84",
X"160c83c8",
X"98335281",
X"aa722784",
X"3881750c",
X"83c89833",
X"5271bb26",
X"8438ff75",
X"0c83c89c",
X"335281aa",
X"72278638",
X"810b8416",
X"0c83c89c",
X"335271bb",
X"268638ff",
X"0b84160c",
X"80577394",
X"2eaa3887",
X"80903387",
X"80913387",
X"80923370",
X"81ff0672",
X"74060687",
X"80933371",
X"06810651",
X"52545454",
X"72772e09",
X"81068338",
X"81577688",
X"160c7580",
X"2eb03875",
X"812a7081",
X"06778106",
X"3184170c",
X"5275832a",
X"76822a71",
X"81067181",
X"0631770c",
X"53537584",
X"2a810688",
X"160c7585",
X"2a81068c",
X"160c883d",
X"0d04fe3d",
X"0d747654",
X"527151fc",
X"cf3f7281",
X"2ea23881",
X"73268d38",
X"72822ea8",
X"3872832e",
X"9c38e639",
X"7108e238",
X"841208dd",
X"38881208",
X"d838a539",
X"88120881",
X"2e9e3891",
X"39881208",
X"812e9538",
X"71089138",
X"8412088c",
X"388c1208",
X"812e0981",
X"06ffb238",
X"843d0d04",
X"fb3d0d78",
X"0284059f",
X"05335556",
X"800b81e5",
X"d0565381",
X"732b7406",
X"5271802e",
X"83388152",
X"74708205",
X"56227073",
X"902b0790",
X"809c0c51",
X"81135372",
X"882e0981",
X"06d93880",
X"5383c8b0",
X"13335170",
X"81ff2ebf",
X"38701081",
X"e3f00570",
X"22535171",
X"81ff2eaf",
X"38807074",
X"18703370",
X"1081e3f0",
X"05702251",
X"51515355",
X"5571712e",
X"96388114",
X"5473862e",
X"098106f1",
X"38719080",
X"9c0c7483",
X"c8a40c81",
X"13537286",
X"2e098106",
X"ffab3880",
X"53721670",
X"33515170",
X"81ff2e9f",
X"38701081",
X"e3f00570",
X"22515170",
X"81ff2e8f",
X"387083c8",
X"a40c7084",
X"80800790",
X"809c0c81",
X"13537286",
X"2e098106",
X"cc388053",
X"72165170",
X"3383c8b0",
X"14348113",
X"5372862e",
X"098106ec",
X"38873d0d",
X"0404fe3d",
X"0d750284",
X"05930533",
X"81065252",
X"70883871",
X"9080940c",
X"8e397081",
X"2e098106",
X"86387190",
X"80980c84",
X"3d0d04fb",
X"3d0d7898",
X"2b70982c",
X"7b982b70",
X"982c0290",
X"059f0533",
X"810683c8",
X"cc117033",
X"70982b70",
X"982c5158",
X"5c5a5651",
X"55515470",
X"742e0981",
X"06943883",
X"c8ac1233",
X"70982b70",
X"982c5152",
X"5670732e",
X"b1387375",
X"347283c8",
X"ac133483",
X"c8ad3383",
X"c8cd3371",
X"982b7190",
X"2b0783c8",
X"ac337088",
X"2b720783",
X"c8cc3371",
X"079080b8",
X"0c525953",
X"5452873d",
X"0d04fe3d",
X"0d748111",
X"33713371",
X"882b0783",
X"c0800c53",
X"51843d0d",
X"0483c8b8",
X"3383c080",
X"0c0483c0",
X"8c080283",
X"c08c0cf5",
X"3d0d83c0",
X"8c088805",
X"0883c08c",
X"088f0533",
X"83c08c08",
X"92052202",
X"8c057390",
X"0583c08c",
X"08e8050c",
X"83c08c08",
X"f8050c83",
X"c08c08f0",
X"050c83c0",
X"8c08ec05",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08f005",
X"0883c08c",
X"08e0050c",
X"83c08c08",
X"fc050c83",
X"c08c08f0",
X"05088927",
X"8a38890b",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"05088605",
X"87fffc06",
X"83c08c08",
X"e0050c02",
X"83c08c08",
X"e0050831",
X"0d853d70",
X"5583c08c",
X"08ec0508",
X"5483c08c",
X"08f00508",
X"5383c08c",
X"08f40508",
X"5283c08c",
X"08e4050c",
X"80e7b93f",
X"83c08008",
X"81ff0683",
X"c08c08e4",
X"050883c0",
X"8c08ec05",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"e0050880",
X"2e8c3883",
X"c08c08f8",
X"05080d89",
X"c83983c0",
X"8c08f005",
X"08802e89",
X"a63883c0",
X"8c08ec05",
X"08810533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508842e",
X"a938840b",
X"83c08c08",
X"e0050825",
X"88c73883",
X"c08c08e0",
X"0508852e",
X"859b3883",
X"c08c08e0",
X"0508a12e",
X"87ad3888",
X"ac39800b",
X"83c08c08",
X"ec050885",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08fc050c",
X"83c08c08",
X"e0050883",
X"2e098106",
X"88833883",
X"c08c08e8",
X"05088105",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e0050881",
X"2687e638",
X"810b83c0",
X"8c08e005",
X"0880d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08fc",
X"050c83c0",
X"8c08ec05",
X"08820533",
X"83c08c08",
X"e0050887",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088b",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"e005088c",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088d",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"e005088e",
X"052383c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088a",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"70940508",
X"fcffff06",
X"7194050c",
X"83c08c08",
X"e0050c83",
X"c08c08ec",
X"05088605",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"f4050c83",
X"c08c08e0",
X"050883c0",
X"8c08fc05",
X"082e0981",
X"06b63883",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c83",
X"c08c08fc",
X"050883c0",
X"8c08e005",
X"088b0534",
X"83c08c08",
X"ec050887",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"812e8f38",
X"83c08c08",
X"e0050882",
X"2eb73884",
X"8c3983c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c820b",
X"83c08c08",
X"e005088a",
X"053483d9",
X"3983c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08fc0508",
X"83c08c08",
X"e005088a",
X"053483a1",
X"3983c08c",
X"08fc0508",
X"802e8395",
X"3883c08c",
X"08ec0508",
X"83053383",
X"0683c08c",
X"08e0050c",
X"83c08c08",
X"e0050883",
X"2e098106",
X"82f33883",
X"c08c08ec",
X"05088205",
X"3370982b",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c83c0",
X"8c08e005",
X"08802582",
X"cc3883c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c83c0",
X"8c08ec05",
X"08860533",
X"83c08c08",
X"e0050880",
X"d6053483",
X"c08c08e0",
X"05088405",
X"83c08c08",
X"ec050882",
X"05338f06",
X"83c08c08",
X"e4050c83",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0883c08c",
X"08e00508",
X"3483c08c",
X"08ec0508",
X"84053383",
X"c08c08e0",
X"05088105",
X"34800b83",
X"c08c08e0",
X"05088205",
X"3483c08c",
X"08e00508",
X"08ff83ff",
X"06828007",
X"83c08c08",
X"e005080c",
X"83c08c08",
X"e8050881",
X"05338105",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"050883c0",
X"8c08e805",
X"08810534",
X"81833983",
X"c08c08fc",
X"0508802e",
X"80f73883",
X"c08c08ec",
X"05088605",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e00508a2",
X"2e098106",
X"80d73883",
X"c08c08ec",
X"05088805",
X"3383c08c",
X"08ec0508",
X"87053371",
X"82802905",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c5283c0",
X"8c08e405",
X"0c83c08c",
X"08f4050c",
X"83c08c08",
X"e4050883",
X"c08c08e0",
X"05088805",
X"2383c08c",
X"08ec0508",
X"3383c08c",
X"08f00508",
X"71317083",
X"ffff0683",
X"c08c08f0",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08ec0508",
X"0583c08c",
X"08ec050c",
X"f6d03983",
X"c08c08f8",
X"05080d83",
X"c08c08f0",
X"050883c0",
X"8c08e005",
X"0c83c08c",
X"08f80508",
X"0d83c08c",
X"08e00508",
X"83c0800c",
X"8d3d0d83",
X"c08c0c04",
X"83c08c08",
X"0283c08c",
X"0ce73d0d",
X"83c08c08",
X"88050802",
X"840583c0",
X"8c08e805",
X"0c83c08c",
X"08d4050c",
X"800b83c8",
X"d43483c0",
X"8c08d405",
X"08900583",
X"c08c08c4",
X"050c800b",
X"83c08c08",
X"c4050834",
X"800b83c0",
X"8c08c405",
X"08810534",
X"800b83c0",
X"8c08c805",
X"0c83c08c",
X"08c80508",
X"80d82983",
X"c08c08c4",
X"05080583",
X"c08c08ff",
X"b8050c80",
X"0b83c08c",
X"08ffb805",
X"0880d805",
X"0c83c08c",
X"08ffb805",
X"08840583",
X"c08c08ff",
X"b8050c83",
X"c08c08c8",
X"050883c0",
X"8c08ffb8",
X"05083488",
X"0b83c08c",
X"08ffb805",
X"08810534",
X"800b83c0",
X"8c08ffb8",
X"05088205",
X"3483c08c",
X"08ffb805",
X"0808ffa1",
X"ff06a080",
X"0783c08c",
X"08ffb805",
X"080c83c0",
X"8c08c805",
X"08810570",
X"81ff0683",
X"c08c08c8",
X"050c83c0",
X"8c08ffb8",
X"050c810b",
X"83c08c08",
X"c8050827",
X"fedb3883",
X"c08c08ec",
X"05705483",
X"c08c08cc",
X"050c9252",
X"83c08c08",
X"d4050851",
X"80dae03f",
X"83c08008",
X"81ff0670",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffbc0508",
X"91d93883",
X"c08c08f4",
X"0551f1ca",
X"3f83c080",
X"0883ffff",
X"0683c08c",
X"08f60552",
X"83c08c08",
X"e0050cf1",
X"b13f83c0",
X"800883ff",
X"ff0683c0",
X"8c08fd05",
X"3383c08c",
X"08ffbc05",
X"0883c08c",
X"08c8050c",
X"83c08c08",
X"c0050c83",
X"c08c08dc",
X"050c83c0",
X"8c08c805",
X"0883c08c",
X"08c00508",
X"2780fe38",
X"83c08c08",
X"cc050854",
X"83c08c08",
X"c8050853",
X"895283c0",
X"8c08d405",
X"085180d9",
X"e73f83c0",
X"800881ff",
X"0683c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffbc05",
X"0883eb38",
X"83c08c08",
X"ee0551f0",
X"b13f83c0",
X"800883ff",
X"ff065383",
X"c08c08c8",
X"05085283",
X"c08c08d4",
X"050851f0",
X"b53f83c0",
X"8c08c805",
X"08810570",
X"81ff0683",
X"c08c08c8",
X"050c83c0",
X"8c08ffb8",
X"050cfef2",
X"3983c08c",
X"08c40508",
X"81053383",
X"c08c08c0",
X"050c83c0",
X"8c08c005",
X"08839e38",
X"83c08c08",
X"c0050883",
X"c08c08ff",
X"b8050c83",
X"c08c08e0",
X"050888de",
X"2e098106",
X"8b38810b",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"dc050885",
X"8e2e0981",
X"0682c538",
X"817083c0",
X"8c08ffb8",
X"05080683",
X"c08c08ff",
X"b8050c83",
X"c08c08c8",
X"050c83c0",
X"8c08ffb8",
X"0508802e",
X"829e3883",
X"c08c08c8",
X"050883c0",
X"8c08c405",
X"08810534",
X"83c08c08",
X"c0050883",
X"c08c08c4",
X"05088705",
X"3483c08c",
X"08c00508",
X"83c08c08",
X"c405088b",
X"053483c0",
X"8c08c005",
X"0883c08c",
X"08c40508",
X"8c053483",
X"0b83c08c",
X"08c40508",
X"8d053483",
X"c08c08c0",
X"050883c0",
X"8c08c405",
X"088e0523",
X"830b83c0",
X"8c08c405",
X"088a0534",
X"83c08c08",
X"c4050894",
X"05088380",
X"800783c0",
X"8c08c405",
X"0894050c",
X"83c8b833",
X"7083c08c",
X"08c80508",
X"0583c08c",
X"08ffb805",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffb805",
X"0883c8b8",
X"3483c08c",
X"08ffbc05",
X"0883c08c",
X"08c40508",
X"94053483",
X"c08c08c8",
X"050883c0",
X"8c08c405",
X"0880d605",
X"3483c08c",
X"08c80508",
X"83c08c08",
X"c4050884",
X"05348e0b",
X"83c08c08",
X"c4050885",
X"053483c0",
X"8c08c005",
X"0883c08c",
X"08c40508",
X"86053483",
X"c08c08c4",
X"05088405",
X"08ff83ff",
X"06828007",
X"83c08c08",
X"c4050884",
X"050ca239",
X"81db0b83",
X"c08c08ff",
X"b8050c8c",
X"d63983c0",
X"8c08ffbc",
X"050883c0",
X"8c08ffb8",
X"050c8cc3",
X"3983c08c",
X"08f10533",
X"5283c08c",
X"08d40508",
X"5180d5ec",
X"3f800b83",
X"c08c08c4",
X"05088105",
X"3383c08c",
X"08ffb805",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"c8050883",
X"c08c08ff",
X"b8050827",
X"8aca3883",
X"c08c08c8",
X"050880d8",
X"297083c0",
X"8c08c405",
X"08057088",
X"05708305",
X"3383c08c",
X"08ffb805",
X"0c83c08c",
X"08cc050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"d8050c83",
X"c08c08ff",
X"b8050888",
X"893883c0",
X"8c08ffbc",
X"05088d05",
X"3383c08c",
X"08d0050c",
X"83c08c08",
X"d0050887",
X"ed3883c0",
X"8c08cc05",
X"08220284",
X"05718605",
X"87fffc06",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"e4050c83",
X"c08c08c0",
X"050c0283",
X"c08c08ff",
X"b8050831",
X"0d893d70",
X"5983c08c",
X"08c00508",
X"5883c08c",
X"08ffbc05",
X"08870533",
X"5783c08c",
X"08ffb805",
X"0ca25583",
X"c08c08d0",
X"05085486",
X"53818152",
X"83c08c08",
X"d4050851",
X"80c89f3f",
X"83c08008",
X"81ff0683",
X"c08c08d0",
X"050c83c0",
X"8c08d005",
X"0881c038",
X"83c08c08",
X"ffbc0508",
X"96055383",
X"c08c08c0",
X"05085283",
X"c08c08ff",
X"b8050851",
X"abd73f83",
X"c0800881",
X"ff0683c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"0508802e",
X"81853883",
X"c08c08ff",
X"bc050894",
X"0583c08c",
X"08ffbc05",
X"08960533",
X"70862a83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08c0",
X"050c83c0",
X"8c08ffb8",
X"0508832e",
X"09810680",
X"c63883c0",
X"8c08ffb8",
X"050883c0",
X"8c08cc05",
X"08820534",
X"83c8b833",
X"70810583",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"b8050883",
X"c8b83483",
X"c08c08ff",
X"bc050883",
X"c08c08c0",
X"05083483",
X"c08c08e4",
X"05080d83",
X"c08c08d0",
X"050881ff",
X"0683c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffbc05",
X"08fbe338",
X"83c08c08",
X"d8050883",
X"c08c08c4",
X"05080588",
X"05708205",
X"335183c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"0508832e",
X"09810680",
X"e33883c0",
X"8c08ffbc",
X"050883c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"05088105",
X"7081ff06",
X"5183c08c",
X"08ffb805",
X"0c810b83",
X"c08c08ff",
X"b8050827",
X"dd38800b",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"81057081",
X"ff065183",
X"c08c08ff",
X"b8050c97",
X"0b83c08c",
X"08ffb805",
X"0827dd38",
X"83c08c08",
X"e0050880",
X"f9327030",
X"70802551",
X"5183c08c",
X"08ffb805",
X"0c83c08c",
X"08dc0508",
X"912e0981",
X"0680f938",
X"83c08c08",
X"ffb80508",
X"802e80ec",
X"3883c08c",
X"08c80508",
X"80e23885",
X"0b83c08c",
X"08c40508",
X"a60534a0",
X"0b83c08c",
X"08c40508",
X"a7053485",
X"0b83c08c",
X"08c40508",
X"a8053480",
X"c00b83c0",
X"8c08c405",
X"08a90534",
X"860b83c0",
X"8c08c405",
X"08aa0534",
X"900b83c0",
X"8c08c405",
X"08ab0534",
X"860b83c0",
X"8c08c405",
X"08ac0534",
X"a00b83c0",
X"8c08c405",
X"08ad0534",
X"83c08c08",
X"e0050889",
X"d8327030",
X"70802551",
X"5183c08c",
X"08ffb805",
X"0c83c08c",
X"08dc0508",
X"83edec2e",
X"09810680",
X"f6388170",
X"83c08c08",
X"ffb80508",
X"0683c08c",
X"08ffb805",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffb805",
X"08802e80",
X"ce3883c0",
X"8c08c805",
X"0880c438",
X"840b83c0",
X"8c08c405",
X"08aa0534",
X"80c00b83",
X"c08c08c4",
X"0508ab05",
X"34840b83",
X"c08c08c4",
X"0508ac05",
X"34900b83",
X"c08c08c4",
X"0508ad05",
X"3483c08c",
X"08ffbc05",
X"0883c08c",
X"08c40508",
X"8c053483",
X"c08c08e0",
X"050880f9",
X"32703070",
X"80255151",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"dc050886",
X"2e098106",
X"80c33881",
X"7083c08c",
X"08ffb805",
X"080683c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb8",
X"0508802e",
X"9c3883c0",
X"8c08c805",
X"08933883",
X"c08c08ff",
X"bc050883",
X"c08c08c4",
X"05088d05",
X"3483c08c",
X"08e00508",
X"b4b43270",
X"30708025",
X"515183c0",
X"8c08ffb8",
X"050c83c0",
X"8c08dc05",
X"0890892e",
X"098106a2",
X"3883c08c",
X"08ffb805",
X"08802e96",
X"3883c08c",
X"08c80508",
X"8d38820b",
X"83c08c08",
X"c405088d",
X"053483c0",
X"8c08c805",
X"0880d829",
X"83c08c08",
X"c4050805",
X"70840570",
X"83053383",
X"c08c08ff",
X"b8050c83",
X"c08c08cc",
X"050c83c0",
X"8c08c005",
X"0c805880",
X"5783c08c",
X"08ffb805",
X"08568055",
X"80548a53",
X"a15283c0",
X"8c08d405",
X"085180c0",
X"d13f83c0",
X"800881ff",
X"06703070",
X"9f2a5183",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"bc0508a0",
X"2e8c3883",
X"c08c08ff",
X"b80508f5",
X"dd3883c0",
X"8c08c005",
X"088b0533",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"802eb338",
X"83c08c08",
X"cc050883",
X"053383c0",
X"8c08ffb8",
X"050c8058",
X"805783c0",
X"8c08ffb8",
X"05085680",
X"5580548b",
X"53a15283",
X"c08c08d4",
X"050851bf",
X"cd3f83c0",
X"8c08c805",
X"08810570",
X"81ff0683",
X"c08c08c4",
X"05088105",
X"335283c0",
X"8c08c805",
X"0c83c08c",
X"08ffb805",
X"0cf5a539",
X"800b83c0",
X"8c08c805",
X"0c83c08c",
X"08c80508",
X"80d82983",
X"c08c08d4",
X"05080570",
X"9a053383",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050882",
X"2e098106",
X"bd3883c0",
X"8c08ffb8",
X"05089705",
X"3383c8d4",
X"5983c08c",
X"08ffb805",
X"0c815783",
X"c08c08ff",
X"b8050856",
X"83c08c08",
X"ffbc0508",
X"55805489",
X"53a15283",
X"c08c08d4",
X"050851be",
X"a93f83c0",
X"8c08c805",
X"08810570",
X"81ff0683",
X"c08c08c8",
X"050c83c0",
X"8c08ffb8",
X"050c810b",
X"83c08c08",
X"c8050827",
X"fee73881",
X"0b83c08c",
X"08c40508",
X"34800b83",
X"c08c08ff",
X"b8050c83",
X"c08c08e8",
X"05080d83",
X"c08c08ff",
X"b8050883",
X"c0800c9b",
X"3d0d83c0",
X"8c0c04f4",
X"3d0d901f",
X"59800b81",
X"1a33555b",
X"7a742781",
X"ad387a80",
X"d829198a",
X"11335555",
X"73832e09",
X"81068188",
X"38941533",
X"57805276",
X"51de8b3f",
X"80538052",
X"7651deab",
X"3fb2ab3f",
X"83c08008",
X"5c805877",
X"81c4291c",
X"87113355",
X"5573802e",
X"80c03874",
X"0881e3e4",
X"2e098106",
X"b5388075",
X"5b567580",
X"d8291a9a",
X"11335555",
X"73832e09",
X"81069238",
X"a4157033",
X"55557674",
X"278738ff",
X"14547375",
X"34811670",
X"81ff0657",
X"54817627",
X"d1388118",
X"7081ff06",
X"59548778",
X"27ffa438",
X"83c8b833",
X"ff055473",
X"83c8b834",
X"811b7081",
X"ff06811b",
X"335f5c54",
X"7c7b26fe",
X"d538800b",
X"83c0800c",
X"8e3d0d04",
X"83c08c08",
X"0283c08c",
X"0ce63d0d",
X"83c08c08",
X"88050802",
X"84057190",
X"05703370",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"cc050c83",
X"c08c08dc",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08ffa405",
X"08802e9f",
X"8c38800b",
X"83c08c08",
X"cc050881",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08d405",
X"0c83c08c",
X"08d40508",
X"83c08c08",
X"ffa40508",
X"259ed438",
X"83c08c08",
X"d4050880",
X"d82983c0",
X"8c08cc05",
X"08058405",
X"70860533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffa40508",
X"802e9de0",
X"38afd73f",
X"83c08c08",
X"ffbc0508",
X"80d40508",
X"83c08008",
X"269dc938",
X"0283c08c",
X"08ffbc05",
X"08810533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"d8050c83",
X"c08c08ff",
X"a4050883",
X"c08c08fc",
X"052383c0",
X"8c08ffa4",
X"05088605",
X"83fc0683",
X"c08c08ff",
X"a4050c02",
X"83c08c08",
X"ffa40508",
X"310d853d",
X"705583c0",
X"8c08fc05",
X"5483c08c",
X"08ffbc05",
X"085383c0",
X"8c08e005",
X"085283c0",
X"8c08c005",
X"0cb7ab3f",
X"83c08008",
X"81ff0683",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a405089c",
X"923883c0",
X"8c08ffbc",
X"05088705",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e80",
X"d53883c0",
X"8c08ffbc",
X"05088605",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08822e09",
X"8106b338",
X"83c08c08",
X"fc052283",
X"c08c08ff",
X"a4050c87",
X"0b83c08c",
X"08ffa405",
X"08279738",
X"83c08c08",
X"c0050882",
X"055283c0",
X"8c08c005",
X"083351d7",
X"c73f83c0",
X"8c08ffbc",
X"05088605",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08832e09",
X"81069afb",
X"3883c08c",
X"08ffbc05",
X"08920583",
X"c08c08ff",
X"bc050889",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08c405",
X"0c83c08c",
X"08ffa405",
X"08832eb6",
X"3883c08c",
X"08c40508",
X"82053383",
X"c08c08fc",
X"052283c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa8",
X"050883c0",
X"8c08ffac",
X"0508269a",
X"9638800b",
X"83c08c08",
X"e4050c80",
X"0b83c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa405",
X"08832e09",
X"810688c1",
X"3883c08c",
X"08c00508",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffb005",
X"082e0981",
X"0687fa38",
X"83c08c08",
X"c0050881",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508942e",
X"09810687",
X"d83883c0",
X"8c08c005",
X"08820533",
X"70810683",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"b005082e",
X"8a38880b",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"a8050881",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e91",
X"3883c08c",
X"08e40508",
X"840783c0",
X"8c08e405",
X"0c83c08c",
X"08ffa805",
X"08822a70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e913883",
X"c08c08e4",
X"05088207",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"a8050883",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e91",
X"3883c08c",
X"08e40508",
X"810783c0",
X"8c08e405",
X"0c83c08c",
X"08c00508",
X"83053370",
X"982b83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"05088025",
X"913883c0",
X"8c08e405",
X"08900783",
X"c08c08e4",
X"050c83c0",
X"8c08ffa8",
X"050881ff",
X"0670852a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa40508",
X"802e9138",
X"83c08c08",
X"e40508a0",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"ffa80508",
X"842a7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"923883c0",
X"8c08e405",
X"0880c007",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"a8050886",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e92",
X"3883c08c",
X"08e40508",
X"81800783",
X"c08c08e4",
X"050c83c0",
X"8c08ffa8",
X"05088106",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9238",
X"83c08c08",
X"e4050882",
X"800783c0",
X"8c08e405",
X"0c83c08c",
X"08ffa805",
X"08812a70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e923883",
X"c08c08e4",
X"05088480",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"c0050884",
X"05337098",
X"2b83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa405",
X"08802592",
X"3883c08c",
X"08e40508",
X"88800783",
X"c08c08e4",
X"050c83c0",
X"8c08c005",
X"08850533",
X"70982b83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050880",
X"25923883",
X"c08c08e4",
X"05089080",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"c0050882",
X"05337081",
X"ff067085",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa405",
X"08802e92",
X"3883c08c",
X"08e40508",
X"a0800783",
X"c08c08e4",
X"050c83c0",
X"8c08ffa8",
X"0508842a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9338",
X"83c08c08",
X"e4050880",
X"c0800783",
X"c08c08e4",
X"050c83c0",
X"8c08ffa8",
X"0508862a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9338",
X"83c08c08",
X"e4050881",
X"80800783",
X"c08c08e4",
X"050c83c0",
X"8c08ffac",
X"0508982b",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"80259338",
X"83c08c08",
X"e4050882",
X"80800783",
X"c08c08e4",
X"050c83c0",
X"8c08c005",
X"08870533",
X"70982b83",
X"c08c08c0",
X"05088905",
X"3370982b",
X"70982c73",
X"982c8180",
X"05545153",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa80508",
X"83c08c08",
X"f8052380",
X"ff0b83c0",
X"8c08ffa4",
X"05083183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08fa",
X"052384d9",
X"39800b83",
X"c08c08e4",
X"050c8180",
X"0b83c08c",
X"08f80523",
X"81800b83",
X"c08c08fa",
X"052384b9",
X"3983c08c",
X"08ffb005",
X"081083c0",
X"8c0805f8",
X"0583c08c",
X"08ffb005",
X"08842983",
X"c08c08ff",
X"b0050810",
X"0583c08c",
X"08c40508",
X"05708405",
X"703383c0",
X"8c08c005",
X"08057033",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffb80508",
X"2383c08c",
X"08ffa805",
X"08810533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"902e0981",
X"06be3883",
X"c08c08ff",
X"a8050833",
X"83c08c08",
X"c0050805",
X"81057033",
X"70828029",
X"83c08c08",
X"ffb40508",
X"05515183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"b8050823",
X"83c08c08",
X"ffac0508",
X"86052283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a80508a2",
X"3883c08c",
X"08ffac05",
X"08880522",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"81ff2e80",
X"e53883c0",
X"8c08ffb8",
X"05082270",
X"83c08c08",
X"ffa80508",
X"31708280",
X"29713183",
X"c08c08ff",
X"ac050888",
X"05227083",
X"c08c08ff",
X"a8050831",
X"70733553",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffb805",
X"082383c0",
X"8c08ffb0",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa4050c",
X"810b83c0",
X"8c08ffb0",
X"050827fc",
X"e038800b",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffb00508",
X"1083c08c",
X"08c40508",
X"05709005",
X"703383c0",
X"8c08c005",
X"08057033",
X"72810533",
X"70720651",
X"535183c0",
X"8c08ffa8",
X"050c5183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e9b3890",
X"0b83c08c",
X"08ffb005",
X"082b83c0",
X"8c08e405",
X"080783c0",
X"8c08e405",
X"0c83c08c",
X"08ffb005",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a4050c97",
X"0b83c08c",
X"08ffb005",
X"0827fef4",
X"3883c08c",
X"08f80522",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"bf269138",
X"83c08c08",
X"e4050882",
X"0783c08c",
X"08e4050c",
X"81c00b83",
X"c08c08ff",
X"a4050827",
X"913883c0",
X"8c08e405",
X"08810783",
X"c08c08e4",
X"050c83c0",
X"8c08fa05",
X"2283c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08bf2691",
X"3883c08c",
X"08e40508",
X"880783c0",
X"8c08e405",
X"0c81c00b",
X"83c08c08",
X"ffa40508",
X"27913883",
X"c08c08e4",
X"05088407",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"bc050890",
X"053383c0",
X"8c08e405",
X"0883c08c",
X"08ffa405",
X"0c83c08c",
X"08c4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffbc0508",
X"8c05082e",
X"85e03883",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"bc05088c",
X"050c83c0",
X"8c08ffbc",
X"05088905",
X"3383c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa805",
X"08802e85",
X"9a3883c0",
X"8c08e405",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffa40508",
X"8f0683c0",
X"8c08e405",
X"0c83c08c",
X"08ffb005",
X"0c83c08c",
X"08d0050c",
X"83c08c08",
X"ffa80508",
X"822e0981",
X"0681c238",
X"800b83c0",
X"8c08ffa4",
X"0508862a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffa80508",
X"2e8c3881",
X"c00b83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffb0",
X"0508872a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9438",
X"83c08c08",
X"ffa80508",
X"81903283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"b0050884",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e94",
X"3883c08c",
X"08ffa805",
X"0880d032",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffb00508",
X"83c08c08",
X"ffa80508",
X"3283c08c",
X"08ffb005",
X"0c800b83",
X"c08c08f0",
X"050c800b",
X"83c08c08",
X"f4052380",
X"0b81e5e0",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffb805",
X"082e82d3",
X"3883c08c",
X"08f00581",
X"e5e00b83",
X"c08c08ff",
X"ac050c83",
X"c08c08c8",
X"050c83c0",
X"8c08ffac",
X"05083383",
X"c08c08ff",
X"ac050881",
X"05338172",
X"2b81722b",
X"077083c0",
X"8c08ffb0",
X"05080652",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffa80508",
X"2e098106",
X"81be3883",
X"c08c08ff",
X"b8050885",
X"2680f638",
X"83c08c08",
X"ffac0508",
X"82053370",
X"81ff0683",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050880",
X"2e80ca38",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"ffb80508",
X"81057081",
X"ff0683c0",
X"8c08c805",
X"08730553",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffa40508",
X"3483c08c",
X"08ffac05",
X"08830533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9d38",
X"810b83c0",
X"8c08ffa4",
X"05082b83",
X"c08c08d0",
X"05080807",
X"83c08c08",
X"d005080c",
X"83c08c08",
X"ffac0508",
X"84057033",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa40508",
X"fdc83883",
X"c08c08f0",
X"05528051",
X"c28e3f83",
X"c08c08e4",
X"05085283",
X"c08c08c4",
X"050851c3",
X"e13f83c0",
X"8c08fb05",
X"33708180",
X"0a29810a",
X"0570982c",
X"5583c08c",
X"08ffa405",
X"0c83c08c",
X"08f90533",
X"7081800a",
X"29810a05",
X"70982c55",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"c4050853",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa8050c",
X"c3b93f83",
X"c08c08ff",
X"bc050888",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"84e13883",
X"c08c08ff",
X"bc050890",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"05088126",
X"84c13880",
X"7081e698",
X"0b81e698",
X"0b810533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffb40508",
X"2e81ae38",
X"83c08c08",
X"ffac0508",
X"842983c0",
X"8c08ffa8",
X"05080570",
X"3383c08c",
X"08c00508",
X"05703372",
X"81053370",
X"72065153",
X"5183c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802eaa",
X"38810b83",
X"c08c08ff",
X"ac05082b",
X"83c08c08",
X"ffb40508",
X"077083ff",
X"ff0683c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffac",
X"05088105",
X"7081ff06",
X"81e69871",
X"84297105",
X"70810533",
X"515383c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508fed4",
X"3883c08c",
X"08ffbc05",
X"088a0522",
X"83c08c08",
X"c0050c83",
X"c08c08ff",
X"b4050883",
X"c08c08c0",
X"05082e82",
X"ae38800b",
X"83c08c08",
X"e8050c80",
X"0b83c08c",
X"08ec0523",
X"807083c0",
X"8c08e805",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffb0050c",
X"81af3983",
X"c08c08ff",
X"b4050883",
X"c08c08ff",
X"ac05082c",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e80e7",
X"3883c08c",
X"08ffb005",
X"0883c08c",
X"08ffb005",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"b8050873",
X"0583c08c",
X"08ffbc05",
X"08900533",
X"83c08c08",
X"ffac0508",
X"84290553",
X"5383c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa805",
X"0881e69a",
X"053383c0",
X"8c08ffa4",
X"05083483",
X"c08c08ff",
X"ac050881",
X"057081ff",
X"0683c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa405",
X"0c8f0b83",
X"c08c08ff",
X"ac050827",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb00508",
X"85268c38",
X"83c08c08",
X"ffa40508",
X"fea93883",
X"c08c08e8",
X"05528051",
X"ffbcbd3f",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffbc0508",
X"8a052383",
X"c08c08ff",
X"bc050880",
X"d2053383",
X"c08c08ff",
X"bc050880",
X"d4050805",
X"83c08c08",
X"ffbc0508",
X"80d4050c",
X"83c08c08",
X"d805080d",
X"83c08c08",
X"d4050881",
X"800a2981",
X"800a0570",
X"982c83c0",
X"8c08cc05",
X"08810533",
X"83c08c08",
X"ffa8050c",
X"5183c08c",
X"08d4050c",
X"83c08c08",
X"ffa80508",
X"83c08c08",
X"d4050824",
X"e1ae3880",
X"0b83c08c",
X"08ffa805",
X"0c83c08c",
X"08dc0508",
X"0d83c08c",
X"08ffa805",
X"0883c080",
X"0c9c3d0d",
X"83c08c0c",
X"04e93d0d",
X"696c0288",
X"0580ea05",
X"225c5a5b",
X"80707141",
X"5e58ff78",
X"797a7b7c",
X"7d464c4a",
X"45405d43",
X"62993d34",
X"62028405",
X"80dd0534",
X"77792280",
X"ffff0654",
X"45727923",
X"79782e88",
X"87387a70",
X"81055c33",
X"70842a71",
X"8c067082",
X"2a5a5656",
X"8306ff1b",
X"7083ffff",
X"065c5456",
X"80547574",
X"2e91387a",
X"7081055c",
X"33ff1b70",
X"83ffff06",
X"5c545481",
X"76279b38",
X"7381ff06",
X"7b708105",
X"5d335574",
X"82802905",
X"ff1b7083",
X"ffff065c",
X"54548276",
X"27aa3873",
X"83ffff06",
X"7b708105",
X"5d337090",
X"2b72077d",
X"7081055f",
X"3370982b",
X"7207fe1f",
X"7083ffff",
X"06405252",
X"52525454",
X"7e802e80",
X"c4387686",
X"f738748a",
X"2e098106",
X"9438811f",
X"7081ff06",
X"811e7081",
X"ff065f52",
X"405386dc",
X"39748c2e",
X"09810686",
X"d338ff1f",
X"7081ff06",
X"ff1e7081",
X"ff065f52",
X"40537b63",
X"2586bd38",
X"ff4386b8",
X"3976812e",
X"83bb3876",
X"81248938",
X"76802e8d",
X"3886a539",
X"76822e84",
X"a638869c",
X"39f81553",
X"72842684",
X"95387284",
X"2981e6d8",
X"05537208",
X"0464802e",
X"80cd3878",
X"22838080",
X"06537283",
X"80802e09",
X"8106bc38",
X"80567564",
X"27a43875",
X"1e7083ff",
X"ff067710",
X"1b901172",
X"832a5851",
X"57515373",
X"75347287",
X"0681712b",
X"51537281",
X"16348116",
X"7081ff06",
X"57539776",
X"27cc387f",
X"84074080",
X"0b993d43",
X"56611670",
X"3370982b",
X"70982c51",
X"51515380",
X"732480fb",
X"38607329",
X"1e7083ff",
X"ff067a22",
X"83808006",
X"52585372",
X"8380802e",
X"09810680",
X"de386088",
X"32703070",
X"72078025",
X"63903270",
X"30707207",
X"80257307",
X"53545851",
X"55537380",
X"2ebd3876",
X"87065372",
X"b6387584",
X"29761005",
X"79118411",
X"79832a57",
X"57515373",
X"75346081",
X"16346586",
X"14236688",
X"14237587",
X"387f8107",
X"408d3975",
X"812e0981",
X"0685387f",
X"82074081",
X"167081ff",
X"06575381",
X"7627fee5",
X"38636129",
X"1e7083ff",
X"ff065f53",
X"80704642",
X"ff028405",
X"80dd0534",
X"ff0b993d",
X"3483f539",
X"811c7081",
X"ff065d53",
X"80427381",
X"2e098106",
X"8e387781",
X"800a2981",
X"800a0558",
X"80d33973",
X"802e8938",
X"73822e09",
X"81068d38",
X"7c81800a",
X"2981800a",
X"055da439",
X"815f83b8",
X"39ff1c70",
X"81ff065d",
X"537b6325",
X"8338ff43",
X"7c802e92",
X"387c8180",
X"0a2981ff",
X"0a055d7c",
X"982c5d83",
X"93397780",
X"2e923877",
X"81800a29",
X"81ff0a05",
X"5877982c",
X"5882fd39",
X"7753839e",
X"39748926",
X"80f43874",
X"842981e6",
X"ec055372",
X"08047387",
X"2e82e138",
X"73852e82",
X"db387388",
X"2e82d538",
X"738c2e82",
X"cf387389",
X"2e098106",
X"86388145",
X"82c23973",
X"812e0981",
X"0682b938",
X"62802582",
X"b3387b98",
X"2b70982c",
X"514382a8",
X"397383ff",
X"ff064682",
X"9f397383",
X"ffff0647",
X"82963973",
X"81ff0641",
X"828e3973",
X"811a3482",
X"87397381",
X"ff064481",
X"ff397e53",
X"82a03974",
X"812e81e3",
X"38748124",
X"89387480",
X"2e8d3881",
X"e7397482",
X"2e81d838",
X"81de3974",
X"567b8338",
X"81567453",
X"73862e09",
X"81069738",
X"75810653",
X"72802e8e",
X"38782282",
X"ffff06fe",
X"80800753",
X"b6397b83",
X"38815373",
X"822e0981",
X"06973872",
X"81065372",
X"802e8e38",
X"782281ff",
X"ff068180",
X"80075393",
X"397b9638",
X"fc145372",
X"81268e38",
X"7822ff80",
X"80075372",
X"792380e5",
X"39805573",
X"812e0981",
X"06833873",
X"55775377",
X"802e8938",
X"74810653",
X"7280ca38",
X"72d01554",
X"55728126",
X"83388155",
X"77802eb9",
X"38748106",
X"5372802e",
X"b0387822",
X"83808006",
X"53728380",
X"802e0981",
X"069f3873",
X"b02e0981",
X"06873861",
X"993d3491",
X"3973b12e",
X"09810689",
X"38610284",
X"0580dd05",
X"34618105",
X"538c3961",
X"74318105",
X"53843961",
X"14537283",
X"ffff0642",
X"79f7fb38",
X"7d832a53",
X"72821a34",
X"78228380",
X"80065372",
X"8380802e",
X"09810688",
X"3881537f",
X"872e8338",
X"80537283",
X"c0800c99",
X"3d0d04fd",
X"3d0d7583",
X"11338212",
X"3371982b",
X"71902b07",
X"81143370",
X"882b7207",
X"75337107",
X"83c0800c",
X"52535456",
X"5452853d",
X"0d04f63d",
X"0d02b705",
X"33028405",
X"bb053302",
X"8805bf05",
X"335b5b5b",
X"80588057",
X"78882b7a",
X"07568055",
X"7a548153",
X"a3527c51",
X"92c83f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f63d",
X"0d02b705",
X"33028405",
X"bb053302",
X"8805bf05",
X"335b5b5b",
X"80588057",
X"78882b7a",
X"07568055",
X"7a548353",
X"a3527c51",
X"928c3f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f73d",
X"0d02b305",
X"33028405",
X"b6052260",
X"5a585680",
X"55805480",
X"5381a352",
X"7b5191de",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8b3d0d04",
X"ee3d0d64",
X"90115c5c",
X"807b3480",
X"0b841c0c",
X"800b881c",
X"34810b89",
X"1c34880b",
X"8a1c3480",
X"0b8b1c34",
X"881b08c1",
X"06810788",
X"1c0c8f3d",
X"70545d88",
X"527b519c",
X"8e3f83c0",
X"800881ff",
X"06705b59",
X"7881a938",
X"903d335e",
X"81db5a7d",
X"892e0981",
X"06819938",
X"7c539252",
X"7b519be7",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"8182387c",
X"58885778",
X"56a95578",
X"54865381",
X"a0527b51",
X"90cc3f83",
X"c0800881",
X"ff06705b",
X"597880e0",
X"3802ba05",
X"337b347c",
X"5478537d",
X"527b519b",
X"cf3f83c0",
X"800881ff",
X"06705b59",
X"7880c138",
X"02bd0533",
X"527b519b",
X"e73f83c0",
X"800881ff",
X"06705b59",
X"78aa3881",
X"7b335a5a",
X"79792699",
X"38805479",
X"5388527b",
X"51fdbb3f",
X"811a7081",
X"ff067c33",
X"525b59e4",
X"39810b88",
X"1c34805a",
X"7983c080",
X"0c943d0d",
X"04800b83",
X"c0800c04",
X"f93d0d79",
X"028405ab",
X"05338e3d",
X"70545858",
X"58ffb1ca",
X"3f8a3d8a",
X"0551ffb1",
X"c13f7551",
X"fc8d3f83",
X"c0800884",
X"86812ebe",
X"3883c080",
X"08848681",
X"26993883",
X"c0800884",
X"82802e80",
X"e63883c0",
X"80088482",
X"812e9f38",
X"81b43983",
X"c0800880",
X"c082832e",
X"80f43883",
X"c0800880",
X"c086832e",
X"80e83881",
X"993983c0",
X"a4335580",
X"5674762e",
X"09810681",
X"8b387454",
X"76539152",
X"7751fbd6",
X"3f745476",
X"53905277",
X"51fbcb3f",
X"74547653",
X"84527751",
X"fbfc3f81",
X"0b83c0a4",
X"3481b156",
X"80de3980",
X"54765391",
X"527751fb",
X"a93f8054",
X"76539052",
X"7751fb9e",
X"3f800b83",
X"c0a43476",
X"52871833",
X"5197923f",
X"b5398054",
X"76539452",
X"7751fb82",
X"3f805476",
X"53905277",
X"51faf73f",
X"7551ffaf",
X"f53f83c0",
X"8008892a",
X"81065376",
X"52871833",
X"5190c93f",
X"800b83c0",
X"a4348056",
X"7583c080",
X"0c893d0d",
X"04f23d0d",
X"6090115a",
X"58800b88",
X"1a337159",
X"56567476",
X"2e82a538",
X"82ac3f84",
X"190883c0",
X"80082682",
X"95387833",
X"5a810b8e",
X"3d23903d",
X"f81155f4",
X"05539918",
X"5277518a",
X"e13f83c0",
X"800881ff",
X"06705755",
X"74772e09",
X"810681d9",
X"38863974",
X"5681d239",
X"81568257",
X"8e3d3377",
X"06557480",
X"2ebb3880",
X"0b8d3d34",
X"903df005",
X"54845375",
X"527751fa",
X"cd3f83c0",
X"800881ff",
X"0655749d",
X"387b5375",
X"527751fc",
X"e73f83c0",
X"800881ff",
X"06557481",
X"b12e818b",
X"3874ffb3",
X"38761081",
X"fc068117",
X"7081ff06",
X"58565787",
X"7627ffa8",
X"38815675",
X"7a2680eb",
X"38800b8d",
X"3d348c3d",
X"70555784",
X"53755277",
X"51f9f73f",
X"83c08008",
X"81ff0655",
X"7480c138",
X"7651ffad",
X"f13f83c0",
X"80088287",
X"06557482",
X"812e0981",
X"06aa3802",
X"ae053381",
X"07557402",
X"8405ae05",
X"347b5375",
X"527751fb",
X"eb3f83c0",
X"800881ff",
X"06557481",
X"b12e9038",
X"74feb838",
X"81167081",
X"ff065755",
X"ff913980",
X"567581ff",
X"0656973f",
X"83c08008",
X"8fd00584",
X"1a0c7557",
X"7683c080",
X"0c903d0d",
X"0404803d",
X"0d9080a0",
X"08708a2c",
X"83c0800c",
X"51823d0d",
X"040483c8",
X"d80b83c0",
X"800c04fd",
X"3d0d7577",
X"5454800b",
X"83c8b834",
X"728a3890",
X"90800b84",
X"150c9039",
X"72812e09",
X"81068838",
X"9098800b",
X"84150c84",
X"140883c8",
X"d00c800b",
X"88150c80",
X"0b8c150c",
X"83c8d008",
X"53820b87",
X"80143487",
X"e851ff90",
X"893f83c8",
X"d0085380",
X"0b881434",
X"83c8d008",
X"53810b87",
X"80143483",
X"c8d00853",
X"800b8c14",
X"3483c8d0",
X"0853800b",
X"a4143491",
X"7434800b",
X"83c0a834",
X"800b83c0",
X"ac34800b",
X"83c0b034",
X"80547381",
X"c42983c8",
X"dc055380",
X"0b831434",
X"81147081",
X"ff065553",
X"877427e6",
X"38853d0d",
X"04fe3d0d",
X"74768211",
X"3370bf06",
X"81712bff",
X"05565151",
X"52539071",
X"278338ff",
X"52765171",
X"712383c8",
X"d0085187",
X"13339012",
X"34800b83",
X"c0ac3480",
X"0b83c0b0",
X"34881333",
X"8a143352",
X"5271802e",
X"aa387081",
X"ff065184",
X"52708338",
X"70527183",
X"c0ac348a",
X"13337030",
X"70802584",
X"2b708807",
X"51515253",
X"7083c0b0",
X"34903970",
X"81ff0651",
X"70833898",
X"527183c0",
X"b034800b",
X"83c0800c",
X"843d0d04",
X"f13d0d61",
X"6568028c",
X"0580cb05",
X"33029005",
X"80ce0522",
X"02940580",
X"d6052242",
X"40415a40",
X"40fd8f3f",
X"83c08008",
X"a788055b",
X"8070715b",
X"5b528394",
X"3983c8d0",
X"08517d94",
X"123483c0",
X"ac338107",
X"55807054",
X"567f8626",
X"80ea387f",
X"842981e7",
X"a00583c8",
X"d0085351",
X"70080480",
X"0b841334",
X"a1397733",
X"70307080",
X"25837131",
X"51515253",
X"70841334",
X"8d39810b",
X"841334b8",
X"39830b84",
X"13348170",
X"5456ad39",
X"810b8413",
X"34a23977",
X"33703070",
X"80258371",
X"31515152",
X"53708413",
X"34807833",
X"52527083",
X"38815271",
X"78348153",
X"74880755",
X"83c0b033",
X"83c8d008",
X"5257810b",
X"81d01234",
X"83c8d008",
X"51810b81",
X"9012347e",
X"802eae38",
X"72802ea9",
X"387eff1e",
X"52547083",
X"ffff0653",
X"7283ffff",
X"2e973873",
X"70810555",
X"3383c8d0",
X"08535170",
X"81c01334",
X"ff1351de",
X"3983c8d0",
X"08a81133",
X"53517688",
X"123483c8",
X"d0085174",
X"713481ff",
X"52913983",
X"c8d008a0",
X"11337081",
X"06515253",
X"708f38fb",
X"813f7a83",
X"c0800826",
X"e6388188",
X"39810ba0",
X"143483c8",
X"d008a811",
X"3380ff06",
X"70780752",
X"53517080",
X"2e80ed38",
X"71862a70",
X"81065151",
X"70802e91",
X"38807833",
X"52537083",
X"38815372",
X"783480e0",
X"3971842a",
X"70810651",
X"5170802e",
X"9b388119",
X"7083ffff",
X"067d3070",
X"9f2a5152",
X"5a51787c",
X"2e098106",
X"af38a439",
X"71832a70",
X"81065151",
X"70802e93",
X"38811a70",
X"81ff065b",
X"5179832e",
X"09810690",
X"388a3971",
X"a3065170",
X"802e8538",
X"71519239",
X"f9e83f7a",
X"83c08008",
X"26fce238",
X"7181bf06",
X"517083c0",
X"800c913d",
X"0d04f63d",
X"0d02b305",
X"33028405",
X"b7053302",
X"8805ba05",
X"22595959",
X"800b8c3d",
X"348c3dfc",
X"05568055",
X"80547653",
X"77527851",
X"fbf23f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f33d",
X"0d7f6264",
X"028c0580",
X"c2052272",
X"22811533",
X"425f415e",
X"59598078",
X"237d5378",
X"33528151",
X"ffa03f83",
X"c0800881",
X"ff065675",
X"802e8638",
X"755481ad",
X"3983c8d0",
X"08a81133",
X"821b3370",
X"862a7081",
X"0673982b",
X"5351575c",
X"56577980",
X"25833881",
X"5673762e",
X"873881f0",
X"54818239",
X"818c1733",
X"7081ff06",
X"79227d71",
X"31902b70",
X"902c7009",
X"709f2c72",
X"06705252",
X"53515357",
X"57547574",
X"24833875",
X"55748480",
X"8029fc80",
X"80057090",
X"2c515574",
X"ff2e9438",
X"83c8d008",
X"81801133",
X"5154737c",
X"7081055e",
X"34db3977",
X"22760554",
X"73782379",
X"09709f2a",
X"70810682",
X"1c3381bf",
X"0671862b",
X"07515151",
X"5473821a",
X"347c7626",
X"8a387722",
X"547a7426",
X"febb3880",
X"547383c0",
X"800c8f3d",
X"0d04f93d",
X"0d7a5780",
X"0b893d23",
X"893dfc05",
X"53765279",
X"51f8da3f",
X"83c08008",
X"81ff0670",
X"57557496",
X"387c547b",
X"53883d22",
X"527651fd",
X"e53f83c0",
X"800881ff",
X"06567583",
X"c0800c89",
X"3d0d04f0",
X"3d0d6266",
X"02880580",
X"ce052241",
X"5d5e8002",
X"840580d2",
X"05227f81",
X"0533ff11",
X"5a5d5a5d",
X"81da5876",
X"bf2680e9",
X"3878802e",
X"80e1387a",
X"58787b27",
X"83387858",
X"821e3370",
X"872a585a",
X"76923d34",
X"923dfc05",
X"5677557b",
X"547e537d",
X"33528251",
X"f8de3f83",
X"c0800881",
X"ff065d80",
X"0b923d33",
X"585a7680",
X"2e833881",
X"5a821e33",
X"80ff067a",
X"872b0757",
X"76821f34",
X"7c913878",
X"78317083",
X"ffff0679",
X"1e5e5a57",
X"ff9b397c",
X"587783c0",
X"800c923d",
X"0d04f83d",
X"0d7b0284",
X"05b20522",
X"5858800b",
X"8a3d238a",
X"3dfc0553",
X"77527a51",
X"f6f73f83",
X"c0800881",
X"ff067057",
X"55749638",
X"7d547653",
X"893d2252",
X"7751feaf",
X"3f83c080",
X"0881ff06",
X"567583c0",
X"800c8a3d",
X"0d04ec3d",
X"0d666e02",
X"880580df",
X"0533028c",
X"0580e305",
X"33029005",
X"80e70533",
X"02940580",
X"eb053302",
X"980580ee",
X"05224143",
X"415f5c40",
X"570280f2",
X"0522963d",
X"23963df0",
X"05538417",
X"70537752",
X"59f6863f",
X"83c08008",
X"81ff0658",
X"7781e538",
X"777a8180",
X"06584080",
X"77258338",
X"81407994",
X"3d347b02",
X"840580c9",
X"05347c02",
X"840580ca",
X"05347d02",
X"840580cb",
X"05347a95",
X"3d347a88",
X"2a577602",
X"840580cd",
X"0534953d",
X"22577602",
X"840580ce",
X"05347688",
X"2a577602",
X"840580cf",
X"05347792",
X"3d34963d",
X"ec115757",
X"8855f417",
X"54923d22",
X"53775277",
X"51f6953f",
X"83c08008",
X"81ff0658",
X"7780ed38",
X"7e802e80",
X"cb38923d",
X"22790858",
X"587f802e",
X"9c387681",
X"80800779",
X"0c7e5496",
X"3dfc0553",
X"7783ffff",
X"06527851",
X"f9fc3f99",
X"39768280",
X"8007790c",
X"7e54953d",
X"22537783",
X"ffff0652",
X"7851fc8f",
X"3f83c080",
X"0881ff06",
X"58779d38",
X"923d2253",
X"80527f30",
X"70802584",
X"71315351",
X"57f9873f",
X"83c08008",
X"81ff0658",
X"7783c080",
X"0c963d0d",
X"04f63d0d",
X"7c028405",
X"b705335b",
X"5b805880",
X"57805680",
X"55795485",
X"5380527a",
X"51fda33f",
X"83c08008",
X"81ff0659",
X"78853879",
X"871c3478",
X"83c0800c",
X"8c3d0d04",
X"f93d0d02",
X"a7053302",
X"8405ab05",
X"33028805",
X"af053358",
X"5957800b",
X"83c8df33",
X"54547274",
X"2e9f3881",
X"147081ff",
X"06555373",
X"872681b6",
X"387381c4",
X"2983c8dc",
X"05831133",
X"515372e3",
X"387381c4",
X"2983c8d8",
X"0555800b",
X"87163476",
X"88163475",
X"8a163477",
X"89163480",
X"750c83c8",
X"d0088c16",
X"0c800b84",
X"1634880b",
X"85163480",
X"0b861634",
X"841508ff",
X"a1ff06a0",
X"80078416",
X"0c811470",
X"81ff0653",
X"537451fe",
X"bc3f83c0",
X"800881ff",
X"06705553",
X"7280cd38",
X"8a397308",
X"750c7254",
X"80c23972",
X"81eba855",
X"5681eba8",
X"08802eb2",
X"38758429",
X"14700876",
X"53700851",
X"5454722d",
X"83c08008",
X"81ff0653",
X"72802ece",
X"38811670",
X"81ff0681",
X"eba87184",
X"29115356",
X"57537208",
X"d0388054",
X"7383c080",
X"0c893d0d",
X"04f93d0d",
X"7957800b",
X"84180883",
X"c8d00c58",
X"f08c3f88",
X"170883c0",
X"80082783",
X"ed38effe",
X"3f83c080",
X"08810588",
X"180c83c8",
X"d008b811",
X"337081ff",
X"06515154",
X"73812ea4",
X"38738124",
X"88387378",
X"2e8a38b8",
X"3973822e",
X"9538b139",
X"763381f0",
X"06547390",
X"2ea63891",
X"7734a139",
X"73587633",
X"81f00654",
X"73902e09",
X"81069138",
X"efac3f83",
X"c0800881",
X"c8058c18",
X"0ca07734",
X"80567581",
X"c42983c8",
X"df113355",
X"5573802e",
X"aa3883c8",
X"d8157008",
X"56547480",
X"2e9d3888",
X"1508802e",
X"96388c14",
X"0883c8d0",
X"082e0981",
X"06893873",
X"51881508",
X"54732d81",
X"167081ff",
X"06575487",
X"7627ffba",
X"38763354",
X"73b02e81",
X"993873b0",
X"248f3873",
X"912eab38",
X"73a02e80",
X"f53882a6",
X"397380d0",
X"2e81e438",
X"7380d024",
X"8b387380",
X"c02e8199",
X"38828f39",
X"7381802e",
X"81fb3882",
X"85398056",
X"7581c429",
X"83c8dc11",
X"83113356",
X"59557380",
X"2ea83883",
X"c8d81570",
X"08565474",
X"802e9b38",
X"8c140883",
X"c8d0082e",
X"0981068e",
X"38735184",
X"15085473",
X"2d800b83",
X"19348116",
X"7081ff06",
X"57548776",
X"27ffb938",
X"92773481",
X"b539edc6",
X"3f8c1708",
X"83c08008",
X"2781a738",
X"b0773481",
X"a13983c8",
X"d0085480",
X"0b8c1534",
X"83c8d008",
X"54840b88",
X"153480c0",
X"7734ed9a",
X"3f83c080",
X"08b2058c",
X"180c80fa",
X"39ed8b3f",
X"8c170883",
X"c0800827",
X"80ec3883",
X"c8d00854",
X"810b8c15",
X"3483c8d0",
X"0854800b",
X"88153483",
X"c8d00854",
X"880ba015",
X"34ecdf3f",
X"83c08008",
X"94058c18",
X"0c80d077",
X"34bc3983",
X"c8d008a0",
X"11337083",
X"2a708106",
X"51515555",
X"73802ea6",
X"38880ba0",
X"1634ecb2",
X"3f8c1708",
X"83c08008",
X"279438ff",
X"8077348e",
X"39775380",
X"528051fa",
X"8b3fff90",
X"773483c8",
X"d008a011",
X"3370832a",
X"70810651",
X"51555573",
X"802e8638",
X"880ba016",
X"34893d0d",
X"04f43d0d",
X"02bb0533",
X"028405bf",
X"05335d5d",
X"800b83c8",
X"dc0b83c8",
X"d80b8c11",
X"72718814",
X"755c5a5b",
X"5f5c595b",
X"58831533",
X"5372802e",
X"81883873",
X"33537c73",
X"2e098106",
X"80fc3881",
X"1433537b",
X"732e0981",
X"0680ef38",
X"750883c8",
X"d0082e09",
X"810680e2",
X"38805675",
X"81c42983",
X"c8e01170",
X"33831e33",
X"5b575553",
X"74782e09",
X"81069738",
X"83c8e413",
X"0879082e",
X"0981068a",
X"38811433",
X"527451fe",
X"f83f8116",
X"7081ff06",
X"57538776",
X"27c53880",
X"77085454",
X"72742e91",
X"38765184",
X"13085372",
X"2d83c080",
X"0881ff06",
X"54800b83",
X"1b347353",
X"a9398118",
X"81c41681",
X"c41681c4",
X"1981c41f",
X"81c41e81",
X"c41d6081",
X"c405415d",
X"5e5f5956",
X"56588778",
X"25feca38",
X"80537283",
X"c0800c8e",
X"3d0d04f8",
X"3d0d02ae",
X"05227d59",
X"57805681",
X"55805486",
X"53818052",
X"7a51f4ee",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8a3d0d04",
X"f73d0d02",
X"b2052202",
X"8405b705",
X"33605a5b",
X"57805682",
X"55795486",
X"53818052",
X"7b51f4be",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8b3d0d04",
X"f83d0d02",
X"af053359",
X"80588057",
X"80568055",
X"78548953",
X"80527a51",
X"f4943f83",
X"c0800881",
X"ff0683c0",
X"800c8a3d",
X"0d04ffb8",
X"3d0d80cb",
X"3d087053",
X"81ea9452",
X"56febc92",
X"3f83c080",
X"0880f338",
X"7551feb5",
X"fd3f83ff",
X"ff0b83c0",
X"80082580",
X"e1387551",
X"feb5fc3f",
X"83c08008",
X"5583c080",
X"0880cf38",
X"82805383",
X"c0800852",
X"8a3d7052",
X"57fef9bb",
X"3f745275",
X"51feb4ec",
X"3f805980",
X"ca3dfdfc",
X"05548280",
X"53765275",
X"51feb2f2",
X"3f811555",
X"7488802e",
X"098106e1",
X"38805275",
X"51feb4c4",
X"3f800b83",
X"d4fc0c75",
X"83d4f80c",
X"8739800b",
X"83d4f80c",
X"80ca3d0d",
X"04ff3d0d",
X"73700853",
X"51029305",
X"33723470",
X"08810571",
X"0c833d0d",
X"04ffb83d",
X"0d80cb3d",
X"70708405",
X"52085856",
X"83d4f808",
X"802e80fa",
X"388a3d70",
X"5a765577",
X"5481d8c5",
X"5380cb3d",
X"fdfc0552",
X"55fee190",
X"3f805280",
X"ca3dfdfc",
X"0551ffad",
X"3f83d4fc",
X"085283d4",
X"f80851fe",
X"b3ca3f80",
X"587451fe",
X"ded23f80",
X"ca3dfdf8",
X"055483c0",
X"80085374",
X"5283d4f8",
X"0851feb1",
X"c53f83d4",
X"fc081883",
X"d4fc0c80",
X"ca3dfdf8",
X"05548153",
X"81eaa052",
X"83d4f808",
X"51feb1a6",
X"3f83d4fc",
X"081883d4",
X"fc0c80ca",
X"3d0d0483",
X"c08c0802",
X"83c08c0c",
X"fd3d0d80",
X"5383c08c",
X"088c0508",
X"5283c08c",
X"08880508",
X"5183d43f",
X"83c08008",
X"7083c080",
X"0c54853d",
X"0d83c08c",
X"0c0483c0",
X"8c080283",
X"c08c0cfd",
X"3d0d8153",
X"83c08c08",
X"8c050852",
X"83c08c08",
X"88050851",
X"83a13f83",
X"c0800870",
X"83c0800c",
X"54853d0d",
X"83c08c0c",
X"0483c08c",
X"080283c0",
X"8c0cf93d",
X"0d800b83",
X"c08c08fc",
X"050c83c0",
X"8c088805",
X"088025b9",
X"3883c08c",
X"08880508",
X"3083c08c",
X"0888050c",
X"800b83c0",
X"8c08f405",
X"0c83c08c",
X"08fc0508",
X"8a38810b",
X"83c08c08",
X"f4050c83",
X"c08c08f4",
X"050883c0",
X"8c08fc05",
X"0c83c08c",
X"088c0508",
X"8025b938",
X"83c08c08",
X"8c050830",
X"83c08c08",
X"8c050c80",
X"0b83c08c",
X"08f0050c",
X"83c08c08",
X"fc05088a",
X"38810b83",
X"c08c08f0",
X"050c83c0",
X"8c08f005",
X"0883c08c",
X"08fc050c",
X"805383c0",
X"8c088c05",
X"085283c0",
X"8c088805",
X"085181df",
X"3f83c080",
X"087083c0",
X"8c08f805",
X"0c5483c0",
X"8c08fc05",
X"08802e90",
X"3883c08c",
X"08f80508",
X"3083c08c",
X"08f8050c",
X"83c08c08",
X"f8050870",
X"83c0800c",
X"54893d0d",
X"83c08c0c",
X"0483c08c",
X"080283c0",
X"8c0cfb3d",
X"0d800b83",
X"c08c08fc",
X"050c83c0",
X"8c088805",
X"08802599",
X"3883c08c",
X"08880508",
X"3083c08c",
X"0888050c",
X"810b83c0",
X"8c08fc05",
X"0c83c08c",
X"088c0508",
X"80259038",
X"83c08c08",
X"8c050830",
X"83c08c08",
X"8c050c81",
X"5383c08c",
X"088c0508",
X"5283c08c",
X"08880508",
X"51bd3f83",
X"c0800870",
X"83c08c08",
X"f8050c54",
X"83c08c08",
X"fc050880",
X"2e903883",
X"c08c08f8",
X"05083083",
X"c08c08f8",
X"050c83c0",
X"8c08f805",
X"087083c0",
X"800c5487",
X"3d0d83c0",
X"8c0c0483",
X"c08c0802",
X"83c08c0c",
X"fd3d0d81",
X"0b83c08c",
X"08fc050c",
X"800b83c0",
X"8c08f805",
X"0c83c08c",
X"088c0508",
X"83c08c08",
X"88050827",
X"b93883c0",
X"8c08fc05",
X"08802eae",
X"38800b83",
X"c08c088c",
X"050824a2",
X"3883c08c",
X"088c0508",
X"1083c08c",
X"088c050c",
X"83c08c08",
X"fc050810",
X"83c08c08",
X"fc050cff",
X"b83983c0",
X"8c08fc05",
X"08802e80",
X"e13883c0",
X"8c088c05",
X"0883c08c",
X"08880508",
X"26ad3883",
X"c08c0888",
X"050883c0",
X"8c088c05",
X"083183c0",
X"8c088805",
X"0c83c08c",
X"08f80508",
X"83c08c08",
X"fc050807",
X"83c08c08",
X"f8050c83",
X"c08c08fc",
X"0508812a",
X"83c08c08",
X"fc050c83",
X"c08c088c",
X"0508812a",
X"83c08c08",
X"8c050cff",
X"953983c0",
X"8c089005",
X"08802e93",
X"3883c08c",
X"08880508",
X"7083c08c",
X"08f4050c",
X"51913983",
X"c08c08f8",
X"05087083",
X"c08c08f4",
X"050c5183",
X"c08c08f4",
X"050883c0",
X"800c853d",
X"0d83c08c",
X"0c0483c0",
X"8c080283",
X"c08c0cff",
X"3d0d800b",
X"83c08c08",
X"fc050c83",
X"c08c0888",
X"05088106",
X"ff117009",
X"7083c08c",
X"088c0508",
X"0683c08c",
X"08fc0508",
X"1183c08c",
X"08fc050c",
X"83c08c08",
X"88050881",
X"2a83c08c",
X"0888050c",
X"83c08c08",
X"8c050810",
X"83c08c08",
X"8c050c51",
X"51515183",
X"c08c0888",
X"0508802e",
X"8438ffab",
X"3983c08c",
X"08fc0508",
X"7083c080",
X"0c51833d",
X"0d83c08c",
X"0c04fc3d",
X"0d767079",
X"7b555555",
X"558f7227",
X"8c387275",
X"07830651",
X"70802ea9",
X"38ff1252",
X"71ff2e98",
X"38727081",
X"05543374",
X"70810556",
X"34ff1252",
X"71ff2e09",
X"8106ea38",
X"7483c080",
X"0c863d0d",
X"04745172",
X"70840554",
X"08717084",
X"05530c72",
X"70840554",
X"08717084",
X"05530c72",
X"70840554",
X"08717084",
X"05530c72",
X"70840554",
X"08717084",
X"05530cf0",
X"1252718f",
X"26c93883",
X"72279538",
X"72708405",
X"54087170",
X"8405530c",
X"fc125271",
X"8326ed38",
X"7054ff81",
X"39000000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"70704740",
X"0c704268",
X"0c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"0000309d",
X"000030de",
X"000030fe",
X"00003122",
X"0000312e",
X"00003138",
X"00003cb0",
X"000046e3",
X"000047ac",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3a00",
X"0c0c3b00",
X"0a0a0005",
X"0b0b0005",
X"06060005",
X"07070004",
X"04044500",
X"05054400",
X"0e0f2900",
X"08080004",
X"09090004",
X"0a0f4300",
X"090f4200",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"000058dd",
X"00005be4",
X"000059f0",
X"00005be4",
X"00005a2d",
X"00005a7e",
X"00005abd",
X"00005ac6",
X"00005be4",
X"00005be4",
X"00005be4",
X"00005be4",
X"00005acf",
X"00005ad7",
X"00005ade",
X"00005ce4",
X"00005ddd",
X"00005ef1",
X"000061e3",
X"000061fe",
X"000061ea",
X"000061fe",
X"00006205",
X"00006210",
X"00006217",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"41545800",
X"63686f6f",
X"73652000",
X"66696c65",
X"20202573",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"25782e48",
X"75622e20",
X"25642070",
X"6f727473",
X"00000000",
X"25782e48",
X"49440000",
X"204d6f75",
X"73650000",
X"204b6579",
X"626f6172",
X"64000000",
X"204a6f79",
X"73746963",
X"6b3a2564",
X"00000000",
X"31364b00",
X"556e6b6e",
X"6f776e20",
X"74797065",
X"206f6620",
X"63617274",
X"72696467",
X"65210000",
X"41353200",
X"43415200",
X"42494e00",
X"31366b20",
X"63617274",
X"20747970",
X"65000000",
X"4c656674",
X"20666f72",
X"206f6e65",
X"20636869",
X"70000000",
X"52696768",
X"7420666f",
X"72207477",
X"6f206368",
X"69700000",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a257300",
X"526f7461",
X"74652055",
X"5342206a",
X"6f797374",
X"69636b73",
X"00000000",
X"45786974",
X"00000000",
X"35323030",
X"2e726f6d",
X"00000000",
X"524f4d00",
X"4d454d00",
X"2f757362",
X"2e6c6f67",
X"00000000",
X"0a000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"01000000",
X"00000000",
X"00007394",
X"000071e4",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"35323030",
X"00000000",
X"2f617461",
X"72353230",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
