-- megafunction wizard: %ALTREMOTE_UPDATE%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altremote_update 

-- ============================================================
-- File Name: remote_update.vhd
-- Megafunction Name(s):
-- 			altremote_update
--
-- Simulation Library Files(s):
-- 			cycloneive;lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altremote_update CBX_AUTO_BLACKBOX="ALL" check_app_pof="false" DEVICE_FAMILY="Cyclone IV E" in_data_width=22 operation_mode="remote" out_data_width=29 busy clock data_in data_out param read_param read_source reconfig reset reset_timer write_param
--VERSION_BEGIN 13.0 cbx_altremote_update 2013:06:12:18:04:00:SJ cbx_cycloneii 2013:06:12:18:04:00:SJ cbx_lpm_add_sub 2013:06:12:18:04:00:SJ cbx_lpm_compare 2013:06:12:18:04:00:SJ cbx_lpm_counter 2013:06:12:18:04:00:SJ cbx_lpm_decode 2013:06:12:18:04:00:SJ cbx_lpm_shiftreg 2013:06:12:18:04:00:SJ cbx_mgl 2013:06:12:18:04:42:SJ cbx_stratix 2013:06:12:18:04:00:SJ cbx_stratixii 2013:06:12:18:04:00:SJ  VERSION_END

 LIBRARY cycloneive;
 USE cycloneive.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = cycloneive_rublock 1 lpm_counter 2 reg 61 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  remote_update_rmtupdt_51n IS 
	 PORT 
	 ( 
		 busy	:	OUT  STD_LOGIC;
		 clock	:	IN  STD_LOGIC;
		 data_in	:	IN  STD_LOGIC_VECTOR (21 DOWNTO 0) := (OTHERS => '0');
		 data_out	:	OUT  STD_LOGIC_VECTOR (28 DOWNTO 0);
		 param	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0');
		 read_param	:	IN  STD_LOGIC := '0';
		 read_source	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0) := (OTHERS => '0');
		 reconfig	:	IN  STD_LOGIC := '0';
		 reset	:	IN  STD_LOGIC;
		 reset_timer	:	IN  STD_LOGIC := '0';
		 write_param	:	IN  STD_LOGIC := '0'
	 ); 
 END remote_update_rmtupdt_51n;

 ARCHITECTURE RTL OF remote_update_rmtupdt_51n IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "suppress_da_rule_internal=c104;suppress_da_rule_internal=C101;suppress_da_rule_internal=C103";

	 SIGNAL	 check_busy_dffe	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe1a0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe1a1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dffe1a_ena	:	STD_LOGIC_VECTOR(1 DOWNTO 0);
	 SIGNAL	 dffe2a0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe2a1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe2a2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dffe2a_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL	 dffe3a0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe3a1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe3a2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dffe3a_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL	 dffe7a	:	STD_LOGIC_VECTOR(28 DOWNTO 0)
	 -- synopsys translate_off
	  := "00000000000000000000000000000"
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dffe7a_ena	:	STD_LOGIC_VECTOR(28 DOWNTO 0);
	 SIGNAL	 dffe8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe9a	:	STD_LOGIC_VECTOR(6 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dffe9a_ena	:	STD_LOGIC_VECTOR(6 DOWNTO 0);
	 SIGNAL	 idle_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 idle_write_wait	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_init_counter_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_init_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_post_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_pre_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_source_update_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_init_counter_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_init_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_load_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_post_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_pre_data_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_source_update_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 write_wait_state	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_cntr5_w_lg_w_q_range38w41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr5_w_lg_w_q_range39w40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr5_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cntr5_w_q_range38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr5_w_q_range39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr6_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_sd4_regout	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w807w810w813w816w818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w807w810w846w847w848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w807w827w828w829w830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w821w822w823w824w825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w821w822w823w891w892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w821w822w850w851w852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w821w855w856w857w858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w821w855w913w914w915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w832w833w881w882w883w884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w832w833w834w835w836w837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w832w833w834w905w906w907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w832w894w895w896w897w898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w832w894w917w918w919w920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w874w875w876w877w879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w874w900w901w902w903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w840w886w887w888w889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w840w841w842w843w844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w840w841w909w910w911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w860w868w869w870w871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w860w861w862w863w864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w804w807w810w813w816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w804w807w810w846w847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w804w807w827w828w829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w804w821w822w823w824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w804w821w822w823w891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w804w821w822w850w851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w804w821w855w856w857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w804w821w855w913w914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w832w833w881w882w883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w832w833w834w835w836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w832w833w834w905w906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w832w894w895w896w897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w832w894w917w918w919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w874w875w876w877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w874w900w901w902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w840w886w887w888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w840w841w842w843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w840w841w909w910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w860w868w869w870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w860w861w862w863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w804w807w810w813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w804w807w810w846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w804w807w827w828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w804w821w822w823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w804w821w822w850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w804w821w855w856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w804w821w855w913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w832w833w881w882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w832w833w834w835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w832w833w834w905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w832w894w895w896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w832w894w917w918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w874w875w876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w874w900w901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w840w886w887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w840w841w842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w840w841w909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w860w868w869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w860w861w862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w804w807w810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w804w807w827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w804w821w822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w804w821w855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w832w833w881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w832w833w834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w832w894w895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w832w894w917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w874w875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w874w900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w840w886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w840w841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w860w868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w860w861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w804w807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w804w821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w832w833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w832w894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_idle955w956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rsource_load12w13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rsource_load12w20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rsource_load12w24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rsource_load12w30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rsource_load12w34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable100w134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_source_update1013w1014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_data972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_init_counter968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_post978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_pre_data967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_load15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_load22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_load26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_load32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_load36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rublock_regout_reg1019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_data990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_init_counter987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_post_data996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_pre_data986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range800w873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range800w839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w4w_range1040w1041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w4w_range1044w1045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bit_counter_all_done989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bit_counter_param_start_match966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_data931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_init935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_init_counter933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_post930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_pre_data932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_source_update934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_load12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_update_done963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_select_shift_nloop1018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w1w954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w2w953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_width_counter_all_done970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_width_counter_param_width_match971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_data925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_init929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_init_counter928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_load923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_post_data924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_pre_data926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_source_update927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_wait922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_wsource_update_done983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range800w801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range802w803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range805w806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range808w809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range811w812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range814w815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range817w878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_idle955w956w957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w4w_range1040w1041w1042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w4w_range1044w1045w1046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable98w99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_source_update1013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_load17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_load8w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  bit_counter_all_done :	STD_LOGIC;
	 SIGNAL  bit_counter_clear :	STD_LOGIC;
	 SIGNAL  bit_counter_enable :	STD_LOGIC;
	 SIGNAL  bit_counter_param_start :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  bit_counter_param_start_match :	STD_LOGIC;
	 SIGNAL  combine_port :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  global_gnd :	STD_LOGIC;
	 SIGNAL  global_vcc :	STD_LOGIC;
	 SIGNAL  idle :	STD_LOGIC;
	 SIGNAL  param_decoder_param_latch :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  param_decoder_select :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  power_up :	STD_LOGIC;
	 SIGNAL  read_data :	STD_LOGIC;
	 SIGNAL  read_init :	STD_LOGIC;
	 SIGNAL  read_init_counter :	STD_LOGIC;
	 SIGNAL  read_post :	STD_LOGIC;
	 SIGNAL  read_pre_data :	STD_LOGIC;
	 SIGNAL  read_source_update :	STD_LOGIC;
	 SIGNAL  rsource_load :	STD_LOGIC;
	 SIGNAL  rsource_parallel_in :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  rsource_serial_out :	STD_LOGIC;
	 SIGNAL  rsource_shift_enable :	STD_LOGIC;
	 SIGNAL  rsource_state_par_ini :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rsource_update_done :	STD_LOGIC;
	 SIGNAL  rublock_captnupdt :	STD_LOGIC;
	 SIGNAL  rublock_clock :	STD_LOGIC;
	 SIGNAL  rublock_reconfig :	STD_LOGIC;
	 SIGNAL  rublock_reconfig_st :	STD_LOGIC;
	 SIGNAL  rublock_regin :	STD_LOGIC;
	 SIGNAL  rublock_regout :	STD_LOGIC;
	 SIGNAL  rublock_regout_reg :	STD_LOGIC;
	 SIGNAL  rublock_shiftnld :	STD_LOGIC;
	 SIGNAL  select_shift_nloop :	STD_LOGIC;
	 SIGNAL  shift_reg_clear :	STD_LOGIC;
	 SIGNAL  shift_reg_load_enable :	STD_LOGIC;
	 SIGNAL  shift_reg_serial_in :	STD_LOGIC;
	 SIGNAL  shift_reg_serial_out :	STD_LOGIC;
	 SIGNAL  shift_reg_shift_enable :	STD_LOGIC;
	 SIGNAL  start_bit_decoder_out :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  start_bit_decoder_param_select :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  w1w :	STD_LOGIC;
	 SIGNAL  w2w :	STD_LOGIC;
	 SIGNAL  w4w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  w52w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  w82w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  width_counter_all_done :	STD_LOGIC;
	 SIGNAL  width_counter_clear :	STD_LOGIC;
	 SIGNAL  width_counter_enable :	STD_LOGIC;
	 SIGNAL  width_counter_param_width :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  width_counter_param_width_match :	STD_LOGIC;
	 SIGNAL  width_decoder_out :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  width_decoder_param_select :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  write_data :	STD_LOGIC;
	 SIGNAL  write_init :	STD_LOGIC;
	 SIGNAL  write_init_counter :	STD_LOGIC;
	 SIGNAL  write_load :	STD_LOGIC;
	 SIGNAL  write_post_data :	STD_LOGIC;
	 SIGNAL  write_pre_data :	STD_LOGIC;
	 SIGNAL  write_source_update :	STD_LOGIC;
	 SIGNAL  write_wait :	STD_LOGIC;
	 SIGNAL  wsource_state_par_ini :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wsource_update_done :	STD_LOGIC;
	 SIGNAL  wire_w_data_in_range103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rsource_parallel_in_range14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rsource_state_par_ini_range21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rsource_state_par_ini_range25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w4w_range1040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w4w_range1044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_wsource_state_par_ini_range31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_wsource_state_par_ini_range35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  cycloneive_rublock
	 PORT
	 ( 
		captnupdt	:	IN STD_LOGIC;
		clk	:	IN STD_LOGIC;
		rconfig	:	IN STD_LOGIC;
		regin	:	IN STD_LOGIC;
		regout	:	OUT STD_LOGIC;
		rsttimer	:	IN STD_LOGIC;
		shiftnld	:	IN STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w807w810w813w816w818w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w804w807w810w813w816w(0) AND wire_w_param_decoder_param_latch_range817w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w807w810w846w847w848w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w804w807w810w846w847w(0) AND wire_w_param_decoder_param_latch_range817w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w807w827w828w829w830w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w804w807w827w828w829w(0) AND wire_w_param_decoder_param_latch_range817w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w821w822w823w824w825w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w804w821w822w823w824w(0) AND wire_w_param_decoder_param_latch_range817w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w821w822w823w891w892w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w804w821w822w823w891w(0) AND wire_w_lg_w_param_decoder_param_latch_range817w878w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w821w822w850w851w852w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w804w821w822w850w851w(0) AND wire_w_param_decoder_param_latch_range817w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w821w855w856w857w858w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w804w821w855w856w857w(0) AND wire_w_param_decoder_param_latch_range817w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w821w855w913w914w915w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w804w821w855w913w914w(0) AND wire_w_param_decoder_param_latch_range817w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w832w833w881w882w883w884w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w832w833w881w882w883w(0) AND wire_w_lg_w_param_decoder_param_latch_range817w878w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w832w833w834w835w836w837w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w832w833w834w835w836w(0) AND wire_w_param_decoder_param_latch_range817w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w832w833w834w905w906w907w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w832w833w834w905w906w(0) AND wire_w_param_decoder_param_latch_range817w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w832w894w895w896w897w898w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w832w894w895w896w897w(0) AND wire_w_lg_w_param_decoder_param_latch_range817w878w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w832w894w917w918w919w920w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w832w894w917w918w919w(0) AND wire_w_param_decoder_param_latch_range817w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w874w875w876w877w879w(0) <= wire_w_lg_w_lg_w_lg_w874w875w876w877w(0) AND wire_w_lg_w_param_decoder_param_latch_range817w878w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w874w900w901w902w903w(0) <= wire_w_lg_w_lg_w_lg_w874w900w901w902w(0) AND wire_w_param_decoder_param_latch_range817w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w840w886w887w888w889w(0) <= wire_w_lg_w_lg_w_lg_w840w886w887w888w(0) AND wire_w_lg_w_param_decoder_param_latch_range817w878w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w840w841w842w843w844w(0) <= wire_w_lg_w_lg_w_lg_w840w841w842w843w(0) AND wire_w_param_decoder_param_latch_range817w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w840w841w909w910w911w(0) <= wire_w_lg_w_lg_w_lg_w840w841w909w910w(0) AND wire_w_param_decoder_param_latch_range817w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w860w868w869w870w871w(0) <= wire_w_lg_w_lg_w_lg_w860w868w869w870w(0) AND wire_w_param_decoder_param_latch_range817w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w860w861w862w863w864w(0) <= wire_w_lg_w_lg_w_lg_w860w861w862w863w(0) AND wire_w_param_decoder_param_latch_range817w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w804w807w810w813w816w(0) <= wire_w_lg_w_lg_w_lg_w804w807w810w813w(0) AND wire_w_lg_w_param_decoder_param_latch_range814w815w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w804w807w810w846w847w(0) <= wire_w_lg_w_lg_w_lg_w804w807w810w846w(0) AND wire_w_lg_w_param_decoder_param_latch_range814w815w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w804w807w827w828w829w(0) <= wire_w_lg_w_lg_w_lg_w804w807w827w828w(0) AND wire_w_lg_w_param_decoder_param_latch_range814w815w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w804w821w822w823w824w(0) <= wire_w_lg_w_lg_w_lg_w804w821w822w823w(0) AND wire_w_lg_w_param_decoder_param_latch_range814w815w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w804w821w822w823w891w(0) <= wire_w_lg_w_lg_w_lg_w804w821w822w823w(0) AND wire_w_param_decoder_param_latch_range814w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w804w821w822w850w851w(0) <= wire_w_lg_w_lg_w_lg_w804w821w822w850w(0) AND wire_w_lg_w_param_decoder_param_latch_range814w815w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w804w821w855w856w857w(0) <= wire_w_lg_w_lg_w_lg_w804w821w855w856w(0) AND wire_w_lg_w_param_decoder_param_latch_range814w815w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w804w821w855w913w914w(0) <= wire_w_lg_w_lg_w_lg_w804w821w855w913w(0) AND wire_w_lg_w_param_decoder_param_latch_range814w815w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w832w833w881w882w883w(0) <= wire_w_lg_w_lg_w_lg_w832w833w881w882w(0) AND wire_w_param_decoder_param_latch_range814w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w832w833w834w835w836w(0) <= wire_w_lg_w_lg_w_lg_w832w833w834w835w(0) AND wire_w_lg_w_param_decoder_param_latch_range814w815w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w832w833w834w905w906w(0) <= wire_w_lg_w_lg_w_lg_w832w833w834w905w(0) AND wire_w_lg_w_param_decoder_param_latch_range814w815w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w832w894w895w896w897w(0) <= wire_w_lg_w_lg_w_lg_w832w894w895w896w(0) AND wire_w_param_decoder_param_latch_range814w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w832w894w917w918w919w(0) <= wire_w_lg_w_lg_w_lg_w832w894w917w918w(0) AND wire_w_lg_w_param_decoder_param_latch_range814w815w(0);
	wire_w_lg_w_lg_w_lg_w874w875w876w877w(0) <= wire_w_lg_w_lg_w874w875w876w(0) AND wire_w_param_decoder_param_latch_range814w(0);
	wire_w_lg_w_lg_w_lg_w874w900w901w902w(0) <= wire_w_lg_w_lg_w874w900w901w(0) AND wire_w_lg_w_param_decoder_param_latch_range814w815w(0);
	wire_w_lg_w_lg_w_lg_w840w886w887w888w(0) <= wire_w_lg_w_lg_w840w886w887w(0) AND wire_w_param_decoder_param_latch_range814w(0);
	wire_w_lg_w_lg_w_lg_w840w841w842w843w(0) <= wire_w_lg_w_lg_w840w841w842w(0) AND wire_w_lg_w_param_decoder_param_latch_range814w815w(0);
	wire_w_lg_w_lg_w_lg_w840w841w909w910w(0) <= wire_w_lg_w_lg_w840w841w909w(0) AND wire_w_lg_w_param_decoder_param_latch_range814w815w(0);
	wire_w_lg_w_lg_w_lg_w860w868w869w870w(0) <= wire_w_lg_w_lg_w860w868w869w(0) AND wire_w_lg_w_param_decoder_param_latch_range814w815w(0);
	wire_w_lg_w_lg_w_lg_w860w861w862w863w(0) <= wire_w_lg_w_lg_w860w861w862w(0) AND wire_w_lg_w_param_decoder_param_latch_range814w815w(0);
	wire_w_lg_w_lg_w_lg_w804w807w810w813w(0) <= wire_w_lg_w_lg_w804w807w810w(0) AND wire_w_lg_w_param_decoder_param_latch_range811w812w(0);
	wire_w_lg_w_lg_w_lg_w804w807w810w846w(0) <= wire_w_lg_w_lg_w804w807w810w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w804w807w827w828w(0) <= wire_w_lg_w_lg_w804w807w827w(0) AND wire_w_lg_w_param_decoder_param_latch_range811w812w(0);
	wire_w_lg_w_lg_w_lg_w804w821w822w823w(0) <= wire_w_lg_w_lg_w804w821w822w(0) AND wire_w_lg_w_param_decoder_param_latch_range811w812w(0);
	wire_w_lg_w_lg_w_lg_w804w821w822w850w(0) <= wire_w_lg_w_lg_w804w821w822w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w804w821w855w856w(0) <= wire_w_lg_w_lg_w804w821w855w(0) AND wire_w_lg_w_param_decoder_param_latch_range811w812w(0);
	wire_w_lg_w_lg_w_lg_w804w821w855w913w(0) <= wire_w_lg_w_lg_w804w821w855w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w832w833w881w882w(0) <= wire_w_lg_w_lg_w832w833w881w(0) AND wire_w_lg_w_param_decoder_param_latch_range811w812w(0);
	wire_w_lg_w_lg_w_lg_w832w833w834w835w(0) <= wire_w_lg_w_lg_w832w833w834w(0) AND wire_w_lg_w_param_decoder_param_latch_range811w812w(0);
	wire_w_lg_w_lg_w_lg_w832w833w834w905w(0) <= wire_w_lg_w_lg_w832w833w834w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w832w894w895w896w(0) <= wire_w_lg_w_lg_w832w894w895w(0) AND wire_w_lg_w_param_decoder_param_latch_range811w812w(0);
	wire_w_lg_w_lg_w_lg_w832w894w917w918w(0) <= wire_w_lg_w_lg_w832w894w917w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w874w875w876w(0) <= wire_w_lg_w874w875w(0) AND wire_w_lg_w_param_decoder_param_latch_range811w812w(0);
	wire_w_lg_w_lg_w874w900w901w(0) <= wire_w_lg_w874w900w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w840w886w887w(0) <= wire_w_lg_w840w886w(0) AND wire_w_lg_w_param_decoder_param_latch_range811w812w(0);
	wire_w_lg_w_lg_w840w841w842w(0) <= wire_w_lg_w840w841w(0) AND wire_w_lg_w_param_decoder_param_latch_range811w812w(0);
	wire_w_lg_w_lg_w840w841w909w(0) <= wire_w_lg_w840w841w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w860w868w869w(0) <= wire_w_lg_w860w868w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w860w861w862w(0) <= wire_w_lg_w860w861w(0) AND wire_w_lg_w_param_decoder_param_latch_range811w812w(0);
	wire_w_lg_w_lg_w804w807w810w(0) <= wire_w_lg_w804w807w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w804w807w827w(0) <= wire_w_lg_w804w807w(0) AND wire_w_param_decoder_param_latch_range808w(0);
	wire_w_lg_w_lg_w804w821w822w(0) <= wire_w_lg_w804w821w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w804w821w855w(0) <= wire_w_lg_w804w821w(0) AND wire_w_param_decoder_param_latch_range808w(0);
	wire_w_lg_w_lg_w832w833w881w(0) <= wire_w_lg_w832w833w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w832w833w834w(0) <= wire_w_lg_w832w833w(0) AND wire_w_param_decoder_param_latch_range808w(0);
	wire_w_lg_w_lg_w832w894w895w(0) <= wire_w_lg_w832w894w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w832w894w917w(0) <= wire_w_lg_w832w894w(0) AND wire_w_param_decoder_param_latch_range808w(0);
	wire_w_lg_w874w875w(0) <= wire_w874w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w874w900w(0) <= wire_w874w(0) AND wire_w_param_decoder_param_latch_range808w(0);
	wire_w_lg_w840w886w(0) <= wire_w840w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w840w841w(0) <= wire_w840w(0) AND wire_w_param_decoder_param_latch_range808w(0);
	wire_w_lg_w860w868w(0) <= wire_w860w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w860w861w(0) <= wire_w860w(0) AND wire_w_param_decoder_param_latch_range808w(0);
	wire_w_lg_w804w807w(0) <= wire_w804w(0) AND wire_w_lg_w_param_decoder_param_latch_range805w806w(0);
	wire_w_lg_w804w821w(0) <= wire_w804w(0) AND wire_w_param_decoder_param_latch_range805w(0);
	wire_w_lg_w832w833w(0) <= wire_w832w(0) AND wire_w_lg_w_param_decoder_param_latch_range805w806w(0);
	wire_w_lg_w832w894w(0) <= wire_w832w(0) AND wire_w_param_decoder_param_latch_range805w(0);
	wire_w_lg_w_lg_idle955w956w(0) <= wire_w_lg_idle955w(0) AND wire_w_lg_w2w953w(0);
	wire_w874w(0) <= wire_w_lg_w_param_decoder_param_latch_range800w873w(0) AND wire_w_lg_w_param_decoder_param_latch_range805w806w(0);
	wire_w840w(0) <= wire_w_lg_w_param_decoder_param_latch_range800w839w(0) AND wire_w_lg_w_param_decoder_param_latch_range805w806w(0);
	wire_w860w(0) <= wire_w_lg_w_param_decoder_param_latch_range800w839w(0) AND wire_w_param_decoder_param_latch_range805w(0);
	wire_w_lg_w_lg_rsource_load12w13w(0) <= wire_w_lg_rsource_load12w(0) AND dffe1a1;
	wire_w_lg_w_lg_rsource_load12w20w(0) <= wire_w_lg_rsource_load12w(0) AND dffe2a1;
	wire_w_lg_w_lg_rsource_load12w24w(0) <= wire_w_lg_rsource_load12w(0) AND dffe2a2;
	wire_w_lg_w_lg_rsource_load12w30w(0) <= wire_w_lg_rsource_load12w(0) AND dffe3a1;
	wire_w_lg_w_lg_rsource_load12w34w(0) <= wire_w_lg_rsource_load12w(0) AND dffe3a2;
	wire_w_lg_w_lg_shift_reg_load_enable100w102w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(1);
	wire_w_lg_w_lg_shift_reg_load_enable100w138w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(10);
	wire_w_lg_w_lg_shift_reg_load_enable100w142w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(11);
	wire_w_lg_w_lg_shift_reg_load_enable100w146w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(12);
	wire_w_lg_w_lg_shift_reg_load_enable100w150w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(13);
	wire_w_lg_w_lg_shift_reg_load_enable100w154w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(14);
	wire_w_lg_w_lg_shift_reg_load_enable100w158w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(15);
	wire_w_lg_w_lg_shift_reg_load_enable100w162w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(16);
	wire_w_lg_w_lg_shift_reg_load_enable100w166w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(17);
	wire_w_lg_w_lg_shift_reg_load_enable100w170w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(18);
	wire_w_lg_w_lg_shift_reg_load_enable100w174w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(19);
	wire_w_lg_w_lg_shift_reg_load_enable100w106w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(2);
	wire_w_lg_w_lg_shift_reg_load_enable100w178w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(20);
	wire_w_lg_w_lg_shift_reg_load_enable100w182w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(21);
	wire_w_lg_w_lg_shift_reg_load_enable100w186w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(22);
	wire_w_lg_w_lg_shift_reg_load_enable100w110w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(3);
	wire_w_lg_w_lg_shift_reg_load_enable100w114w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(4);
	wire_w_lg_w_lg_shift_reg_load_enable100w118w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(5);
	wire_w_lg_w_lg_shift_reg_load_enable100w122w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(6);
	wire_w_lg_w_lg_shift_reg_load_enable100w126w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(7);
	wire_w_lg_w_lg_shift_reg_load_enable100w130w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(8);
	wire_w_lg_w_lg_shift_reg_load_enable100w134w(0) <= wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(9);
	wire_w804w(0) <= wire_w_lg_w_param_decoder_param_latch_range800w801w(0) AND wire_w_lg_w_param_decoder_param_latch_range802w803w(0);
	wire_w832w(0) <= wire_w_lg_w_param_decoder_param_latch_range800w801w(0) AND wire_w_param_decoder_param_latch_range802w(0);
	wire_w_lg_w_lg_read_source_update1013w1014w(0) <= wire_w_lg_read_source_update1013w(0) AND rsource_serial_out;
	wire_w_lg_idle955w(0) <= idle AND wire_w_lg_w1w954w(0);
	wire_w_lg_read_data972w(0) <= read_data AND wire_w_lg_width_counter_param_width_match971w(0);
	wire_w_lg_read_init_counter968w(0) <= read_init_counter AND wire_w_lg_bit_counter_param_start_match966w(0);
	wire_w_lg_read_post978w(0) <= read_post AND wire_w_lg_width_counter_all_done970w(0);
	wire_w_lg_read_pre_data967w(0) <= read_pre_data AND wire_w_lg_bit_counter_param_start_match966w(0);
	wire_w_lg_rsource_load15w(0) <= rsource_load AND wire_w_rsource_parallel_in_range14w(0);
	wire_w_lg_rsource_load22w(0) <= rsource_load AND wire_w_rsource_state_par_ini_range21w(0);
	wire_w_lg_rsource_load26w(0) <= rsource_load AND wire_w_rsource_state_par_ini_range25w(0);
	wire_w_lg_rsource_load32w(0) <= rsource_load AND wire_w_wsource_state_par_ini_range31w(0);
	wire_w_lg_rsource_load36w(0) <= rsource_load AND wire_w_wsource_state_par_ini_range35w(0);
	wire_w_lg_rublock_regout_reg1019w(0) <= rublock_regout_reg AND wire_w_lg_select_shift_nloop1018w(0);
	wire_w_lg_shift_reg_load_enable104w(0) <= shift_reg_load_enable AND wire_w_data_in_range103w(0);
	wire_w_lg_shift_reg_load_enable144w(0) <= shift_reg_load_enable AND wire_w_data_in_range143w(0);
	wire_w_lg_shift_reg_load_enable148w(0) <= shift_reg_load_enable AND wire_w_data_in_range147w(0);
	wire_w_lg_shift_reg_load_enable152w(0) <= shift_reg_load_enable AND wire_w_data_in_range151w(0);
	wire_w_lg_shift_reg_load_enable156w(0) <= shift_reg_load_enable AND wire_w_data_in_range155w(0);
	wire_w_lg_shift_reg_load_enable160w(0) <= shift_reg_load_enable AND wire_w_data_in_range159w(0);
	wire_w_lg_shift_reg_load_enable164w(0) <= shift_reg_load_enable AND wire_w_data_in_range163w(0);
	wire_w_lg_shift_reg_load_enable168w(0) <= shift_reg_load_enable AND wire_w_data_in_range167w(0);
	wire_w_lg_shift_reg_load_enable172w(0) <= shift_reg_load_enable AND wire_w_data_in_range171w(0);
	wire_w_lg_shift_reg_load_enable176w(0) <= shift_reg_load_enable AND wire_w_data_in_range175w(0);
	wire_w_lg_shift_reg_load_enable180w(0) <= shift_reg_load_enable AND wire_w_data_in_range179w(0);
	wire_w_lg_shift_reg_load_enable108w(0) <= shift_reg_load_enable AND wire_w_data_in_range107w(0);
	wire_w_lg_shift_reg_load_enable184w(0) <= shift_reg_load_enable AND wire_w_data_in_range183w(0);
	wire_w_lg_shift_reg_load_enable188w(0) <= shift_reg_load_enable AND wire_w_data_in_range187w(0);
	wire_w_lg_shift_reg_load_enable112w(0) <= shift_reg_load_enable AND wire_w_data_in_range111w(0);
	wire_w_lg_shift_reg_load_enable116w(0) <= shift_reg_load_enable AND wire_w_data_in_range115w(0);
	wire_w_lg_shift_reg_load_enable120w(0) <= shift_reg_load_enable AND wire_w_data_in_range119w(0);
	wire_w_lg_shift_reg_load_enable124w(0) <= shift_reg_load_enable AND wire_w_data_in_range123w(0);
	wire_w_lg_shift_reg_load_enable128w(0) <= shift_reg_load_enable AND wire_w_data_in_range127w(0);
	wire_w_lg_shift_reg_load_enable132w(0) <= shift_reg_load_enable AND wire_w_data_in_range131w(0);
	wire_w_lg_shift_reg_load_enable136w(0) <= shift_reg_load_enable AND wire_w_data_in_range135w(0);
	wire_w_lg_shift_reg_load_enable140w(0) <= shift_reg_load_enable AND wire_w_data_in_range139w(0);
	wire_w_lg_write_data990w(0) <= write_data AND wire_w_lg_width_counter_param_width_match971w(0);
	wire_w_lg_write_init_counter987w(0) <= write_init_counter AND wire_w_lg_bit_counter_param_start_match966w(0);
	wire_w_lg_write_post_data996w(0) <= write_post_data AND wire_w_lg_bit_counter_all_done989w(0);
	wire_w_lg_write_pre_data986w(0) <= write_pre_data AND wire_w_lg_bit_counter_param_start_match966w(0);
	wire_w_lg_w_param_decoder_param_latch_range800w873w(0) <= wire_w_param_decoder_param_latch_range800w(0) AND wire_w_lg_w_param_decoder_param_latch_range802w803w(0);
	wire_w_lg_w_param_decoder_param_latch_range800w839w(0) <= wire_w_param_decoder_param_latch_range800w(0) AND wire_w_param_decoder_param_latch_range802w(0);
	wire_w_lg_w_w4w_range1040w1041w(0) <= wire_w_w4w_range1040w(0) AND w1w;
	wire_w_lg_w_w4w_range1044w1045w(0) <= wire_w_w4w_range1044w(0) AND w1w;
	wire_w_lg_bit_counter_all_done989w(0) <= NOT bit_counter_all_done;
	wire_w_lg_bit_counter_param_start_match966w(0) <= NOT bit_counter_param_start_match;
	wire_w_lg_idle936w(0) <= NOT idle;
	wire_w_lg_read_data931w(0) <= NOT read_data;
	wire_w_lg_read_init935w(0) <= NOT read_init;
	wire_w_lg_read_init_counter933w(0) <= NOT read_init_counter;
	wire_w_lg_read_post930w(0) <= NOT read_post;
	wire_w_lg_read_pre_data932w(0) <= NOT read_pre_data;
	wire_w_lg_read_source_update934w(0) <= NOT read_source_update;
	wire_w_lg_rsource_load12w(0) <= NOT rsource_load;
	wire_w_lg_rsource_update_done963w(0) <= NOT rsource_update_done;
	wire_w_lg_select_shift_nloop1018w(0) <= NOT select_shift_nloop;
	wire_w_lg_shift_reg_load_enable100w(0) <= NOT shift_reg_load_enable;
	wire_w_lg_w1w954w(0) <= NOT w1w;
	wire_w_lg_w2w953w(0) <= NOT w2w;
	wire_w_lg_width_counter_all_done970w(0) <= NOT width_counter_all_done;
	wire_w_lg_width_counter_param_width_match971w(0) <= NOT width_counter_param_width_match;
	wire_w_lg_write_data925w(0) <= NOT write_data;
	wire_w_lg_write_init929w(0) <= NOT write_init;
	wire_w_lg_write_init_counter928w(0) <= NOT write_init_counter;
	wire_w_lg_write_load923w(0) <= NOT write_load;
	wire_w_lg_write_post_data924w(0) <= NOT write_post_data;
	wire_w_lg_write_pre_data926w(0) <= NOT write_pre_data;
	wire_w_lg_write_source_update927w(0) <= NOT write_source_update;
	wire_w_lg_write_wait922w(0) <= NOT write_wait;
	wire_w_lg_wsource_update_done983w(0) <= NOT wsource_update_done;
	wire_w_lg_w_param_decoder_param_latch_range800w801w(0) <= NOT wire_w_param_decoder_param_latch_range800w(0);
	wire_w_lg_w_param_decoder_param_latch_range802w803w(0) <= NOT wire_w_param_decoder_param_latch_range802w(0);
	wire_w_lg_w_param_decoder_param_latch_range805w806w(0) <= NOT wire_w_param_decoder_param_latch_range805w(0);
	wire_w_lg_w_param_decoder_param_latch_range808w809w(0) <= NOT wire_w_param_decoder_param_latch_range808w(0);
	wire_w_lg_w_param_decoder_param_latch_range811w812w(0) <= NOT wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_param_decoder_param_latch_range814w815w(0) <= NOT wire_w_param_decoder_param_latch_range814w(0);
	wire_w_lg_w_param_decoder_param_latch_range817w878w(0) <= NOT wire_w_param_decoder_param_latch_range817w(0);
	wire_w_lg_w_lg_w_lg_idle955w956w957w(0) <= wire_w_lg_w_lg_idle955w956w(0) OR write_wait;
	wire_w_lg_w_lg_w_w4w_range1040w1041w1042w(0) <= wire_w_lg_w_w4w_range1040w1041w(0) OR w2w;
	wire_w_lg_w_lg_w_w4w_range1044w1045w1046w(0) <= wire_w_lg_w_w4w_range1044w1045w(0) OR w2w;
	wire_w_lg_w_lg_shift_reg_load_enable98w99w(0) <= wire_w_lg_shift_reg_load_enable98w(0) OR shift_reg_clear;
	wire_w_lg_read_source_update1013w(0) <= read_source_update OR write_source_update;
	wire_w_lg_rsource_load17w(0) <= rsource_load OR global_vcc;
	wire_w_lg_rsource_load8w(0) <= rsource_load OR rsource_shift_enable;
	wire_w_lg_shift_reg_load_enable98w(0) <= shift_reg_load_enable OR shift_reg_shift_enable;
	bit_counter_all_done <= ((((wire_cntr5_w_lg_w_q_range38w41w(0) AND (NOT wire_cntr5_q(2))) AND wire_cntr5_q(3)) AND (NOT wire_cntr5_q(4))) AND wire_cntr5_q(5));
	bit_counter_clear <= (rsource_update_done OR wsource_update_done);
	bit_counter_enable <= (((((((((rsource_update_done OR wsource_update_done) OR read_init_counter) OR write_init_counter) OR read_pre_data) OR write_pre_data) OR read_data) OR write_data) OR read_post) OR write_post_data);
	bit_counter_param_start <= start_bit_decoder_out;
	bit_counter_param_start_match <= ((((((NOT w52w(0)) AND (NOT w52w(1))) AND (NOT w52w(2))) AND (NOT w52w(3))) AND (NOT w52w(4))) AND (NOT w52w(5)));
	busy <= wire_w_lg_idle936w(0);
	combine_port <= ( read_param & write_param & read_source & param);
	data_out <= dffe7a;
	global_gnd <= '0';
	global_vcc <= '1';
	idle <= idle_state;
	param_decoder_param_latch <= dffe9a;
	param_decoder_select <= ( wire_w_lg_w_lg_w_lg_w_lg_w_lg_w832w894w917w918w919w920w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w821w855w913w914w915w & wire_w_lg_w_lg_w_lg_w_lg_w840w841w909w910w911w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w832w833w834w905w906w907w & wire_w_lg_w_lg_w_lg_w_lg_w874w900w901w902w903w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w832w894w895w896w897w898w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w821w822w823w891w892w & wire_w_lg_w_lg_w_lg_w_lg_w840w886w887w888w889w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w832w833w881w882w883w884w & wire_w_lg_w_lg_w_lg_w_lg_w874w875w876w877w879w & wire_w_lg_w_lg_w_lg_w_lg_w860w868w869w870w871w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w821w822w850w851w852w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w807w810w846w847w848w & wire_w_lg_w_lg_w_lg_w_lg_w860w861w862w863w864w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w821w855w856w857w858w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w807w827w828w829w830w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w821w822w850w851w852w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w807w810w846w847w848w & wire_w_lg_w_lg_w_lg_w_lg_w840w841w842w843w844w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w832w833w834w835w836w837w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w807w827w828w829w830w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w821w822w823w824w825w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w804w807w810w813w816w818w);
	power_up <= ((((((((((((((wire_w_lg_idle936w(0) AND wire_w_lg_read_init935w(0)) AND wire_w_lg_read_source_update934w(0)) AND wire_w_lg_read_init_counter933w(0)) AND wire_w_lg_read_pre_data932w(0)) AND wire_w_lg_read_data931w(0)) AND wire_w_lg_read_post930w(0)) AND wire_w_lg_write_init929w(0)) AND wire_w_lg_write_init_counter928w(0)) AND wire_w_lg_write_source_update927w(0)) AND wire_w_lg_write_pre_data926w(0)) AND wire_w_lg_write_data925w(0)) AND wire_w_lg_write_post_data924w(0)) AND wire_w_lg_write_load923w(0)) AND wire_w_lg_write_wait922w(0));
	read_data <= read_data_state;
	read_init <= read_init_state;
	read_init_counter <= read_init_counter_state;
	read_post <= read_post_state;
	read_pre_data <= read_pre_data_state;
	read_source_update <= read_source_update_state;
	rsource_load <= (idle AND (write_param OR read_param));
	rsource_parallel_in <= ( wire_w_lg_w_lg_w_w4w_range1044w1045w1046w & wire_w_lg_w_lg_w_w4w_range1040w1041w1042w);
	rsource_serial_out <= dffe1a0;
	rsource_shift_enable <= wire_w_lg_read_source_update1013w(0);
	rsource_state_par_ini <= ( read_param & global_gnd & global_gnd);
	rsource_update_done <= dffe2a0;
	rublock_captnupdt <= wire_w_lg_write_load923w(0);
	rublock_clock <= (NOT (clock OR idle_write_wait));
	rublock_reconfig <= rublock_reconfig_st;
	rublock_reconfig_st <= (idle AND reconfig);
	rublock_regin <= ((((wire_w_lg_rublock_regout_reg1019w(0) AND wire_w_lg_read_source_update934w(0)) AND wire_w_lg_write_source_update927w(0)) OR (((shift_reg_serial_out AND select_shift_nloop) AND wire_w_lg_read_source_update934w(0)) AND wire_w_lg_write_source_update927w(0))) OR wire_w_lg_w_lg_read_source_update1013w1014w(0));
	rublock_regout <= wire_sd4_regout;
	rublock_regout_reg <= dffe8;
	rublock_shiftnld <= (((((((read_pre_data OR write_pre_data) OR read_data) OR write_data) OR read_post) OR write_post_data) OR read_source_update) OR write_source_update);
	select_shift_nloop <= (wire_w_lg_read_data972w(0) OR wire_w_lg_write_data990w(0));
	shift_reg_clear <= rsource_update_done;
	shift_reg_load_enable <= (idle AND write_param);
	shift_reg_serial_in <= (rublock_regout_reg AND select_shift_nloop);
	shift_reg_serial_out <= dffe7a(0);
	shift_reg_shift_enable <= (((read_data OR write_data) OR read_post) OR write_post_data);
	start_bit_decoder_out <= ((((((((((((((((((((((( "0" & start_bit_decoder_param_select(0) & start_bit_decoder_param_select(0) & start_bit_decoder_param_select(0) & start_bit_decoder_param_select(0) & "0") OR ( "0" & "0" & "0" & "0" & "0" & "0")) OR ( "0" & start_bit_decoder_param_select(2) & start_bit_decoder_param_select(2) & start_bit_decoder_param_select(2) & start_bit_decoder_param_select(2) & "0")) OR ( "0" & "0" & "0" & "0" & "0" & "0")) OR ( "0" & start_bit_decoder_param_select(4) & start_bit_decoder_param_select(4) & start_bit_decoder_param_select(4) & "0" & start_bit_decoder_param_select(4))) OR ( "0" & start_bit_decoder_param_select(5) & start_bit_decoder_param_select(5) & start_bit_decoder_param_select(5) & start_bit_decoder_param_select(5) & "0")) OR ( "0" & "0" & "0" & "0" & "0" & "0")) OR ( "0" & start_bit_decoder_param_select(7) & start_bit_decoder_param_select(7) & "0" & "0" & "0")) OR ( "0" & "0" & "0" & "0" & "0" & "0")) OR ( "0" & start_bit_decoder_param_select(9) & start_bit_decoder_param_select(9) & "0" & start_bit_decoder_param_select(9) & "0")) OR ( "0" & start_bit_decoder_param_select(10) & start_bit_decoder_param_select(10) & "0" & "0" & "0")) OR ( "0" & "0" & "0" & "0" & "0" & "0")) OR ( "0" & start_bit_decoder_param_select(12) & start_bit_decoder_param_select(12) & "0" & start_bit_decoder_param_select(12) & "0")) OR ( start_bit_decoder_param_select(13) & "0" & "0" & start_bit_decoder_param_select(13) & "0" & start_bit_decoder_param_select(13))) OR ( "0" & "0" & "0" & "0" & "0" & "0")) OR ( start_bit_decoder_param_select(15) & "0" & "0" & "0" & start_bit_decoder_param_select(15) & start_bit_decoder_param_select(15))) OR ( "0" & "0" & start_bit_decoder_param_select(16) & start_bit_decoder_param_select(16) & "0" & "0")) OR ( start_bit_decoder_param_select(17) & "0" & "0" & start_bit_decoder_param_select(17) & "0" & "0")) OR ( start_bit_decoder_param_select(18) & "0" & "0" & start_bit_decoder_param_select(18) & "0" & start_bit_decoder_param_select(18))) OR ( "0" & "0" & "0" & "0" & "0" & "0"
)) OR ( start_bit_decoder_param_select(20) & "0" & "0" & "0" & start_bit_decoder_param_select(20) & start_bit_decoder_param_select(20))) OR ( "0" & "0" & start_bit_decoder_param_select(21) & start_bit_decoder_param_select(21) & "0" & "0")) OR ( start_bit_decoder_param_select(22) & "0" & "0" & start_bit_decoder_param_select(22) & "0" & "0"));
	start_bit_decoder_param_select <= param_decoder_select;
	w1w <= read_param;
	w2w <= write_param;
	w4w <= read_source;
	w52w <= (wire_cntr5_q XOR bit_counter_param_start);
	w82w <= (wire_cntr6_q XOR width_counter_param_width);
	width_counter_all_done <= (((((NOT wire_cntr6_q(0)) AND (NOT wire_cntr6_q(1))) AND wire_cntr6_q(2)) AND wire_cntr6_q(3)) AND wire_cntr6_q(4));
	width_counter_clear <= (rsource_update_done OR wsource_update_done);
	width_counter_enable <= ((read_data OR write_data) OR read_post);
	width_counter_param_width <= width_decoder_out;
	width_counter_param_width_match <= (((((NOT w82w(0)) AND (NOT w82w(1))) AND (NOT w82w(2))) AND (NOT w82w(3))) AND (NOT w82w(4)));
	width_decoder_out <= ((((((((((((((((((((((( "0" & "0" & "0" & width_decoder_param_select(0) & "0") OR ( width_decoder_param_select(1) & width_decoder_param_select(1) & "0" & "0" & "0")) OR ( "0" & "0" & "0" & width_decoder_param_select(2) & "0")) OR ( width_decoder_param_select(3) & width_decoder_param_select(3) & width_decoder_param_select(3) & "0" & width_decoder_param_select(3))) OR ( "0" & "0" & "0" & "0" & width_decoder_param_select(4))) OR ( "0" & "0" & "0" & width_decoder_param_select(5) & "0")) OR ( width_decoder_param_select(6) & width_decoder_param_select(6) & "0" & "0" & "0")) OR ( "0" & "0" & "0" & width_decoder_param_select(7) & "0")) OR ( width_decoder_param_select(8) & width_decoder_param_select(8) & "0" & "0" & "0")) OR ( "0" & "0" & width_decoder_param_select(9) & "0" & width_decoder_param_select(9))) OR ( "0" & "0" & "0" & width_decoder_param_select(10) & "0")) OR ( width_decoder_param_select(11) & width_decoder_param_select(11) & "0" & "0" & "0")) OR ( "0" & "0" & width_decoder_param_select(12) & "0" & width_decoder_param_select(12))) OR ( "0" & "0" & "0" & "0" & width_decoder_param_select(13))) OR ( "0" & width_decoder_param_select(14) & width_decoder_param_select(14) & "0" & "0")) OR ( "0" & "0" & "0" & "0" & width_decoder_param_select(15))) OR ( width_decoder_param_select(16) & "0" & width_decoder_param_select(16) & width_decoder_param_select(16) & "0")) OR ( "0" & "0" & "0" & "0" & width_decoder_param_select(17))) OR ( "0" & "0" & "0" & "0" & width_decoder_param_select(18))) OR ( "0" & width_decoder_param_select(19) & width_decoder_param_select(19) & "0" & "0")) OR ( "0" & "0" & "0" & "0" & width_decoder_param_select(20))) OR ( width_decoder_param_select(21) & "0" & width_decoder_param_select(21) & width_decoder_param_select(21) & "0")) OR ( "0" & "0" & "0" & "0" & width_decoder_param_select(22)));
	width_decoder_param_select <= param_decoder_select;
	write_data <= write_data_state;
	write_init <= write_init_state;
	write_init_counter <= write_init_counter_state;
	write_load <= write_load_state;
	write_post_data <= write_post_data_state;
	write_pre_data <= write_pre_data_state;
	write_source_update <= write_source_update_state;
	write_wait <= write_wait_state;
	wsource_state_par_ini <= ( write_param & global_gnd & global_gnd);
	wsource_update_done <= dffe3a0;
	wire_w_data_in_range103w(0) <= data_in(0);
	wire_w_data_in_range143w(0) <= data_in(10);
	wire_w_data_in_range147w(0) <= data_in(11);
	wire_w_data_in_range151w(0) <= data_in(12);
	wire_w_data_in_range155w(0) <= data_in(13);
	wire_w_data_in_range159w(0) <= data_in(14);
	wire_w_data_in_range163w(0) <= data_in(15);
	wire_w_data_in_range167w(0) <= data_in(16);
	wire_w_data_in_range171w(0) <= data_in(17);
	wire_w_data_in_range175w(0) <= data_in(18);
	wire_w_data_in_range179w(0) <= data_in(19);
	wire_w_data_in_range107w(0) <= data_in(1);
	wire_w_data_in_range183w(0) <= data_in(20);
	wire_w_data_in_range187w(0) <= data_in(21);
	wire_w_data_in_range111w(0) <= data_in(2);
	wire_w_data_in_range115w(0) <= data_in(3);
	wire_w_data_in_range119w(0) <= data_in(4);
	wire_w_data_in_range123w(0) <= data_in(5);
	wire_w_data_in_range127w(0) <= data_in(6);
	wire_w_data_in_range131w(0) <= data_in(7);
	wire_w_data_in_range135w(0) <= data_in(8);
	wire_w_data_in_range139w(0) <= data_in(9);
	wire_w_param_decoder_param_latch_range800w(0) <= param_decoder_param_latch(0);
	wire_w_param_decoder_param_latch_range802w(0) <= param_decoder_param_latch(1);
	wire_w_param_decoder_param_latch_range805w(0) <= param_decoder_param_latch(2);
	wire_w_param_decoder_param_latch_range808w(0) <= param_decoder_param_latch(3);
	wire_w_param_decoder_param_latch_range811w(0) <= param_decoder_param_latch(4);
	wire_w_param_decoder_param_latch_range814w(0) <= param_decoder_param_latch(5);
	wire_w_param_decoder_param_latch_range817w(0) <= param_decoder_param_latch(6);
	wire_w_rsource_parallel_in_range14w(0) <= rsource_parallel_in(0);
	wire_w_rsource_state_par_ini_range21w(0) <= rsource_state_par_ini(0);
	wire_w_rsource_state_par_ini_range25w(0) <= rsource_state_par_ini(1);
	wire_w_w4w_range1040w(0) <= w4w(0);
	wire_w_w4w_range1044w(0) <= w4w(1);
	wire_w_wsource_state_par_ini_range31w(0) <= wsource_state_par_ini(0);
	wire_w_wsource_state_par_ini_range35w(0) <= wsource_state_par_ini(1);
	check_busy_dffe <= (OTHERS => '0');
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe1a0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe1a_ena(0) = '1') THEN dffe1a0 <= (wire_w_lg_rsource_load15w(0) OR wire_w_lg_w_lg_rsource_load12w13w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe1a1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe1a_ena(1) = '1') THEN dffe1a1 <= (rsource_parallel_in(1) AND rsource_load);
			END IF;
		END IF;
	END PROCESS;
	loop0 : FOR i IN 0 TO 1 GENERATE
		wire_dffe1a_ena(i) <= wire_w_lg_rsource_load8w(0);
	END GENERATE loop0;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe2a0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe2a_ena(0) = '1') THEN dffe2a0 <= (wire_w_lg_rsource_load22w(0) OR wire_w_lg_w_lg_rsource_load12w20w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe2a1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe2a_ena(1) = '1') THEN dffe2a1 <= (wire_w_lg_rsource_load26w(0) OR wire_w_lg_w_lg_rsource_load12w24w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe2a2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe2a_ena(2) = '1') THEN dffe2a2 <= (rsource_state_par_ini(2) AND rsource_load);
			END IF;
		END IF;
	END PROCESS;
	loop1 : FOR i IN 0 TO 2 GENERATE
		wire_dffe2a_ena(i) <= wire_w_lg_rsource_load17w(0);
	END GENERATE loop1;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe3a0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe3a_ena(0) = '1') THEN dffe3a0 <= (wire_w_lg_rsource_load32w(0) OR wire_w_lg_w_lg_rsource_load12w30w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe3a1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe3a_ena(1) = '1') THEN dffe3a1 <= (wire_w_lg_rsource_load36w(0) OR wire_w_lg_w_lg_rsource_load12w34w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe3a2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe3a_ena(2) = '1') THEN dffe3a2 <= (wsource_state_par_ini(2) AND rsource_load);
			END IF;
		END IF;
	END PROCESS;
	loop2 : FOR i IN 0 TO 2 GENERATE
		wire_dffe3a_ena(i) <= wire_w_lg_rsource_load17w(0);
	END GENERATE loop2;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(0) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(0) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(0) <= '0';
				ELSE dffe7a(0) <= (wire_w_lg_shift_reg_load_enable104w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w102w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(1) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(1) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(1) <= '0';
				ELSE dffe7a(1) <= (wire_w_lg_shift_reg_load_enable108w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w106w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(2) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(2) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(2) <= '0';
				ELSE dffe7a(2) <= (wire_w_lg_shift_reg_load_enable112w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w110w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(3) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(3) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(3) <= '0';
				ELSE dffe7a(3) <= (wire_w_lg_shift_reg_load_enable116w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w114w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(4) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(4) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(4) <= '0';
				ELSE dffe7a(4) <= (wire_w_lg_shift_reg_load_enable120w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w118w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(5) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(5) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(5) <= '0';
				ELSE dffe7a(5) <= (wire_w_lg_shift_reg_load_enable124w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w122w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(6) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(6) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(6) <= '0';
				ELSE dffe7a(6) <= (wire_w_lg_shift_reg_load_enable128w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w126w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(7) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(7) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(7) <= '0';
				ELSE dffe7a(7) <= (wire_w_lg_shift_reg_load_enable132w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w130w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(8) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(8) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(8) <= '0';
				ELSE dffe7a(8) <= (wire_w_lg_shift_reg_load_enable136w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w134w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(9) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(9) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(9) <= '0';
				ELSE dffe7a(9) <= (wire_w_lg_shift_reg_load_enable140w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w138w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(10) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(10) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(10) <= '0';
				ELSE dffe7a(10) <= (wire_w_lg_shift_reg_load_enable144w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w142w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(11) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(11) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(11) <= '0';
				ELSE dffe7a(11) <= (wire_w_lg_shift_reg_load_enable148w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w146w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(12) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(12) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(12) <= '0';
				ELSE dffe7a(12) <= (wire_w_lg_shift_reg_load_enable152w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w150w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(13) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(13) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(13) <= '0';
				ELSE dffe7a(13) <= (wire_w_lg_shift_reg_load_enable156w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w154w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(14) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(14) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(14) <= '0';
				ELSE dffe7a(14) <= (wire_w_lg_shift_reg_load_enable160w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w158w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(15) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(15) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(15) <= '0';
				ELSE dffe7a(15) <= (wire_w_lg_shift_reg_load_enable164w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w162w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(16) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(16) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(16) <= '0';
				ELSE dffe7a(16) <= (wire_w_lg_shift_reg_load_enable168w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w166w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(17) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(17) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(17) <= '0';
				ELSE dffe7a(17) <= (wire_w_lg_shift_reg_load_enable172w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w170w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(18) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(18) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(18) <= '0';
				ELSE dffe7a(18) <= (wire_w_lg_shift_reg_load_enable176w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w174w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(19) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(19) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(19) <= '0';
				ELSE dffe7a(19) <= (wire_w_lg_shift_reg_load_enable180w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w178w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(20) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(20) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(20) <= '0';
				ELSE dffe7a(20) <= (wire_w_lg_shift_reg_load_enable184w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w182w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(21) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(21) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(21) <= '0';
				ELSE dffe7a(21) <= (wire_w_lg_shift_reg_load_enable188w(0) OR wire_w_lg_w_lg_shift_reg_load_enable100w186w(0));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(22) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(22) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(22) <= '0';
				ELSE dffe7a(22) <= (wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(23));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(23) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(23) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(23) <= '0';
				ELSE dffe7a(23) <= (wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(24));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(24) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(24) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(24) <= '0';
				ELSE dffe7a(24) <= (wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(25));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(25) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(25) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(25) <= '0';
				ELSE dffe7a(25) <= (wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(26));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(26) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(26) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(26) <= '0';
				ELSE dffe7a(26) <= (wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(27));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(27) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(27) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(27) <= '0';
				ELSE dffe7a(27) <= (wire_w_lg_shift_reg_load_enable100w(0) AND dffe7a(28));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7a(28) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(28) = '1') THEN 
				IF (shift_reg_clear = '1') THEN dffe7a(28) <= '0';
				ELSE dffe7a(28) <= (wire_w_lg_shift_reg_load_enable100w(0) AND shift_reg_serial_in);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	loop3 : FOR i IN 0 TO 28 GENERATE
		wire_dffe7a_ena(i) <= wire_w_lg_w_lg_shift_reg_load_enable98w99w(0);
	END GENERATE loop3;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe8 <= rublock_regout;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe9a(0) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe9a_ena(0) = '1') THEN dffe9a(0) <= combine_port(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe9a(1) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe9a_ena(1) = '1') THEN dffe9a(1) <= combine_port(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe9a(2) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe9a_ena(2) = '1') THEN dffe9a(2) <= combine_port(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe9a(3) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe9a_ena(3) = '1') THEN dffe9a(3) <= combine_port(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe9a(4) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe9a_ena(4) = '1') THEN dffe9a(4) <= combine_port(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe9a(5) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe9a_ena(5) = '1') THEN dffe9a(5) <= combine_port(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe9a(6) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe9a_ena(6) = '1') THEN dffe9a(6) <= combine_port(6);
			END IF;
		END IF;
	END PROCESS;
	loop4 : FOR i IN 0 TO 6 GENERATE
		wire_dffe9a_ena(i) <= (idle AND (write_param OR read_param));
	END GENERATE loop4;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN idle_state <= '1';
		ELSIF (clock = '1' AND clock'event) THEN idle_state <= (((wire_w_lg_w_lg_w_lg_idle955w956w957w(0) OR (read_data AND width_counter_all_done)) OR (read_post AND width_counter_all_done)) OR power_up);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN idle_write_wait <= '0';
		ELSIF (clock = '1' AND clock'event) THEN idle_write_wait <= ((((wire_w_lg_w_lg_w_lg_idle955w956w957w(0) OR (read_data AND width_counter_all_done)) OR (read_post AND width_counter_all_done)) OR power_up) AND write_load);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_data_state <= (((read_init_counter AND bit_counter_param_start_match) OR (read_pre_data AND bit_counter_param_start_match)) OR (wire_w_lg_read_data972w(0) AND wire_w_lg_width_counter_all_done970w(0)));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_init_counter_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_init_counter_state <= rsource_update_done;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_init_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_init_state <= (idle AND read_param);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_post_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_post_state <= (((read_data AND width_counter_param_width_match) AND wire_w_lg_width_counter_all_done970w(0)) OR wire_w_lg_read_post978w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_pre_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_pre_data_state <= (wire_w_lg_read_init_counter968w(0) OR wire_w_lg_read_pre_data967w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN read_source_update_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN read_source_update_state <= ((read_init OR read_source_update) AND wire_w_lg_rsource_update_done963w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_data_state <= (((write_init_counter AND bit_counter_param_start_match) OR (write_pre_data AND bit_counter_param_start_match)) OR (wire_w_lg_write_data990w(0) AND wire_w_lg_bit_counter_all_done989w(0)));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_init_counter_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_init_counter_state <= wsource_update_done;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_init_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_init_state <= (idle AND write_param);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_load_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_load_state <= ((write_data AND bit_counter_all_done) OR (write_post_data AND bit_counter_all_done));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_post_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_post_data_state <= (((write_data AND width_counter_param_width_match) AND wire_w_lg_bit_counter_all_done989w(0)) OR wire_w_lg_write_post_data996w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_pre_data_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_pre_data_state <= (wire_w_lg_write_init_counter987w(0) OR wire_w_lg_write_pre_data986w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_source_update_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_source_update_state <= ((write_init OR write_source_update) AND wire_w_lg_wsource_update_done983w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN write_wait_state <= '0';
		ELSIF (clock = '1' AND clock'event) THEN write_wait_state <= write_load;
		END IF;
	END PROCESS;
	wire_cntr5_w_lg_w_q_range38w41w(0) <= wire_cntr5_w_q_range38w(0) AND wire_cntr5_w_lg_w_q_range39w40w(0);
	wire_cntr5_w_lg_w_q_range39w40w(0) <= NOT wire_cntr5_w_q_range39w(0);
	wire_cntr5_w_q_range38w(0) <= wire_cntr5_q(0);
	wire_cntr5_w_q_range39w(0) <= wire_cntr5_q(1);
	cntr5 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 6
	  )
	  PORT MAP ( 
		aclr => reset,
		clock => clock,
		cnt_en => bit_counter_enable,
		q => wire_cntr5_q,
		sclr => bit_counter_clear
	  );
	cntr6 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 5
	  )
	  PORT MAP ( 
		aclr => reset,
		clock => clock,
		cnt_en => width_counter_enable,
		q => wire_cntr6_q,
		sclr => width_counter_clear
	  );
	sd4 :  cycloneive_rublock
	  PORT MAP ( 
		captnupdt => rublock_captnupdt,
		clk => rublock_clock,
		rconfig => rublock_reconfig,
		regin => rublock_regin,
		regout => wire_sd4_regout,
		rsttimer => reset_timer,
		shiftnld => rublock_shiftnld
	  );

 END RTL; --remote_update_rmtupdt_51n
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY remote_update IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data_in		: IN STD_LOGIC_VECTOR (21 DOWNTO 0);
		param		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		read_param		: IN STD_LOGIC ;
		read_source		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		reconfig		: IN STD_LOGIC ;
		reset		: IN STD_LOGIC ;
		reset_timer		: IN STD_LOGIC ;
		write_param		: IN STD_LOGIC ;
		busy		: OUT STD_LOGIC ;
		data_out		: OUT STD_LOGIC_VECTOR (28 DOWNTO 0)
	);
END remote_update;


ARCHITECTURE RTL OF remote_update IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "altremote_update";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "check_app_pof=false;intended_device_family=Cyclone IV E;in_data_width=22;operation_mode=REMOTE;out_data_width=29;";
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (28 DOWNTO 0);



	COMPONENT remote_update_rmtupdt_51n
	PORT (
			clock	: IN STD_LOGIC ;
			data_in	: IN STD_LOGIC_VECTOR (21 DOWNTO 0);
			read_param	: IN STD_LOGIC ;
			read_source	: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
			busy	: OUT STD_LOGIC ;
			data_out	: OUT STD_LOGIC_VECTOR (28 DOWNTO 0);
			param	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			reconfig	: IN STD_LOGIC ;
			reset	: IN STD_LOGIC ;
			reset_timer	: IN STD_LOGIC ;
			write_param	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	busy    <= sub_wire0;
	data_out    <= sub_wire1(28 DOWNTO 0);

	remote_update_rmtupdt_51n_component : remote_update_rmtupdt_51n
	PORT MAP (
		clock => clock,
		data_in => data_in,
		read_param => read_param,
		read_source => read_source,
		param => param,
		reconfig => reconfig,
		reset => reset,
		reset_timer => reset_timer,
		write_param => write_param,
		busy => sub_wire0,
		data_out => sub_wire1
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: SIM_INIT_PAGE_SELECT_COMBO STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT0_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT1_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT2_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT3_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT4_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_WATCHDOG_VALUE_EDIT STRING "1"
-- Retrieval info: PRIVATE: SUPPORT_WRITE_CHECK STRING "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WATCHDOG_ENABLE_CHECK STRING "0"
-- Retrieval info: CONSTANT: CHECK_APP_POF STRING "false"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: IN_DATA_WIDTH NUMERIC "22"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "REMOTE"
-- Retrieval info: CONSTANT: OUT_DATA_WIDTH NUMERIC "29"
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: data_in 0 0 22 0 INPUT NODEFVAL "data_in[21..0]"
-- Retrieval info: USED_PORT: data_out 0 0 29 0 OUTPUT NODEFVAL "data_out[28..0]"
-- Retrieval info: USED_PORT: param 0 0 3 0 INPUT NODEFVAL "param[2..0]"
-- Retrieval info: USED_PORT: read_param 0 0 0 0 INPUT NODEFVAL "read_param"
-- Retrieval info: USED_PORT: read_source 0 0 2 0 INPUT NODEFVAL "read_source[1..0]"
-- Retrieval info: USED_PORT: reconfig 0 0 0 0 INPUT NODEFVAL "reconfig"
-- Retrieval info: USED_PORT: reset 0 0 0 0 INPUT NODEFVAL "reset"
-- Retrieval info: USED_PORT: reset_timer 0 0 0 0 INPUT NODEFVAL "reset_timer"
-- Retrieval info: USED_PORT: write_param 0 0 0 0 INPUT NODEFVAL "write_param"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @data_in 0 0 22 0 data_in 0 0 22 0
-- Retrieval info: CONNECT: @param 0 0 3 0 param 0 0 3 0
-- Retrieval info: CONNECT: @read_param 0 0 0 0 read_param 0 0 0 0
-- Retrieval info: CONNECT: @read_source 0 0 2 0 read_source 0 0 2 0
-- Retrieval info: CONNECT: @reconfig 0 0 0 0 reconfig 0 0 0 0
-- Retrieval info: CONNECT: @reset 0 0 0 0 reset 0 0 0 0
-- Retrieval info: CONNECT: @reset_timer 0 0 0 0 reset_timer 0 0 0 0
-- Retrieval info: CONNECT: @write_param 0 0 0 0 write_param 0 0 0 0
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: CONNECT: data_out 0 0 29 0 @data_out 0 0 29 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL remote_update.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL remote_update.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL remote_update.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL remote_update.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL remote_update_inst.vhd FALSE
-- Retrieval info: LIB_FILE: cycloneive
-- Retrieval info: LIB_FILE: lpm
