
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80de",
X"bc738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80e1",
X"dc0c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580d8",
X"e92d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580d6fd",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80d0b404",
X"f23d0d60",
X"913dec11",
X"56565990",
X"53f01552",
X"78519488",
X"3f83e080",
X"0880e538",
X"7a902e09",
X"810680dc",
X"3802b305",
X"3380e1e4",
X"0b80e1e4",
X"33575757",
X"8c397477",
X"2e8a3884",
X"16703356",
X"5674f338",
X"75337058",
X"5574802e",
X"80cf3880",
X"0b821722",
X"70832a57",
X"58587775",
X"27bb3896",
X"800a5790",
X"3dec0554",
X"80c08053",
X"76527851",
X"93aa3f83",
X"e0800888",
X"387a80c0",
X"802e8538",
X"80579a39",
X"811880c0",
X"80188218",
X"2270832a",
X"585c5858",
X"747826cb",
X"38811633",
X"577683e0",
X"800c903d",
X"0d04fc3d",
X"0d767052",
X"55b3c63f",
X"83e08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"811451b2",
X"de3f83e0",
X"80083070",
X"83e08008",
X"07802583",
X"e0800c53",
X"863d0d04",
X"fc3d0d76",
X"70525599",
X"ff3f83e0",
X"80085481",
X"5383e080",
X"0880c738",
X"745199c2",
X"3f83e080",
X"080b0b80",
X"e09c5383",
X"e0800852",
X"53ff8f3f",
X"83e08008",
X"a5380b0b",
X"80e0a052",
X"7251fefe",
X"3f83e080",
X"0894380b",
X"0b80e0a4",
X"527251fe",
X"ed3f83e0",
X"8008802e",
X"83388154",
X"73537283",
X"e0800c86",
X"3d0d04fd",
X"3d0d7570",
X"52549998",
X"3f815383",
X"e0800898",
X"38735198",
X"e13f83e0",
X"a0085283",
X"e0800851",
X"feb43f83",
X"e0800853",
X"7283e080",
X"0c853d0d",
X"04e03d0d",
X"a33d0870",
X"525e8f87",
X"3f83e080",
X"0833943d",
X"56547394",
X"3880e49c",
X"52745184",
X"c6397d52",
X"7851928a",
X"3f84d039",
X"7d518eef",
X"3f83e080",
X"08527451",
X"8e9f3f83",
X"e0a80852",
X"933d7052",
X"5d94fa3f",
X"83e08008",
X"59800b83",
X"e0800855",
X"5b83e080",
X"087b2e94",
X"38811b74",
X"525b97fb",
X"3f83e080",
X"085483e0",
X"8008ee38",
X"805aff7a",
X"437a427a",
X"415f7909",
X"709f2c7b",
X"065b547a",
X"7a248438",
X"ff1b5af6",
X"1a700970",
X"9f2c7206",
X"7bff125a",
X"5a525555",
X"80752595",
X"38765197",
X"ba3f83e0",
X"800876ff",
X"18585557",
X"738024ed",
X"38747f2e",
X"8638b998",
X"3f745f78",
X"ff1b7058",
X"5d58807a",
X"25953877",
X"5197903f",
X"83e08008",
X"76ff1858",
X"55587380",
X"24ed3880",
X"0b83e3a8",
X"0c800b83",
X"e3c80c0b",
X"0b80e0a8",
X"518be33f",
X"81800b83",
X"e3c80c0b",
X"0b80e0b0",
X"518bd33f",
X"a80b83e3",
X"a80c7680",
X"2e80e838",
X"83e3a808",
X"77793270",
X"30707207",
X"80257087",
X"2b83e3c8",
X"0c515678",
X"53565696",
X"c33f83e0",
X"8008802e",
X"8a380b0b",
X"80e0b851",
X"8b983f76",
X"5196833f",
X"83e08008",
X"520b0b80",
X"e0ec518b",
X"853f7651",
X"96893f83",
X"e0800883",
X"e3a80855",
X"57757425",
X"8638a816",
X"56f73975",
X"83e3a80c",
X"86f07624",
X"ff943887",
X"980b83e3",
X"a80c7780",
X"2eb73877",
X"5195bf3f",
X"83e08008",
X"78525595",
X"df3f0b0b",
X"80e0c054",
X"83e08008",
X"8f388739",
X"807634fd",
X"96390b0b",
X"80e0bc54",
X"74537352",
X"0b0b80e0",
X"8c518a9e",
X"3f80540b",
X"0b80e094",
X"518a933f",
X"81145473",
X"a82e0981",
X"06ed3886",
X"8da051b5",
X"983f8052",
X"903d7052",
X"5480c3a3",
X"3f835273",
X"5180c39b",
X"3f61802e",
X"80ff387b",
X"5473ff2e",
X"96387880",
X"2e818038",
X"785194df",
X"3f83e080",
X"08ff1555",
X"59e73978",
X"802e80eb",
X"38785194",
X"db3f83e0",
X"8008802e",
X"fc843878",
X"5194a33f",
X"83e08008",
X"520b0b80",
X"e09851ac",
X"813f83e0",
X"8008a438",
X"7c51adb9",
X"3f83e080",
X"085574ff",
X"16565480",
X"7425fbef",
X"38741d70",
X"33555673",
X"af2efec8",
X"38e83978",
X"5193e13f",
X"83e08008",
X"527c51ac",
X"f03ffbcf",
X"397f8829",
X"6010057a",
X"0561055a",
X"fc8039a2",
X"3d0d04fe",
X"3d0d80e3",
X"a4087033",
X"7081ff06",
X"70842a81",
X"32810655",
X"51525371",
X"802e8c38",
X"a8733480",
X"e3a40851",
X"b8713471",
X"83e0800c",
X"843d0d04",
X"fe3d0d80",
X"e3a40870",
X"337081ff",
X"0670852a",
X"81328106",
X"55515253",
X"71802e8c",
X"38987334",
X"80e3a408",
X"51b87134",
X"7183e080",
X"0c843d0d",
X"04803d0d",
X"80e3a008",
X"51937134",
X"80e3ac08",
X"51ff7134",
X"823d0d04",
X"fe3d0d02",
X"93053380",
X"e3a00853",
X"53807234",
X"8a51b2e1",
X"3fd33f80",
X"e3b00852",
X"80f87234",
X"80e3c808",
X"52807234",
X"fa1380e3",
X"d0085353",
X"72723480",
X"e3b80852",
X"80723480",
X"e3c00852",
X"72723480",
X"e3a40852",
X"80723480",
X"e3a40852",
X"b8723484",
X"3d0d04ff",
X"3d0d028f",
X"053380e3",
X"a8085252",
X"717134fe",
X"9e3f83e0",
X"8008802e",
X"f638833d",
X"0d04803d",
X"0d8439bb",
X"bf3ffeb8",
X"3f83e080",
X"08802ef3",
X"3880e3a8",
X"08703370",
X"81ff0683",
X"e0800c51",
X"51823d0d",
X"04803d0d",
X"80e3a008",
X"51a37134",
X"80e3ac08",
X"51ff7134",
X"80e3a408",
X"51a87134",
X"80e3a408",
X"51b87134",
X"823d0d04",
X"803d0d80",
X"e3a00870",
X"337081c0",
X"06703070",
X"802583e0",
X"800c5151",
X"5151823d",
X"0d04ff3d",
X"0d80e3a4",
X"08703370",
X"81ff0670",
X"832a8132",
X"70810651",
X"51515252",
X"70802ee5",
X"38b07234",
X"80e3a408",
X"51b87134",
X"833d0d04",
X"803d0d80",
X"e3dc0870",
X"08810683",
X"e0800c51",
X"823d0d04",
X"fd3d0d75",
X"77545480",
X"73259438",
X"73708105",
X"55335280",
X"e0c45185",
X"a13fff13",
X"53e93985",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"80c1883f",
X"83e08008",
X"7a27ed38",
X"74802e80",
X"e0387452",
X"755180c0",
X"f23f83e0",
X"80087553",
X"76525480",
X"c1983f83",
X"e080087a",
X"53755256",
X"80c0d83f",
X"83e08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"e08008c2",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9c",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fbfd3f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd13f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbad3f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83e0900c",
X"7183e094",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383e090",
X"085283e0",
X"940851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"9aaa5351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fd3d",
X"0d757052",
X"54a3c23f",
X"83e08008",
X"14537274",
X"2e9238ff",
X"13703353",
X"5371af2e",
X"098106ee",
X"38811353",
X"7283e080",
X"0c853d0d",
X"04fd3d0d",
X"75777053",
X"5454c73f",
X"83e08008",
X"732ea138",
X"83e08008",
X"733152ff",
X"125271ff",
X"2e8f3872",
X"70810554",
X"33747081",
X"055634eb",
X"39ff1454",
X"80743485",
X"3d0d0480",
X"3d0d7251",
X"ff903f82",
X"3d0d0471",
X"83e0800c",
X"04803d0d",
X"72518071",
X"34810bbc",
X"120c800b",
X"80c0120c",
X"823d0d04",
X"800b83e2",
X"d408248a",
X"38b9f13f",
X"ff0b83e2",
X"d40c800b",
X"83e0800c",
X"04ff3d0d",
X"735283e0",
X"b008722e",
X"8d38d93f",
X"71519697",
X"3f7183e0",
X"b00c833d",
X"0d04f43d",
X"0d7e6062",
X"5c5a5581",
X"54bc1508",
X"81913874",
X"51cf3f79",
X"58807a25",
X"80f73883",
X"e3840870",
X"892a5783",
X"ff067884",
X"80723156",
X"56577378",
X"25833873",
X"557583e2",
X"d4082e84",
X"38ff893f",
X"83e2d408",
X"8025a638",
X"75892b51",
X"98da3f83",
X"e384088f",
X"3dfc1155",
X"5c548152",
X"f81b5196",
X"c43f7614",
X"83e3840c",
X"7583e2d4",
X"0c745376",
X"527851b8",
X"843f83e0",
X"800883e3",
X"84081683",
X"e3840c78",
X"7631761b",
X"5b595677",
X"8024ff8b",
X"38617a71",
X"0c547554",
X"75802e83",
X"38815473",
X"83e0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"9b3f7651",
X"feaf3f86",
X"3dfc0553",
X"78527751",
X"95e73f79",
X"75710c54",
X"83e08008",
X"5483e080",
X"08802e83",
X"38815473",
X"83e0800c",
X"863d0d04",
X"fe3d0d75",
X"83e2d408",
X"53538072",
X"24893871",
X"732e8438",
X"fdd63f74",
X"51fdea3f",
X"725197ac",
X"3f83e080",
X"085283e0",
X"8008802e",
X"83388152",
X"7183e080",
X"0c843d0d",
X"04803d0d",
X"7280c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d72bc11",
X"0883e080",
X"0c51823d",
X"0d0480c4",
X"0b83e080",
X"0c04fd3d",
X"0d757771",
X"54705355",
X"539f9a3f",
X"82c81308",
X"bc150c82",
X"c0130880",
X"c0150cfc",
X"eb3f7351",
X"93a93f73",
X"83e0b00c",
X"83e08008",
X"5383e080",
X"08802e83",
X"38815372",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"775553fc",
X"bf3f7280",
X"2ea538bc",
X"13085273",
X"519ea43f",
X"83e08008",
X"8f387752",
X"7251ff9a",
X"3f83e080",
X"08538a39",
X"82cc1308",
X"53d83981",
X"537283e0",
X"800c853d",
X"0d04fe3d",
X"0dff0b83",
X"e2d40c74",
X"83e0b40c",
X"7583e2d0",
X"0cb4c83f",
X"83e08008",
X"81ff0652",
X"81537199",
X"3883e2ec",
X"518e933f",
X"83e08008",
X"5283e080",
X"08802e83",
X"38725271",
X"537283e0",
X"800c843d",
X"0d04fa3d",
X"0d787a82",
X"c4120882",
X"c4120870",
X"72245956",
X"56575773",
X"732e0981",
X"06913880",
X"c0165280",
X"c017519c",
X"953f83e0",
X"80085574",
X"83e0800c",
X"883d0d04",
X"f63d0d7c",
X"5b807b71",
X"5c54577a",
X"772e8c38",
X"811a82cc",
X"1408545a",
X"72f63880",
X"5980d939",
X"7a548157",
X"80707b7b",
X"315a5755",
X"ff185374",
X"732580c1",
X"3882cc14",
X"08527351",
X"ff8c3f80",
X"0b83e080",
X"0825a138",
X"82cc1408",
X"82cc1108",
X"82cc160c",
X"7482cc12",
X"0c537580",
X"2e863872",
X"82cc170c",
X"72548057",
X"7382cc15",
X"08811757",
X"5556ffb8",
X"39811959",
X"800bff1b",
X"54547873",
X"25833881",
X"54768132",
X"70750651",
X"5372ff90",
X"388c3d0d",
X"04f73d0d",
X"7b7d5a5a",
X"82d05283",
X"e2d00851",
X"b4913f83",
X"e0800857",
X"f9e23f79",
X"5283e2d8",
X"5195b43f",
X"83e08008",
X"54805383",
X"e0800873",
X"2e098106",
X"82833883",
X"e0b4080b",
X"0b80e098",
X"53705256",
X"9bd33f0b",
X"0b80e098",
X"5280c016",
X"519bc63f",
X"75bc170c",
X"7382c017",
X"0c810b82",
X"c4170c81",
X"0b82c817",
X"0c7382cc",
X"170cff17",
X"82d01755",
X"57819139",
X"83e0c033",
X"70822a70",
X"81065154",
X"55728180",
X"3874812a",
X"81065877",
X"80f63874",
X"842a8106",
X"82c4150c",
X"83e0c033",
X"810682c8",
X"150c7952",
X"73519aed",
X"3f73519b",
X"843f83e0",
X"80081453",
X"af737081",
X"05553472",
X"bc150c83",
X"e0c15272",
X"519ace3f",
X"83e0b808",
X"82c0150c",
X"83e0ce52",
X"80c01451",
X"9abb3f78",
X"802e8d38",
X"7351782d",
X"83e08008",
X"802e9938",
X"7782cc15",
X"0c75802e",
X"86387382",
X"cc170c73",
X"82d015ff",
X"19595556",
X"76802e9b",
X"3883e0b8",
X"5283e2d8",
X"5194aa3f",
X"83e08008",
X"8a3883e0",
X"c1335372",
X"fed23878",
X"802e8938",
X"83e0b408",
X"51fcb93f",
X"83e0b408",
X"537283e0",
X"800c8b3d",
X"0d04ff3d",
X"0d805273",
X"51fdb63f",
X"833d0d04",
X"f03d0d62",
X"705254f6",
X"913f83e0",
X"80087453",
X"873d7053",
X"5555f6b1",
X"3ff7913f",
X"7351d33f",
X"63537452",
X"83e08008",
X"51fab93f",
X"923d0d04",
X"7183e080",
X"0c0480c0",
X"1283e080",
X"0c04803d",
X"0d7282c0",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"cc110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"82c41108",
X"83e0800c",
X"51823d0d",
X"04f93d0d",
X"7983e098",
X"08575781",
X"77278196",
X"38768817",
X"0827818e",
X"38753355",
X"74822e89",
X"3874832e",
X"b33880fe",
X"39745476",
X"1083fe06",
X"5376882a",
X"8c170805",
X"52893dfc",
X"0551aee4",
X"3f83e080",
X"0880df38",
X"029d0533",
X"893d3371",
X"882b0756",
X"5680d139",
X"84547682",
X"2b83fc06",
X"5376872a",
X"8c170805",
X"52893dfc",
X"0551aeb4",
X"3f83e080",
X"08b03802",
X"9f053302",
X"84059e05",
X"3371982b",
X"71902b07",
X"028c059d",
X"05337088",
X"2b72078d",
X"3d337180",
X"fffffe80",
X"06075152",
X"53575856",
X"83398155",
X"7483e080",
X"0c893d0d",
X"04fb3d0d",
X"83e09808",
X"fe198812",
X"08fe0555",
X"56548056",
X"7473278d",
X"38821433",
X"75712994",
X"16080557",
X"537583e0",
X"800c873d",
X"0d04fc3d",
X"0d765280",
X"0b83e098",
X"08703351",
X"52537083",
X"2e098106",
X"91389512",
X"33941333",
X"71982b71",
X"902b0755",
X"55519b12",
X"339a1333",
X"71882b07",
X"740783e0",
X"800c5586",
X"3d0d04fc",
X"3d0d7683",
X"e0980855",
X"55807523",
X"88150853",
X"72812e88",
X"38881408",
X"73268538",
X"8152b239",
X"72903873",
X"33527183",
X"2e098106",
X"85389014",
X"0853728c",
X"160c7280",
X"2e8d3872",
X"51fed63f",
X"83e08008",
X"52853990",
X"14085271",
X"90160c80",
X"527183e0",
X"800c863d",
X"0d04fa3d",
X"0d7883e0",
X"98087122",
X"81057083",
X"ffff0657",
X"54575573",
X"802e8838",
X"90150853",
X"72863883",
X"5280e739",
X"738f0652",
X"7180da38",
X"81139016",
X"0c8c1508",
X"53729038",
X"830b8417",
X"22575273",
X"762780c6",
X"38bf3982",
X"1633ff05",
X"74842a06",
X"5271b238",
X"7251fcb1",
X"3f815271",
X"83e08008",
X"27a83883",
X"5283e080",
X"08881708",
X"279c3883",
X"e080088c",
X"160c83e0",
X"800851fd",
X"bc3f83e0",
X"80089016",
X"0c737523",
X"80527183",
X"e0800c88",
X"3d0d04f2",
X"3d0d6062",
X"64585e5b",
X"75335574",
X"a02e0981",
X"06883881",
X"16704456",
X"ef396270",
X"33565674",
X"af2e0981",
X"06843881",
X"1643800b",
X"881c0c62",
X"70335155",
X"749f2691",
X"387a51fd",
X"d23f83e0",
X"80085680",
X"7d348381",
X"39933d84",
X"1c087058",
X"595f8a55",
X"a0767081",
X"055834ff",
X"155574ff",
X"2e098106",
X"ef388070",
X"5a5c887f",
X"085f5a7b",
X"811d7081",
X"ff066013",
X"703370af",
X"327030a0",
X"73277180",
X"25075151",
X"525b535e",
X"57557480",
X"e73876ae",
X"2e098106",
X"83388155",
X"787a2775",
X"07557480",
X"2e9f3879",
X"88327030",
X"78ae3270",
X"30707307",
X"9f2a5351",
X"57515675",
X"bb388859",
X"8b5affab",
X"3976982b",
X"55748025",
X"873880dd",
X"cc173357",
X"ff9f1755",
X"74992689",
X"38e01770",
X"81ff0658",
X"5578811a",
X"7081ff06",
X"721b535b",
X"57557675",
X"34fef839",
X"7b1e7f0c",
X"805576a0",
X"26833881",
X"55748b19",
X"347a51fc",
X"823f83e0",
X"800880f5",
X"38a0547a",
X"2270852b",
X"83e00654",
X"55901b08",
X"527c51a8",
X"ef3f83e0",
X"80085783",
X"e0800881",
X"81387c33",
X"5574802e",
X"80f4388b",
X"1d337083",
X"2a708106",
X"51565674",
X"b4388b7d",
X"841d0883",
X"e0800859",
X"5b5b58ff",
X"185877ff",
X"2e9a3879",
X"7081055b",
X"33797081",
X"055b3371",
X"71315256",
X"5675802e",
X"e2388639",
X"75802e96",
X"387a51fb",
X"e53fff86",
X"3983e080",
X"085683e0",
X"8008b638",
X"83397656",
X"841b088b",
X"11335155",
X"74a7388b",
X"1d337084",
X"2a708106",
X"51565674",
X"89388356",
X"94398156",
X"90397c51",
X"fa943f83",
X"e0800888",
X"1c0cfd81",
X"397583e0",
X"800c903d",
X"0d04f83d",
X"0d7a7c59",
X"57825483",
X"fe537752",
X"7651a7b4",
X"3f835683",
X"e0800880",
X"ec388117",
X"33773371",
X"882b0756",
X"56825674",
X"82d4d52e",
X"09810680",
X"d4387554",
X"b6537752",
X"7651a788",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"ac388254",
X"80d25377",
X"527651a6",
X"df3f83e0",
X"80089838",
X"81173377",
X"3371882b",
X"0783e080",
X"08525656",
X"748182c6",
X"2e833881",
X"567583e0",
X"800c8a3d",
X"0d04eb3d",
X"0d675a80",
X"0b83e098",
X"0ca6943f",
X"83e08008",
X"81065582",
X"567483ee",
X"38747553",
X"8f3d7053",
X"5759feca",
X"3f83e080",
X"0881ff06",
X"5776812e",
X"09810680",
X"d4389054",
X"83be5374",
X"527551a5",
X"f33f83e0",
X"800880c9",
X"388f3d33",
X"5574802e",
X"80c93802",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"70587b57",
X"5e525e57",
X"5957fdee",
X"3f83e080",
X"0881ff06",
X"5776832e",
X"09810686",
X"38815682",
X"f1397680",
X"2e863886",
X"5682e739",
X"a4548d53",
X"78527551",
X"a58a3f81",
X"5683e080",
X"0882d338",
X"02be0533",
X"028405bd",
X"05337188",
X"2b07595d",
X"77ab3802",
X"80ce0533",
X"02840580",
X"cd053371",
X"982b7190",
X"2b07973d",
X"3370882b",
X"72070294",
X"0580cb05",
X"33710754",
X"525e5759",
X"5602b705",
X"33787129",
X"028805b6",
X"0533028c",
X"05b50533",
X"71882b07",
X"701d707f",
X"8c050c5f",
X"5957595d",
X"8e3d3382",
X"1b3402b9",
X"0533903d",
X"3371882b",
X"075a5c78",
X"841b2302",
X"bb053302",
X"8405ba05",
X"3371882b",
X"07565c74",
X"ab380280",
X"ca053302",
X"840580c9",
X"05337198",
X"2b71902b",
X"07963d33",
X"70882b72",
X"07029405",
X"80c70533",
X"71075152",
X"53575e5c",
X"74763178",
X"3179842a",
X"903d3354",
X"71713153",
X"5656a4f7",
X"3f83e080",
X"08820570",
X"881c0c83",
X"e08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83e0980c",
X"80567583",
X"e0800c97",
X"3d0d04e9",
X"3d0d83e0",
X"98085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e63f83e0",
X"80085483",
X"e0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f48a",
X"3f83e080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383e080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83e09808",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0ea3f",
X"83e08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"843f83e0",
X"80085583",
X"e0800880",
X"2eff8938",
X"83e08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"519fb13f",
X"83e08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83e0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83e09808",
X"55568555",
X"73802e81",
X"e1388114",
X"33810653",
X"84557280",
X"2e81d338",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b7388214",
X"3370892b",
X"56537680",
X"2eb53874",
X"52ff1651",
X"9ff93f83",
X"e08008ff",
X"18765470",
X"5358539f",
X"ea3f83e0",
X"80087326",
X"96387430",
X"70780670",
X"98170c77",
X"7131a417",
X"08525851",
X"538939a0",
X"140870a4",
X"160c5374",
X"7627b938",
X"7251eed9",
X"3f83e080",
X"0853810b",
X"83e08008",
X"278b3888",
X"140883e0",
X"80082688",
X"38800b81",
X"1534b039",
X"83e08008",
X"a4150c98",
X"14081598",
X"150c7575",
X"3156c439",
X"98140816",
X"7098160c",
X"735256ef",
X"c83f83e0",
X"80088c38",
X"83e08008",
X"81153481",
X"55943982",
X"1433ff05",
X"76892a06",
X"83e08008",
X"05a8150c",
X"80557483",
X"e0800c88",
X"3d0d04ef",
X"3d0d6356",
X"855583e0",
X"9808802e",
X"80d23893",
X"3df40584",
X"170c6453",
X"883d7053",
X"765257f1",
X"d23f83e0",
X"80085583",
X"e08008b4",
X"38883d33",
X"5473802e",
X"a13802a7",
X"05337084",
X"2a708106",
X"51555583",
X"5573802e",
X"97387651",
X"eef83f83",
X"e0800888",
X"170c7551",
X"efa93f83",
X"e0800855",
X"7483e080",
X"0c933d0d",
X"04e43d0d",
X"6ea13d08",
X"405e8556",
X"83e09808",
X"802e8485",
X"389e3df4",
X"05841f0c",
X"7e98387d",
X"51eef83f",
X"83e08008",
X"5683ee39",
X"814181f6",
X"39834181",
X"f139933d",
X"7f960541",
X"59807f82",
X"95055e56",
X"756081ff",
X"05348341",
X"901e0876",
X"2e81d338",
X"a0547d22",
X"70852b83",
X"e0065458",
X"901e0852",
X"78519bbc",
X"3f83e080",
X"084183e0",
X"8008ffb8",
X"3878335c",
X"7b802eff",
X"b4388b19",
X"3370bf06",
X"71810652",
X"43557480",
X"2e80de38",
X"7b81bf06",
X"55748f24",
X"80d3389a",
X"19335574",
X"80cb38f3",
X"1d70585d",
X"8156758b",
X"2e098106",
X"85388e56",
X"8b39759a",
X"2e098106",
X"83389c56",
X"75197070",
X"81055233",
X"7133811a",
X"821a5f5b",
X"525b5574",
X"86387977",
X"34853980",
X"df773477",
X"7b57577a",
X"a02e0981",
X"06c03881",
X"567b81e5",
X"32703070",
X"9f2a5151",
X"557bae2e",
X"93387480",
X"2e8e3861",
X"832a7081",
X"06515574",
X"802e9738",
X"7d51ede2",
X"3f83e080",
X"084183e0",
X"80088738",
X"901e08fe",
X"af388060",
X"3475802e",
X"88387c52",
X"7f5183a5",
X"3f60802e",
X"8638800b",
X"901f0c60",
X"5660832e",
X"85386081",
X"d038891f",
X"57901e08",
X"802e81a8",
X"38805675",
X"19703351",
X"5574a02e",
X"a0387485",
X"2e098106",
X"843881e5",
X"55747770",
X"81055934",
X"81167081",
X"ff065755",
X"877627d7",
X"38881933",
X"5574a02e",
X"a938ae77",
X"70810559",
X"34885675",
X"19703351",
X"5574a02e",
X"95387477",
X"70810559",
X"34811670",
X"81ff0657",
X"558a7627",
X"e2388b19",
X"337f8805",
X"349f1933",
X"9e1a3371",
X"982b7190",
X"2b079d1c",
X"3370882b",
X"72079c1e",
X"33710764",
X"0c52991d",
X"33981e33",
X"71882b07",
X"53515357",
X"5956747f",
X"84052397",
X"1933961a",
X"3371882b",
X"07565674",
X"7f860523",
X"8077347d",
X"51ebf33f",
X"83e08008",
X"83327030",
X"7072079f",
X"2c83e080",
X"08065256",
X"56961f33",
X"55748a38",
X"891f5296",
X"1f5181b1",
X"3f7583e0",
X"800c9e3d",
X"0d04fd3d",
X"0d757753",
X"54733351",
X"70893871",
X"33517080",
X"2ea13873",
X"33723352",
X"53727127",
X"8538ff51",
X"94397073",
X"27853881",
X"518b3981",
X"14811353",
X"54d33980",
X"517083e0",
X"800c853d",
X"0d04fd3d",
X"0d757754",
X"54723370",
X"81ff0652",
X"5270802e",
X"a3387181",
X"ff068114",
X"ffbf1253",
X"54527099",
X"268938a0",
X"127081ff",
X"06535171",
X"74708105",
X"5634d239",
X"80743485",
X"3d0d04ff",
X"bd3d0d80",
X"c63d0852",
X"a53d7052",
X"54ffb33f",
X"80c73d08",
X"52853d70",
X"5253ffa6",
X"3f725273",
X"51fedf3f",
X"80c53d0d",
X"04fe3d0d",
X"74765353",
X"71708105",
X"53335170",
X"73708105",
X"553470f0",
X"38843d0d",
X"04fe3d0d",
X"74528072",
X"33525370",
X"732e8d38",
X"81128114",
X"71335354",
X"5270f538",
X"7283e080",
X"0c843d0d",
X"047183e3",
X"9c0c8880",
X"800b83e3",
X"980c8480",
X"800b83e3",
X"a00c04f0",
X"3d0d8380",
X"805683e3",
X"9c081683",
X"e3980817",
X"56547433",
X"743483e3",
X"a0081654",
X"80743481",
X"16567583",
X"80a02e09",
X"8106db38",
X"83d08056",
X"83e39c08",
X"1683e398",
X"08175654",
X"74337434",
X"83e3a008",
X"16548074",
X"34811656",
X"7583d0a0",
X"2e098106",
X"db3883a8",
X"805683e3",
X"9c081683",
X"e3980817",
X"56547433",
X"743483e3",
X"a0081654",
X"80743481",
X"16567583",
X"a8902e09",
X"8106db38",
X"805683e3",
X"9c081683",
X"e3a00817",
X"55557333",
X"75348116",
X"56758180",
X"802e0981",
X"06e43887",
X"833f893d",
X"58a25380",
X"dfcc5277",
X"519d8b3f",
X"80578c80",
X"5683e3a0",
X"08167719",
X"55557333",
X"75348116",
X"81185856",
X"76a22e09",
X"8106e638",
X"80e2e808",
X"54867434",
X"80e2ec08",
X"54807434",
X"80e39c08",
X"54807434",
X"80e38c08",
X"54af7434",
X"80e39808",
X"54bf7434",
X"80e39408",
X"54807434",
X"80e39008",
X"549f7434",
X"80e38808",
X"54807434",
X"80e2f808",
X"54f87434",
X"80e2f008",
X"54767434",
X"80e2e008",
X"54827434",
X"80e2f408",
X"54827434",
X"923d0d04",
X"fe3d0d80",
X"5383e3a0",
X"081383e3",
X"9c081452",
X"52703372",
X"34811353",
X"72818080",
X"2e098106",
X"e4388380",
X"805383e3",
X"a0081383",
X"e39c0814",
X"52527033",
X"72348113",
X"53728380",
X"a02e0981",
X"06e43883",
X"d0805383",
X"e3a00813",
X"83e39c08",
X"14525270",
X"33723481",
X"13537283",
X"d0a02e09",
X"8106e438",
X"83a88053",
X"83e3a008",
X"1383e39c",
X"08145252",
X"70337234",
X"81135372",
X"83a8902e",
X"098106e4",
X"38843d0d",
X"04803d0d",
X"80e3f808",
X"70088106",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"80e3f808",
X"700870fe",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d80e3",
X"f8087008",
X"70812c81",
X"0683e080",
X"0c515182",
X"3d0d04ff",
X"3d0d80e3",
X"f8087008",
X"70fd0676",
X"1007720c",
X"5252833d",
X"0d04803d",
X"0d80e3f8",
X"08700870",
X"822cbf06",
X"83e0800c",
X"5151823d",
X"0d04ff3d",
X"0d80e3f8",
X"08700870",
X"fe830676",
X"822b0772",
X"0c525283",
X"3d0d0480",
X"3d0d80e3",
X"f8087008",
X"70882c87",
X"0683e080",
X"0c515182",
X"3d0d04ff",
X"3d0d80e3",
X"f8087008",
X"70f1ff06",
X"76882b07",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"e3f80870",
X"08708b2c",
X"bf0683e0",
X"800c5151",
X"823d0d04",
X"ff3d0d80",
X"e3f80870",
X"0870f88f",
X"ff06768b",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d80e3f8",
X"08700870",
X"912cbf06",
X"83e0800c",
X"5151823d",
X"0d04ff3d",
X"0d80e3f8",
X"08700870",
X"fc87ffff",
X"0676912b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80e48808",
X"70087088",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04803d0d",
X"80e48808",
X"70087089",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04803d0d",
X"80e48808",
X"7008708a",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04803d0d",
X"80e48808",
X"7008708b",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04fd3d0d",
X"7581e629",
X"872a80e3",
X"e8085473",
X"0c853d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727081",
X"055434ff",
X"1151f039",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708405",
X"540cff11",
X"51f03984",
X"3d0d04fe",
X"3d0d8180",
X"80538052",
X"88800a51",
X"ffb33fa0",
X"80538052",
X"82800a51",
X"c73f843d",
X"0d04803d",
X"0d8151fc",
X"9c3f7280",
X"2e8338d3",
X"3f8151fc",
X"be3f8051",
X"fcb93f80",
X"51fc863f",
X"823d0d04",
X"fd3d0d75",
X"52805480",
X"ff722588",
X"38810bff",
X"80135354",
X"ffbf1251",
X"70992686",
X"38e01252",
X"9e39ff9f",
X"12519971",
X"279538d0",
X"12e01370",
X"54545189",
X"71278838",
X"8f732783",
X"38805273",
X"802e8538",
X"81801252",
X"7181ff06",
X"83e0800c",
X"853d0d04",
X"803d0d84",
X"d8c05180",
X"71708105",
X"53347084",
X"e0c02e09",
X"8106f038",
X"823d0d04",
X"fe3d0d02",
X"97053351",
X"ff863f83",
X"e0800881",
X"ff0683e3",
X"a8085452",
X"8073249b",
X"3883e3c4",
X"08137283",
X"e3c80807",
X"53537173",
X"3483e3a8",
X"08810583",
X"e3a80c84",
X"3d0d04fa",
X"3d0d8280",
X"0a1b5580",
X"57883dfc",
X"05547953",
X"74527851",
X"d5da3f88",
X"3d0d04fe",
X"3d0d83e3",
X"c0085274",
X"51dcbd3f",
X"83e08008",
X"8c387653",
X"755283e3",
X"c00851c7",
X"3f843d0d",
X"04fe3d0d",
X"83e3c008",
X"53755274",
X"51d6fd3f",
X"83e08008",
X"8d387753",
X"765283e3",
X"c00851ff",
X"a23f843d",
X"0d04fd3d",
X"0d83e3c0",
X"0851d5f1",
X"3f83e080",
X"0890802e",
X"098106ad",
X"38805483",
X"c1808053",
X"83e08008",
X"5283e3c0",
X"0851fef3",
X"3f87c180",
X"80143387",
X"c1908015",
X"34811454",
X"7390802e",
X"098106e9",
X"38853d0d",
X"0480e0cc",
X"0b83e080",
X"0c04f73d",
X"0d805a80",
X"59805880",
X"705757fd",
X"e73f800b",
X"83e3a80c",
X"800b83e3",
X"c80c80e0",
X"d051d0d6",
X"3f81800b",
X"83e3c80c",
X"80e0d451",
X"d0c83f80",
X"d00b83e3",
X"a80c7530",
X"70770780",
X"2570872b",
X"83e3c80c",
X"5154f99e",
X"3f83e080",
X"085280e0",
X"dc51d0a2",
X"3f80f80b",
X"83e3a80c",
X"75813270",
X"30707207",
X"80257087",
X"2b83e3c8",
X"0c515555",
X"ff833f83",
X"e0800852",
X"80e0e851",
X"cff83f81",
X"a00b83e3",
X"a80c7582",
X"32703070",
X"72078025",
X"70872b83",
X"e3c80c51",
X"5583e3c0",
X"085255d1",
X"923f83e0",
X"80085280",
X"e0f051cf",
X"c93f81c8",
X"0b83e3a8",
X"0c758332",
X"70307072",
X"07802570",
X"872b83e3",
X"c80c5155",
X"80e0f852",
X"55cfa73f",
X"81f00b83",
X"e3a80c75",
X"84327030",
X"70720780",
X"2570872b",
X"83e3c80c",
X"515580e1",
X"885255cf",
X"853f8298",
X"0b83e3a8",
X"0c758532",
X"70307072",
X"07802570",
X"872b83e3",
X"c80c5155",
X"80e1a052",
X"55cee33f",
X"82c00b83",
X"e3a80c75",
X"86327030",
X"70720780",
X"2570872b",
X"83e3c80c",
X"515580e1",
X"b85255ce",
X"c13f868d",
X"a051f9d1",
X"3f805288",
X"3d705254",
X"87dd3f83",
X"52735187",
X"d63f7816",
X"56758025",
X"85388056",
X"90398676",
X"25853886",
X"56873975",
X"862682db",
X"38758429",
X"80dff005",
X"54730804",
X"f6f03f83",
X"e0800878",
X"56547481",
X"2e098106",
X"893883e0",
X"80081054",
X"903974ff",
X"2e098106",
X"883883e0",
X"8008812c",
X"54907425",
X"85389054",
X"88397380",
X"24833881",
X"547351f6",
X"cd3f828f",
X"39f6e03f",
X"83e08008",
X"18547380",
X"25853880",
X"54883987",
X"74258338",
X"87547351",
X"f6dd3f81",
X"ee397787",
X"3879802e",
X"81e53883",
X"e0a40883",
X"e0a00c8c",
X"830b83e0",
X"a80c83e3",
X"c00851ff",
X"bfab3ffb",
X"b53f81c7",
X"3979802e",
X"81c13883",
X"e09c0883",
X"e0a00c8c",
X"830b83e0",
X"a80c83e3",
X"bc0851ff",
X"bf873f75",
X"832e0981",
X"06943881",
X"80805382",
X"80805283",
X"e3bc0851",
X"fa993f81",
X"87397584",
X"2e098106",
X"af388280",
X"80538180",
X"805283e3",
X"bc0851f9",
X"fe3f8054",
X"84828080",
X"14338481",
X"80801534",
X"81145473",
X"8180802e",
X"098106e8",
X"3880d139",
X"75852e09",
X"810680c8",
X"38805481",
X"80805380",
X"c0805283",
X"e3bc0851",
X"f9c53f82",
X"80805380",
X"c0805283",
X"e3bc0851",
X"f9b53f84",
X"81808014",
X"338481c0",
X"80153484",
X"82808014",
X"338482c0",
X"80153481",
X"14547380",
X"c0802e09",
X"8106dc38",
X"81548c39",
X"79873876",
X"802efac3",
X"38805473",
X"83e0800c",
X"8b3d0d04",
X"ff3d0df5",
X"d43f83e0",
X"8008802e",
X"86388051",
X"80dd39f5",
X"dc3f83e0",
X"800880d1",
X"38f6823f",
X"83e08008",
X"802eaa38",
X"8151f3a1",
X"3fefcc3f",
X"800b83e3",
X"a80cf9f2",
X"3f83e080",
X"0852ff0b",
X"83e3a80c",
X"f1ea3f71",
X"a4387151",
X"f2ff3fa2",
X"39f5b63f",
X"83e08008",
X"802e9738",
X"8151f2ed",
X"3fef983f",
X"ff0b83e3",
X"a80cf1c4",
X"3f8151f6",
X"b93f833d",
X"0d04fc3d",
X"0d908080",
X"52868480",
X"8051cffa",
X"3f83e080",
X"08b83880",
X"e48c51d4",
X"bd3f83e0",
X"800883e3",
X"c0085480",
X"e1c45383",
X"e0800852",
X"55cf993f",
X"83e08008",
X"8438f8aa",
X"3f818080",
X"54828080",
X"5380e1c0",
X"527451f7",
X"f43f8151",
X"f5e43ffe",
X"b73ffc39",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"0280e1d0",
X"0b83e0a4",
X"0c80e1d4",
X"0b83e09c",
X"0c80e1d8",
X"0b83e0ac",
X"0c83e08c",
X"08fc050c",
X"800b83e3",
X"ac0b83e0",
X"8c08f805",
X"0c83e08c",
X"08f4050c",
X"cde83f83",
X"e0800886",
X"05fc0683",
X"e08c08f0",
X"050c0283",
X"e08c08f0",
X"0508310d",
X"833d7083",
X"e08c08f8",
X"05087084",
X"0583e08c",
X"08f8050c",
X"0c51cab1",
X"3f83e08c",
X"08f40508",
X"810583e0",
X"8c08f405",
X"0c83e08c",
X"08f40508",
X"862e0981",
X"06ffad38",
X"86948080",
X"51ecfe3f",
X"ff0b83e3",
X"a80c800b",
X"83e3c80c",
X"84d8c00b",
X"83e3c40c",
X"8151f0cd",
X"3f8151f0",
X"f63f8051",
X"f0f13f81",
X"51f19b3f",
X"8151f1f8",
X"3f8251f1",
X"c23f8051",
X"f2a03f80",
X"c7a45280",
X"51c7f03f",
X"fdcc3f83",
X"e08c08fc",
X"05080d80",
X"0b83e080",
X"0c873d0d",
X"83e08c0c",
X"04fd3d0d",
X"75548074",
X"0c800b84",
X"150c800b",
X"88150c80",
X"e2dc0870",
X"3380e2e0",
X"08703370",
X"822a7081",
X"06703070",
X"72077009",
X"709f2c78",
X"069e0654",
X"51515451",
X"51555254",
X"51807298",
X"06525370",
X"882e0981",
X"06833881",
X"53709832",
X"70307080",
X"25757131",
X"84180c51",
X"51518072",
X"86065253",
X"70822e09",
X"81068338",
X"81537086",
X"32703070",
X"80257571",
X"31770c51",
X"51517194",
X"32703070",
X"80258817",
X"0c515185",
X"3d0d04fe",
X"3d0d7476",
X"54527151",
X"fee73f72",
X"812ea238",
X"8173268d",
X"3872822e",
X"ab387283",
X"2e9f38e6",
X"397108e2",
X"38841208",
X"dd388812",
X"08d838a0",
X"39881208",
X"812e0981",
X"06cc3894",
X"39881208",
X"812e8d38",
X"71088938",
X"84120880",
X"2effb738",
X"843d0d04",
X"fd3d0d75",
X"547383e3",
X"d0082ea7",
X"3880e3ec",
X"0874a00a",
X"07710c80",
X"e3fc0853",
X"53710851",
X"70802ef9",
X"3880730c",
X"71085170",
X"fb387383",
X"e3d00c85",
X"3d0d04ff",
X"0b83e3d0",
X"0c818080",
X"0b83e3cc",
X"0c800b83",
X"e0800c04",
X"fc3d0d76",
X"028405a2",
X"05220288",
X"05a60522",
X"7a545555",
X"55ff9d3f",
X"72802ea3",
X"3883e3cc",
X"08145271",
X"33757081",
X"05573481",
X"147083ff",
X"ff06ff15",
X"7083ffff",
X"06565255",
X"52da3980",
X"0b83e080",
X"0c863d0d",
X"04f73d0d",
X"7b7d7f11",
X"58555980",
X"5573762e",
X"b13883e3",
X"cc088b3d",
X"59577419",
X"703375fc",
X"06197008",
X"5d768306",
X"7b075354",
X"54517271",
X"3479720c",
X"81148116",
X"56547376",
X"2e098106",
X"d938800b",
X"83e0800c",
X"8b3d0d04",
X"fe3d0d80",
X"e3ec0883",
X"e3d00890",
X"0a07710c",
X"80e3fc08",
X"53537108",
X"5170802e",
X"f9388073",
X"0c710851",
X"70fb3884",
X"3d0d0483",
X"e08c0802",
X"83e08c0c",
X"fd3d0d80",
X"5383e08c",
X"088c0508",
X"5283e08c",
X"08880508",
X"5183d43f",
X"83e08008",
X"7083e080",
X"0c54853d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cfd",
X"3d0d8153",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"83a13f83",
X"e0800870",
X"83e0800c",
X"54853d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cf93d",
X"0d800b83",
X"e08c08fc",
X"050c83e0",
X"8c088805",
X"088025b9",
X"3883e08c",
X"08880508",
X"3083e08c",
X"0888050c",
X"800b83e0",
X"8c08f405",
X"0c83e08c",
X"08fc0508",
X"8a38810b",
X"83e08c08",
X"f4050c83",
X"e08c08f4",
X"050883e0",
X"8c08fc05",
X"0c83e08c",
X"088c0508",
X"8025b938",
X"83e08c08",
X"8c050830",
X"83e08c08",
X"8c050c80",
X"0b83e08c",
X"08f0050c",
X"83e08c08",
X"fc05088a",
X"38810b83",
X"e08c08f0",
X"050c83e0",
X"8c08f005",
X"0883e08c",
X"08fc050c",
X"805383e0",
X"8c088c05",
X"085283e0",
X"8c088805",
X"085181df",
X"3f83e080",
X"087083e0",
X"8c08f805",
X"0c5483e0",
X"8c08fc05",
X"08802e90",
X"3883e08c",
X"08f80508",
X"3083e08c",
X"08f8050c",
X"83e08c08",
X"f8050870",
X"83e0800c",
X"54893d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cfb3d",
X"0d800b83",
X"e08c08fc",
X"050c83e0",
X"8c088805",
X"08802599",
X"3883e08c",
X"08880508",
X"3083e08c",
X"0888050c",
X"810b83e0",
X"8c08fc05",
X"0c83e08c",
X"088c0508",
X"80259038",
X"83e08c08",
X"8c050830",
X"83e08c08",
X"8c050c81",
X"5383e08c",
X"088c0508",
X"5283e08c",
X"08880508",
X"51bd3f83",
X"e0800870",
X"83e08c08",
X"f8050c54",
X"83e08c08",
X"fc050880",
X"2e903883",
X"e08c08f8",
X"05083083",
X"e08c08f8",
X"050c83e0",
X"8c08f805",
X"087083e0",
X"800c5487",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"fd3d0d81",
X"0b83e08c",
X"08fc050c",
X"800b83e0",
X"8c08f805",
X"0c83e08c",
X"088c0508",
X"83e08c08",
X"88050827",
X"b93883e0",
X"8c08fc05",
X"08802eae",
X"38800b83",
X"e08c088c",
X"050824a2",
X"3883e08c",
X"088c0508",
X"1083e08c",
X"088c050c",
X"83e08c08",
X"fc050810",
X"83e08c08",
X"fc050cff",
X"b83983e0",
X"8c08fc05",
X"08802e80",
X"e13883e0",
X"8c088c05",
X"0883e08c",
X"08880508",
X"26ad3883",
X"e08c0888",
X"050883e0",
X"8c088c05",
X"083183e0",
X"8c088805",
X"0c83e08c",
X"08f80508",
X"83e08c08",
X"fc050807",
X"83e08c08",
X"f8050c83",
X"e08c08fc",
X"0508812a",
X"83e08c08",
X"fc050c83",
X"e08c088c",
X"0508812a",
X"83e08c08",
X"8c050cff",
X"953983e0",
X"8c089005",
X"08802e93",
X"3883e08c",
X"08880508",
X"7083e08c",
X"08f4050c",
X"51913983",
X"e08c08f8",
X"05087083",
X"e08c08f4",
X"050c5183",
X"e08c08f4",
X"050883e0",
X"800c853d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cff",
X"3d0d800b",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"05088106",
X"ff117009",
X"7083e08c",
X"088c0508",
X"0683e08c",
X"08fc0508",
X"1183e08c",
X"08fc050c",
X"83e08c08",
X"88050881",
X"2a83e08c",
X"0888050c",
X"83e08c08",
X"8c050810",
X"83e08c08",
X"8c050c51",
X"51515183",
X"e08c0888",
X"0508802e",
X"8438ffab",
X"3983e08c",
X"08fc0508",
X"7083e080",
X"0c51833d",
X"0d83e08c",
X"0c04fc3d",
X"0d767079",
X"7b555555",
X"558f7227",
X"8c387275",
X"07830651",
X"70802ea9",
X"38ff1252",
X"71ff2e98",
X"38727081",
X"05543374",
X"70810556",
X"34ff1252",
X"71ff2e09",
X"8106ea38",
X"7483e080",
X"0c863d0d",
X"04745172",
X"70840554",
X"08717084",
X"05530c72",
X"70840554",
X"08717084",
X"05530c72",
X"70840554",
X"08717084",
X"05530c72",
X"70840554",
X"08717084",
X"05530cf0",
X"1252718f",
X"26c93883",
X"72279538",
X"72708405",
X"54087170",
X"8405530c",
X"fc125271",
X"8326ed38",
X"7054ff81",
X"39000000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00002608",
X"00002649",
X"0000266a",
X"00002691",
X"00002691",
X"00002691",
X"00002754",
X"25732025",
X"73000000",
X"20000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"31364b00",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"43617274",
X"72696467",
X"65203332",
X"6b000000",
X"43617274",
X"72696467",
X"65203136",
X"6b206f6e",
X"65206368",
X"69700000",
X"43617274",
X"72696467",
X"65203136",
X"6b207477",
X"6f206368",
X"69700000",
X"45786974",
X"00000000",
X"61636964",
X"35323030",
X"2e726f6d",
X"00000000",
X"524f4d00",
X"42494e00",
X"43415200",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"0001e80a",
X"0001e809",
X"0001e80f",
X"0001d40e",
X"0001d403",
X"0001d402",
X"0001d400",
X"0001d401",
X"0001d409",
X"0001d301",
X"0001d300",
X"0001c010",
X"0001c01b",
X"0001c016",
X"0001c019",
X"0001c018",
X"0001c017",
X"0001c01a",
X"0004007c",
X"00040078",
X"00040074",
X"00040068",
X"00040060",
X"0004005c",
X"00040058",
X"00040054",
X"00040050",
X"0004004c",
X"00040048",
X"00040044",
X"00040040",
X"00040034",
X"00040030",
X"0004002c",
X"00040028",
X"00040024",
X"00040020",
X"0004001c",
X"00040018",
X"00040014",
X"00040010",
X"0004000c",
X"00040008",
X"00040004",
X"00040000",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
