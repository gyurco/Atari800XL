
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f4",
X"b0738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80f8",
X"cc0c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f1",
X"f12d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580f1b0",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80dbfc04",
X"fd3d0d75",
X"705254ae",
X"a73f83e0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83e0",
X"8008732e",
X"a13883e0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183e0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83e2c008",
X"248a38b4",
X"f83fff0b",
X"83e2c00c",
X"800b83e0",
X"800c04ff",
X"3d0d7352",
X"83e09c08",
X"722e8d38",
X"d93f7151",
X"96993f71",
X"83e09c0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"558154bc",
X"15088191",
X"387451cf",
X"3f795880",
X"7a2580f7",
X"3883e2f0",
X"0870892a",
X"5783ff06",
X"78848072",
X"31565657",
X"73782583",
X"38735575",
X"83e2c008",
X"2e8438ff",
X"893f83e2",
X"c0088025",
X"a6387589",
X"2b5198dc",
X"3f83e2f0",
X"088f3dfc",
X"11555c54",
X"8152f81b",
X"5196c63f",
X"761483e2",
X"f00c7583",
X"e2c00c74",
X"53765278",
X"51b3a93f",
X"83e08008",
X"83e2f008",
X"1683e2f0",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8b3861",
X"7a710c54",
X"75547580",
X"2e833881",
X"547383e0",
X"800c8e3d",
X"0d04fc3d",
X"0dfe9b3f",
X"7651feaf",
X"3f863dfc",
X"05537852",
X"775195e9",
X"3f797571",
X"0c5483e0",
X"80085483",
X"e0800880",
X"2e833881",
X"547383e0",
X"800c863d",
X"0d04fe3d",
X"0d7583e2",
X"c0085353",
X"80722489",
X"3871732e",
X"8438fdd6",
X"3f7451fd",
X"ea3f7251",
X"97ae3f83",
X"e0800852",
X"83e08008",
X"802e8338",
X"81527183",
X"e0800c84",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"e0800c51",
X"823d0d04",
X"80c40b83",
X"e0800c04",
X"fd3d0d75",
X"77715470",
X"535553a9",
X"ff3f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfceb3f",
X"735193ab",
X"3f7383e0",
X"9c0c83e0",
X"80085383",
X"e0800880",
X"2e833881",
X"537283e0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcbf3f",
X"72802ea5",
X"38bc1308",
X"527351a9",
X"893f83e0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"e0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83e0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83e2c0",
X"0c7483e0",
X"a00c7583",
X"e2bc0caf",
X"dd3f83e0",
X"800881ff",
X"06528153",
X"71993883",
X"e2d8518e",
X"943f83e0",
X"80085283",
X"e0800880",
X"2e833872",
X"52715372",
X"83e0800c",
X"843d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"51a6fa3f",
X"83e08008",
X"557483e0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"e0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283e2bc",
X"085180e0",
X"b33f83e0",
X"800857f9",
X"e13f7952",
X"83e2c451",
X"95b73f83",
X"e0800854",
X"805383e0",
X"8008732e",
X"09810682",
X"833883e0",
X"a0080b0b",
X"80f5e853",
X"705256a6",
X"b73f0b0b",
X"80f5e852",
X"80c01651",
X"a6aa3f75",
X"bc170c73",
X"82c0170c",
X"810b82c4",
X"170c810b",
X"82c8170c",
X"7382cc17",
X"0cff1782",
X"d0175557",
X"81913983",
X"e0ac3370",
X"822a7081",
X"06515455",
X"72818038",
X"74812a81",
X"06587780",
X"f6387484",
X"2a810682",
X"c4150c83",
X"e0ac3381",
X"0682c815",
X"0c795273",
X"51a5d13f",
X"7351a5e8",
X"3f83e080",
X"081453af",
X"73708105",
X"553472bc",
X"150c83e0",
X"ad527251",
X"a5b23f83",
X"e0a40882",
X"c0150c83",
X"e0ba5280",
X"c01451a5",
X"9f3f7880",
X"2e8d3873",
X"51782d83",
X"e0800880",
X"2e993877",
X"82cc150c",
X"75802e86",
X"387382cc",
X"170c7382",
X"d015ff19",
X"59555676",
X"802e9b38",
X"83e0a452",
X"83e2c451",
X"94ad3f83",
X"e080088a",
X"3883e0ad",
X"335372fe",
X"d2387880",
X"2e893883",
X"e0a00851",
X"fcb83f83",
X"e0a00853",
X"7283e080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb53f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f690",
X"3f83e080",
X"08745387",
X"3d705355",
X"55f6b03f",
X"f7903f73",
X"51d33f63",
X"53745283",
X"e0800851",
X"fab83f92",
X"3d0d0471",
X"83e0800c",
X"0480c012",
X"83e0800c",
X"04803d0d",
X"7282c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"e0800c51",
X"823d0d04",
X"f93d0d79",
X"83e09008",
X"57578177",
X"27819638",
X"76881708",
X"27818e38",
X"75335574",
X"822e8938",
X"74832eb3",
X"3880fe39",
X"74547610",
X"83fe0653",
X"76882a8c",
X"17080552",
X"893dfc05",
X"51aa8b3f",
X"83e08008",
X"80df3802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d13984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"51a9db3f",
X"83e08008",
X"b038029f",
X"05330284",
X"059e0533",
X"71982b71",
X"902b0702",
X"8c059d05",
X"3370882b",
X"72078d3d",
X"337180ff",
X"fffe8006",
X"07515253",
X"57585683",
X"39815574",
X"83e0800c",
X"893d0d04",
X"fb3d0d83",
X"e09008fe",
X"19881208",
X"fe055556",
X"54805674",
X"73278d38",
X"82143375",
X"71299416",
X"08055753",
X"7583e080",
X"0c873d0d",
X"04fc3d0d",
X"7652800b",
X"83e09008",
X"70335152",
X"5370832e",
X"09810691",
X"38951233",
X"94133371",
X"982b7190",
X"2b075555",
X"519b1233",
X"9a133371",
X"882b0774",
X"0783e080",
X"0c55863d",
X"0d04fc3d",
X"0d7683e0",
X"90085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"fed63f83",
X"e0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183e080",
X"0c863d0d",
X"04fa3d0d",
X"7883e090",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fcb13f",
X"81527183",
X"e0800827",
X"a8388352",
X"83e08008",
X"88170827",
X"9c3883e0",
X"80088c16",
X"0c83e080",
X"0851fdbc",
X"3f83e080",
X"0890160c",
X"73752380",
X"527183e0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585e5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"9f269138",
X"7a51fdd2",
X"3f83e080",
X"0856807d",
X"34838139",
X"933d841c",
X"08705859",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"3880705a",
X"5c887f08",
X"5f5a7b81",
X"1d7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535e57",
X"557480e7",
X"3876ae2e",
X"09810683",
X"38815578",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675bb",
X"3888598b",
X"5affab39",
X"76982b55",
X"74802587",
X"3880f3c0",
X"173357ff",
X"9f175574",
X"99268938",
X"e0177081",
X"ff065855",
X"78811a70",
X"81ff0672",
X"1b535b57",
X"55767534",
X"fef8397b",
X"1e7f0c80",
X"5576a026",
X"83388155",
X"748b1934",
X"7a51fc82",
X"3f83e080",
X"0880f538",
X"a0547a22",
X"70852b83",
X"e0065455",
X"901b0852",
X"7c51a496",
X"3f83e080",
X"085783e0",
X"80088181",
X"387c3355",
X"74802e80",
X"f4388b1d",
X"3370832a",
X"70810651",
X"565674b4",
X"388b7d84",
X"1d0883e0",
X"8008595b",
X"5b58ff18",
X"5877ff2e",
X"9a387970",
X"81055b33",
X"79708105",
X"5b337171",
X"31525656",
X"75802ee2",
X"38863975",
X"802e9638",
X"7a51fbe5",
X"3fff8639",
X"83e08008",
X"5683e080",
X"08b63883",
X"39765684",
X"1b088b11",
X"33515574",
X"a7388b1d",
X"3370842a",
X"70810651",
X"56567489",
X"38835694",
X"39815690",
X"397c51fa",
X"943f83e0",
X"8008881c",
X"0cfd8139",
X"7583e080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"51a2db3f",
X"835683e0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"51a2af3f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"7651a286",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583e080",
X"0c8a3d0d",
X"04eb3d0d",
X"675a800b",
X"83e0900c",
X"a1a83f83",
X"e0800881",
X"06558256",
X"7483ef38",
X"7475538f",
X"3d705357",
X"59feca3f",
X"83e08008",
X"81ff0657",
X"76812e09",
X"810680d4",
X"38905483",
X"be537452",
X"7551a19a",
X"3f83e080",
X"0880c938",
X"8f3d3355",
X"74802e80",
X"c93802bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"33710770",
X"587b575e",
X"525e5759",
X"57fdee3f",
X"83e08008",
X"81ff0657",
X"76832e09",
X"81068638",
X"815682f2",
X"3976802e",
X"86388656",
X"82e839a4",
X"548d5378",
X"527551a0",
X"b13f8156",
X"83e08008",
X"82d43802",
X"be053302",
X"8405bd05",
X"3371882b",
X"07595d77",
X"ab380280",
X"ce053302",
X"840580cd",
X"05337198",
X"2b71902b",
X"07973d33",
X"70882b72",
X"07029405",
X"80cb0533",
X"71075452",
X"5e575956",
X"02b70533",
X"78712902",
X"8805b605",
X"33028c05",
X"b5053371",
X"882b0770",
X"1d707f8c",
X"050c5f59",
X"57595d8e",
X"3d33821b",
X"3402b905",
X"33903d33",
X"71882b07",
X"5a5c7884",
X"1b2302bb",
X"05330284",
X"05ba0533",
X"71882b07",
X"565c74ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"07515253",
X"575e5c74",
X"76317831",
X"79842a90",
X"3d335471",
X"71315356",
X"5680d198",
X"3f83e080",
X"08820570",
X"881c0c83",
X"e08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83e0900c",
X"80567583",
X"e0800c97",
X"3d0d04e9",
X"3d0d83e0",
X"90085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e53f83e0",
X"80085483",
X"e0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f489",
X"3f83e080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383e080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83e09008",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0e93f",
X"83e08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"833f83e0",
X"80085583",
X"e0800880",
X"2eff8938",
X"83e08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"519ad73f",
X"83e08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83e0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83e09008",
X"55568555",
X"73802e81",
X"e3388114",
X"33810653",
X"84557280",
X"2e81d538",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b9388214",
X"3370892b",
X"56537680",
X"2eb73874",
X"52ff1651",
X"80cc993f",
X"83e08008",
X"ff187654",
X"70535853",
X"80cc893f",
X"83e08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed63f83",
X"e0800853",
X"810b83e0",
X"8008278b",
X"38881408",
X"83e08008",
X"26883880",
X"0b811534",
X"b03983e0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc53f",
X"83e08008",
X"8c3883e0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683e0",
X"800805a8",
X"150c8055",
X"7483e080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83e09008",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1cf3f",
X"83e08008",
X"5583e080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef5",
X"3f83e080",
X"0888170c",
X"7551efa6",
X"3f83e080",
X"08557483",
X"e0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683e0",
X"9008802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f53f83e0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"96e03f83",
X"e0800841",
X"83e08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"eddf3f83",
X"e0800841",
X"83e08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"8e863f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f03f83e0",
X"80088332",
X"70307072",
X"079f2c83",
X"e0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"8c923f75",
X"83e0800c",
X"9e3d0d04",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"7751e0d2",
X"3f83e080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3380f8d4",
X"0b80f8d4",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"527751e0",
X"813f83e0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583e0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"558b993f",
X"83e08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"8114518a",
X"b13f83e0",
X"80083070",
X"83e08008",
X"07802583",
X"e0800c53",
X"863d0d04",
X"fc3d0d76",
X"705255e6",
X"ee3f83e0",
X"80085481",
X"5383e080",
X"0880c138",
X"7451e6b1",
X"3f83e080",
X"0880f5f8",
X"5383e080",
X"085253ff",
X"913f83e0",
X"8008a138",
X"80f5fc52",
X"7251ff82",
X"3f83e080",
X"08923880",
X"f6805272",
X"51fef33f",
X"83e08008",
X"802e8338",
X"81547353",
X"7283e080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"e68d3f81",
X"5383e080",
X"08983873",
X"51e5d63f",
X"83e38808",
X"5283e080",
X"0851feba",
X"3f83e080",
X"08537283",
X"e0800c85",
X"3d0d04df",
X"3d0da43d",
X"0870525e",
X"dbfb3f83",
X"e0800833",
X"953d5654",
X"73963880",
X"fc905274",
X"5189913f",
X"9a397d52",
X"7851defc",
X"3f84d039",
X"7d51dbe1",
X"3f83e080",
X"08527451",
X"db913f80",
X"43804280",
X"41804083",
X"e3900852",
X"943d7052",
X"5de1e43f",
X"83e08008",
X"59800b83",
X"e0800855",
X"5b83e080",
X"087b2e94",
X"38811b74",
X"525be4e6",
X"3f83e080",
X"085483e0",
X"8008ee38",
X"805aff5f",
X"7909709f",
X"2c7b065b",
X"547a7a24",
X"8438ff1b",
X"5af61a70",
X"09709f2c",
X"72067bff",
X"125a5a52",
X"55558075",
X"25953876",
X"51e4ab3f",
X"83e08008",
X"76ff1858",
X"55577380",
X"24ed3874",
X"7f2e8638",
X"a0bd3f74",
X"5f78ff1b",
X"70585d58",
X"807a2595",
X"387751e4",
X"813f83e0",
X"800876ff",
X"18585558",
X"738024ed",
X"38800b83",
X"e7c00c80",
X"0b83e7e4",
X"0c80f684",
X"518d903f",
X"81800b83",
X"e7e40c80",
X"f68c518d",
X"823fa80b",
X"83e7c00c",
X"76802e80",
X"e43883e7",
X"c0087779",
X"32703070",
X"72078025",
X"70872b83",
X"e7e40c51",
X"56785356",
X"56e3b83f",
X"83e08008",
X"802e8838",
X"80f69451",
X"8cc93f76",
X"51e2fa3f",
X"83e08008",
X"5280f7b4",
X"518cb83f",
X"7651e382",
X"3f83e080",
X"0883e7c0",
X"08555775",
X"74258638",
X"a81656f7",
X"397583e7",
X"c00c86f0",
X"7624ff98",
X"3887980b",
X"83e7c00c",
X"77802eb1",
X"387751e2",
X"b83f83e0",
X"80087852",
X"55e2d83f",
X"80f69c54",
X"83e08008",
X"8d388739",
X"80763481",
X"d03980f6",
X"98547453",
X"735280f5",
X"ec518bd7",
X"3f805480",
X"f5f4518b",
X"ce3f8114",
X"5473a82e",
X"098106ef",
X"38868da0",
X"519cb03f",
X"8052903d",
X"70525780",
X"c1eb3f83",
X"52765180",
X"c1e33f62",
X"818f3861",
X"802e80fb",
X"387b5473",
X"ff2e9638",
X"78802e81",
X"8a387851",
X"e1dc3f83",
X"e08008ff",
X"155559e7",
X"3978802e",
X"80f53878",
X"51e1d83f",
X"83e08008",
X"802efc8e",
X"387851e1",
X"a03f83e0",
X"80085280",
X"f5e85183",
X"e43f83e0",
X"8008a338",
X"7c51859c",
X"3f83e080",
X"085574ff",
X"16565480",
X"7425ae38",
X"741d7033",
X"555673af",
X"2efecd38",
X"e9397851",
X"e0e13f83",
X"e0800852",
X"7c5184d4",
X"3f8f397f",
X"88296010",
X"057a0561",
X"055afc90",
X"3962802e",
X"fbd13880",
X"52765180",
X"c0c33fa3",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067084",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d38a8",
X"0b9088b8",
X"34b80b90",
X"88b83470",
X"83e0800c",
X"823d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"852a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"980b9088",
X"b834b80b",
X"9088b834",
X"7083e080",
X"0c823d0d",
X"04930b90",
X"88bc34ff",
X"0b9088a8",
X"3404ff3d",
X"0d028f05",
X"3352800b",
X"9088bc34",
X"8a5199f7",
X"3fdf3f80",
X"f80b9088",
X"a034800b",
X"90888834",
X"fa125271",
X"90888034",
X"800b9088",
X"98347190",
X"88903490",
X"88b85280",
X"7234b872",
X"34833d0d",
X"04803d0d",
X"028b0533",
X"51709088",
X"b434febf",
X"3f83e080",
X"08802ef6",
X"38823d0d",
X"04803d0d",
X"8439a4ae",
X"3ffed93f",
X"83e08008",
X"802ef338",
X"9088b433",
X"7081ff06",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"a30b9088",
X"bc34ff0b",
X"9088a834",
X"9088b851",
X"a87134b8",
X"7134823d",
X"0d04803d",
X"0d9088bc",
X"337081c0",
X"06703070",
X"802583e0",
X"800c5151",
X"51823d0d",
X"04803d0d",
X"9088b833",
X"7081ff06",
X"70832a81",
X"32708106",
X"51515151",
X"70802ee8",
X"38b00b90",
X"88b834b8",
X"0b9088b8",
X"34823d0d",
X"04803d0d",
X"9080ac08",
X"810683e0",
X"800c823d",
X"0d04fd3d",
X"0d757754",
X"54807325",
X"94387370",
X"81055533",
X"5280f6a0",
X"5187843f",
X"ff1353e9",
X"39853d0d",
X"04fd3d0d",
X"75775354",
X"73335170",
X"89387133",
X"5170802e",
X"a1387333",
X"72335253",
X"72712785",
X"38ff5194",
X"39707327",
X"85388151",
X"8b398114",
X"81135354",
X"d3398051",
X"7083e080",
X"0c853d0d",
X"04fd3d0d",
X"75775454",
X"72337081",
X"ff065252",
X"70802ea3",
X"387181ff",
X"068114ff",
X"bf125354",
X"52709926",
X"8938a012",
X"7081ff06",
X"53517174",
X"70810556",
X"34d23980",
X"7434853d",
X"0d04ffbd",
X"3d0d80c6",
X"3d0852a5",
X"3d705254",
X"ffb33f80",
X"c73d0852",
X"853d7052",
X"53ffa63f",
X"72527351",
X"fedf3f80",
X"c53d0d04",
X"fe3d0d74",
X"76535371",
X"70810553",
X"33517073",
X"70810555",
X"3470f038",
X"843d0d04",
X"fe3d0d74",
X"52807233",
X"52537073",
X"2e8d3881",
X"12811471",
X"33535452",
X"70f53872",
X"83e0800c",
X"843d0d04",
X"f63d0d7c",
X"7e60625a",
X"5d5b5680",
X"59815585",
X"39747a29",
X"55745275",
X"51b8ed3f",
X"83e08008",
X"7a27ee38",
X"74802e80",
X"dd387452",
X"7551b8d8",
X"3f83e080",
X"08755376",
X"5254b8dc",
X"3f83e080",
X"087a5375",
X"5256b8c0",
X"3f83e080",
X"08793070",
X"7b079f2a",
X"70778024",
X"07515154",
X"55728738",
X"83e08008",
X"c5387681",
X"18b01655",
X"58588974",
X"258b38b7",
X"14537a85",
X"3880d714",
X"53727834",
X"811959ff",
X"9f398077",
X"348c3d0d",
X"04f73d0d",
X"7b7d7f62",
X"029005bb",
X"05335759",
X"565a5ab0",
X"58728338",
X"a0587570",
X"70810552",
X"33715954",
X"55903980",
X"74258e38",
X"ff147770",
X"81055933",
X"545472ef",
X"3873ff15",
X"55538073",
X"25893877",
X"52795178",
X"2def3975",
X"33755753",
X"72802e90",
X"38725279",
X"51782d75",
X"70810557",
X"3353ed39",
X"8b3d0d04",
X"ee3d0d64",
X"66696970",
X"70810552",
X"335b4a5c",
X"5e5e7680",
X"2e82f938",
X"76a52e09",
X"810682e0",
X"38807041",
X"67707081",
X"05523371",
X"4a59575f",
X"76b02e09",
X"81068c38",
X"75708105",
X"57337648",
X"57815fd0",
X"17567589",
X"2680da38",
X"76675c59",
X"805c9339",
X"778a2480",
X"c3387b8a",
X"29187b70",
X"81055d33",
X"5a5cd019",
X"7081ff06",
X"58588977",
X"27a438ff",
X"9f197081",
X"ff06ffa9",
X"1b5a5156",
X"85762792",
X"38ffbf19",
X"7081ff06",
X"51567585",
X"268a38c9",
X"19587780",
X"25ffb938",
X"7a477b40",
X"7881ff06",
X"577680e4",
X"2e80e538",
X"7680e424",
X"a7387680",
X"d82e8186",
X"387680d8",
X"24903876",
X"802e81cc",
X"3876a52e",
X"81b63881",
X"b9397680",
X"e32e818c",
X"3881af39",
X"7680f52e",
X"9b387680",
X"f5248b38",
X"7680f32e",
X"81813881",
X"99397680",
X"f82e80ca",
X"38818f39",
X"913d7055",
X"5780538a",
X"5279841b",
X"7108535b",
X"56fc813f",
X"7655ab39",
X"79841b71",
X"08943d70",
X"5b5b525b",
X"56758025",
X"8c387530",
X"56ad7834",
X"0280c105",
X"57765480",
X"538a5275",
X"51fbd53f",
X"77557e54",
X"b839913d",
X"70557780",
X"d8327030",
X"70802556",
X"51585690",
X"5279841b",
X"7108535b",
X"57fbb13f",
X"7555db39",
X"79841b83",
X"1233545b",
X"56983979",
X"841b7108",
X"575b5680",
X"547f537c",
X"527d51fc",
X"9c3f8739",
X"76527d51",
X"7c2d6670",
X"33588105",
X"47fd8339",
X"943d0d04",
X"7283e094",
X"0c7183e0",
X"980c04fb",
X"3d0d883d",
X"70708405",
X"52085754",
X"755383e0",
X"94085283",
X"e0980851",
X"fcc63f87",
X"3d0d04ff",
X"3d0d7370",
X"08535102",
X"93053372",
X"34700881",
X"05710c83",
X"3d0d04fc",
X"3d0d873d",
X"88115578",
X"54bdbb53",
X"51fc993f",
X"8052873d",
X"51d13f86",
X"3d0d04fc",
X"3d0d7655",
X"7483e398",
X"082eaf38",
X"80537451",
X"87c13f83",
X"e0800881",
X"ff06ff14",
X"7081ff06",
X"7230709f",
X"2a515255",
X"53547280",
X"2e843871",
X"dd3873fe",
X"387483e3",
X"980c863d",
X"0d04ff3d",
X"0dff0b83",
X"e3980c84",
X"a53f8151",
X"87853f83",
X"e0800881",
X"ff065271",
X"ee3881d3",
X"3f7183e0",
X"800c833d",
X"0d04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"823f7280",
X"2ea03883",
X"e3ac1433",
X"75708105",
X"57348114",
X"7083ffff",
X"06ff1570",
X"83ffff06",
X"56525552",
X"dd39800b",
X"83e0800c",
X"863d0d04",
X"fc3d0d76",
X"787a1156",
X"53558053",
X"71742e93",
X"38721551",
X"703383e3",
X"ac133481",
X"12811454",
X"52ea3980",
X"0b83e080",
X"0c863d0d",
X"04fd3d0d",
X"905483e3",
X"98085186",
X"f43f83e0",
X"800881ff",
X"06ff1571",
X"30713070",
X"73079f2a",
X"729f2a06",
X"52555255",
X"5372db38",
X"853d0d04",
X"803d0d83",
X"e3a40810",
X"83e39c08",
X"079080a8",
X"0c823d0d",
X"04800b83",
X"e3a40ce4",
X"3f04810b",
X"83e3a40c",
X"db3f04ed",
X"3f047183",
X"e3a00c04",
X"803d0d80",
X"51f43f81",
X"0b83e3a4",
X"0c810b83",
X"e39c0cff",
X"bb3f823d",
X"0d04803d",
X"0d723070",
X"74078025",
X"83e39c0c",
X"51ffa53f",
X"823d0d04",
X"803d0d02",
X"8b053390",
X"80a40c90",
X"80a80870",
X"81065151",
X"70f53890",
X"80a40870",
X"81ff0683",
X"e0800c51",
X"823d0d04",
X"803d0d81",
X"ff51d13f",
X"83e08008",
X"81ff0683",
X"e0800c82",
X"3d0d0480",
X"3d0d7390",
X"2b730790",
X"80b40c82",
X"3d0d0404",
X"fb3d0d78",
X"0284059f",
X"05337098",
X"2b555755",
X"7280259b",
X"387580ff",
X"06568052",
X"80f751e0",
X"3f83e080",
X"0881ff06",
X"54738126",
X"80ff3880",
X"51fee73f",
X"ffa23f81",
X"51fedf3f",
X"ff9a3f75",
X"51feed3f",
X"74982a51",
X"fee63f74",
X"902a7081",
X"ff065253",
X"feda3f74",
X"882a7081",
X"ff065253",
X"fece3f74",
X"81ff0651",
X"fec63f81",
X"557580c0",
X"2e098106",
X"86388195",
X"558d3975",
X"80c82e09",
X"81068438",
X"81875574",
X"51fea53f",
X"8a55fec8",
X"3f83e080",
X"0881ff06",
X"70982b54",
X"54728025",
X"8c38ff15",
X"7081ff06",
X"565374e2",
X"387383e0",
X"800c873d",
X"0d04fa3d",
X"0dfdc53f",
X"8051fdda",
X"3f8a54fe",
X"933fff14",
X"7081ff06",
X"555373f3",
X"38737453",
X"5580c051",
X"fea63f83",
X"e0800881",
X"ff065473",
X"812e0981",
X"06829f38",
X"83aa5280",
X"c851fe8c",
X"3f83e080",
X"0881ff06",
X"5372812e",
X"09810681",
X"a8387454",
X"873d7411",
X"5456fdc8",
X"3f83e080",
X"08733481",
X"147081ff",
X"06555383",
X"7427e538",
X"029a0533",
X"5372812e",
X"09810681",
X"d938029b",
X"05335380",
X"ce905472",
X"81aa2e8d",
X"3881c739",
X"80e4518a",
X"9e3fff14",
X"5473802e",
X"81b83882",
X"0a5281e9",
X"51fda53f",
X"83e08008",
X"81ff0653",
X"72de3872",
X"5280fa51",
X"fd923f83",
X"e0800881",
X"ff065372",
X"81903872",
X"54731653",
X"fcd63f83",
X"e0800873",
X"34811470",
X"81ff0655",
X"53837427",
X"e838873d",
X"3370862a",
X"70810651",
X"54548c55",
X"7280e338",
X"845580de",
X"39745281",
X"e951fccc",
X"3f83e080",
X"0881ff06",
X"53825581",
X"e9568173",
X"27863873",
X"5580c156",
X"80ce9054",
X"8a3980e4",
X"5189903f",
X"ff145473",
X"802ea938",
X"80527551",
X"fc9a3f83",
X"e0800881",
X"ff065372",
X"e1388480",
X"5280d051",
X"fc863f83",
X"e0800881",
X"ff065372",
X"802e8338",
X"80557483",
X"e3a83480",
X"51fb873f",
X"fbc23f88",
X"3d0d04fb",
X"3d0d7754",
X"800b83e3",
X"a8337083",
X"2a708106",
X"51555755",
X"72752e09",
X"81068538",
X"73892b54",
X"735280d1",
X"51fbbd3f",
X"83e08008",
X"81ff0653",
X"72bd3882",
X"b8c054fb",
X"833f83e0",
X"800881ff",
X"06537281",
X"ff2e0981",
X"068938ff",
X"145473e7",
X"389f3972",
X"81fe2e09",
X"81069638",
X"83e7ac52",
X"83e3ac51",
X"faed3ffa",
X"d33ffad0",
X"3f833981",
X"558051fa",
X"893ffac4",
X"3f7481ff",
X"0683e080",
X"0c873d0d",
X"04fb3d0d",
X"7783e3ac",
X"56548151",
X"f9ec3f83",
X"e3a83370",
X"832a7081",
X"06515456",
X"72853873",
X"892b5473",
X"5280d851",
X"fab63f83",
X"e0800881",
X"ff065372",
X"80e43881",
X"ff51f9d4",
X"3f81fe51",
X"f9ce3f84",
X"80537470",
X"81055633",
X"51f9c13f",
X"ff137083",
X"ffff0651",
X"5372eb38",
X"7251f9b0",
X"3f7251f9",
X"ab3ff9d0",
X"3f83e080",
X"089f0653",
X"a7885472",
X"852e8c38",
X"993980e4",
X"5186c83f",
X"ff1454f9",
X"b33f83e0",
X"800881ff",
X"2e843873",
X"e9388051",
X"f8e43ff9",
X"9f3f800b",
X"83e0800c",
X"873d0d04",
X"7183e7b0",
X"0c888080",
X"0b83e7ac",
X"0c848080",
X"0b83e7b4",
X"0c04fd3d",
X"0d777017",
X"557705ff",
X"1a535371",
X"ff2e9438",
X"73708105",
X"55335170",
X"73708105",
X"5534ff12",
X"52e93985",
X"3d0d04fc",
X"3d0d87a6",
X"81557433",
X"83e7b834",
X"a05483a0",
X"805383e7",
X"b0085283",
X"e7ac0851",
X"ffb83fa0",
X"5483a480",
X"5383e7b0",
X"085283e7",
X"ac0851ff",
X"a53f9054",
X"83a88053",
X"83e7b008",
X"5283e7ac",
X"0851ff92",
X"3fa05380",
X"5283e7b4",
X"0883a080",
X"055185a0",
X"3fa05380",
X"5283e7b4",
X"0883a480",
X"05518590",
X"3f905380",
X"5283e7b4",
X"0883a880",
X"05518580",
X"3fff7534",
X"83a08054",
X"805383e7",
X"b0085283",
X"e7b40851",
X"fecc3f80",
X"d0805483",
X"b0805383",
X"e7b00852",
X"83e7b408",
X"51feb73f",
X"86c53fa2",
X"54805383",
X"e7b4088c",
X"80055280",
X"f9c851fe",
X"a13f860b",
X"87a88334",
X"800b87a8",
X"8234800b",
X"87a09a34",
X"af0b87a0",
X"9634bf0b",
X"87a09734",
X"800b87a0",
X"98349f0b",
X"87a09934",
X"800b87a0",
X"9b34e00b",
X"87a88934",
X"a20b87a8",
X"8034830b",
X"87a48f34",
X"820b87a8",
X"8134863d",
X"0d04fd3d",
X"0d83a080",
X"54805383",
X"e7b40852",
X"83e7b008",
X"51fdbf3f",
X"80d08054",
X"83b08053",
X"83e7b408",
X"5283e7b0",
X"0851fdaa",
X"3fa05483",
X"a0805383",
X"e7b40852",
X"83e7b008",
X"51fd973f",
X"a05483a4",
X"805383e7",
X"b4085283",
X"e7b00851",
X"fd843f90",
X"5483a880",
X"5383e7b4",
X"085283e7",
X"b00851fc",
X"f13f83e7",
X"b83387a6",
X"8134853d",
X"0d04803d",
X"0d908090",
X"08810683",
X"e0800c82",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe067607",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"812c8106",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fd06",
X"76100772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087082",
X"2cbf0683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fe8306",
X"76822b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"882c8706",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f1ff",
X"0676882b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70912cbf",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870fc",
X"87ffff06",
X"76912b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"992c8106",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870ffbf",
X"0a067699",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908080",
X"0870882c",
X"810683e0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"80087089",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8a2c8106",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708b2c81",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708c2c",
X"bf0683e0",
X"800c5182",
X"3d0d04fe",
X"3d0d7481",
X"e629872a",
X"9080a00c",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d848080",
X"53805288",
X"800a51ff",
X"b33f8180",
X"80538052",
X"82800a51",
X"c63f843d",
X"0d04803d",
X"0d8151fc",
X"aa3f7280",
X"2e903880",
X"51fdfe3f",
X"cd3f83e7",
X"bc3351fd",
X"f43f8151",
X"fcbb3f80",
X"51fcb63f",
X"8051fc87",
X"3f823d0d",
X"04fd3d0d",
X"75528054",
X"80ff7225",
X"8838810b",
X"ff801353",
X"54ffbf12",
X"51709926",
X"8638e012",
X"52b039ff",
X"9f125199",
X"7127a738",
X"d012e013",
X"54517089",
X"26853872",
X"52983972",
X"8f268538",
X"72528f39",
X"71ba2e09",
X"81068538",
X"9a528339",
X"80527380",
X"2e853881",
X"80125271",
X"81ff0683",
X"e0800c85",
X"3d0d0480",
X"3d0d84d8",
X"c0518071",
X"70810553",
X"347084e0",
X"c02e0981",
X"06f03882",
X"3d0d04fe",
X"3d0d0297",
X"053351fe",
X"f43f83e0",
X"800881ff",
X"0683e7c0",
X"08545280",
X"73249b38",
X"83e7e008",
X"137283e7",
X"e4080753",
X"53717334",
X"83e7c008",
X"810583e7",
X"c00c843d",
X"0d04fa3d",
X"0d82800a",
X"1b558057",
X"883dfc05",
X"54795374",
X"527851ff",
X"bba43f88",
X"3d0d04fe",
X"3d0d83e7",
X"d8085274",
X"51c2883f",
X"83e08008",
X"8c387653",
X"755283e7",
X"d80851c6",
X"3f843d0d",
X"04fe3d0d",
X"83e7d808",
X"53755274",
X"51ffbcc6",
X"3f83e080",
X"088d3877",
X"53765283",
X"e7d80851",
X"ffa03f84",
X"3d0d04fe",
X"3d0d83e7",
X"d80851ff",
X"bbb93f83",
X"e0800881",
X"80802e09",
X"81068838",
X"83c18080",
X"539c3983",
X"e7d80851",
X"ffbb9c3f",
X"83e08008",
X"80d0802e",
X"09810693",
X"3883c1b0",
X"805383e0",
X"80085283",
X"e7d80851",
X"fed43f84",
X"3d0d0480",
X"3d0df9fc",
X"3f83e080",
X"08842980",
X"f9ec0570",
X"0883e080",
X"0c51823d",
X"0d04ed3d",
X"0d804480",
X"43804280",
X"4180705a",
X"5bfdcc3f",
X"800b83e7",
X"c00c800b",
X"83e7e40c",
X"80f6ec51",
X"eac13f81",
X"800b83e7",
X"e40c80f6",
X"f051eab3",
X"3f80d00b",
X"83e7c00c",
X"7830707a",
X"07802570",
X"872b83e7",
X"e40c5155",
X"f8ed3f83",
X"e0800852",
X"80f6f851",
X"ea8d3f80",
X"f80b83e7",
X"c00c7881",
X"32703070",
X"72078025",
X"70872b83",
X"e7e40c51",
X"56569cfa",
X"3f83e080",
X"085280f7",
X"8851e9e3",
X"3f81a00b",
X"83e7c00c",
X"78823270",
X"30707207",
X"80257087",
X"2b83e7e4",
X"0c515656",
X"fec53f83",
X"e0800852",
X"80f79851",
X"e9b93f81",
X"c80b83e7",
X"c00c7883",
X"32703070",
X"72078025",
X"70872b83",
X"e7e40c51",
X"5683e7d8",
X"085256ff",
X"b6973f83",
X"e0800852",
X"80f7a051",
X"e9893f82",
X"980b83e7",
X"c00c810b",
X"83e7c45b",
X"5883e7c0",
X"0883197a",
X"32703070",
X"72078025",
X"70872b83",
X"e7e40c51",
X"578e3d70",
X"55ff1b54",
X"5757579a",
X"bc3f7970",
X"84055b08",
X"51ffb5cd",
X"3f745483",
X"e0800853",
X"775280f7",
X"a851e8bb",
X"3fa81783",
X"e7c00c81",
X"18587785",
X"2e098106",
X"ffaf3883",
X"b80b83e7",
X"c00c7888",
X"32703070",
X"72078025",
X"70872b83",
X"e7e40c51",
X"5656f7b9",
X"3f80f7b8",
X"5583e080",
X"08802e8f",
X"3883e7d4",
X"0851ffb4",
X"f83f83e0",
X"80085574",
X"5280f7c0",
X"51e7e83f",
X"84880b83",
X"e7c00c78",
X"89327030",
X"70720780",
X"2570872b",
X"83e7e40c",
X"515780f7",
X"cc5255e7",
X"c63f868d",
X"a051f8b3",
X"3f805291",
X"3d705255",
X"9def3f83",
X"5274519d",
X"e83f6355",
X"74839c38",
X"61195978",
X"80258538",
X"74599039",
X"89792585",
X"38885987",
X"39788926",
X"82fb3878",
X"822b5580",
X"f5c01508",
X"04f5d43f",
X"83e08008",
X"61575575",
X"812e0981",
X"06893883",
X"e0800810",
X"55903975",
X"ff2e0981",
X"06883883",
X"e0800881",
X"2c559075",
X"25853890",
X"55883974",
X"80248338",
X"81557451",
X"f5ae3f82",
X"b03999c1",
X"3f83e080",
X"08610555",
X"74802585",
X"38805588",
X"39877525",
X"83388755",
X"74518da4",
X"3f828e39",
X"f59e3f83",
X"e0800861",
X"05557480",
X"25853880",
X"55883986",
X"75258338",
X"86557451",
X"f5973f81",
X"ec396087",
X"3862802e",
X"81e33883",
X"e38c0883",
X"e3880cad",
X"e50b83e3",
X"900c83e7",
X"d80851d6",
X"da3ffa8f",
X"3f81c639",
X"60568076",
X"259838ad",
X"840b83e3",
X"900c83e7",
X"b4157008",
X"5255d6bb",
X"3f740852",
X"92397580",
X"25923883",
X"e7b41508",
X"51ffb2bf",
X"3f8052fc",
X"1951b839",
X"62802e81",
X"8c3883e7",
X"b4157008",
X"83e7c408",
X"720c83e7",
X"c40cfc1a",
X"70535155",
X"8bf13f83",
X"e0800856",
X"80518be7",
X"3f83e080",
X"08527451",
X"88803f75",
X"52805187",
X"f93f80d5",
X"39605580",
X"7525b638",
X"83e39408",
X"83e3880c",
X"ade50b83",
X"e3900c83",
X"e7d40851",
X"d5c53f83",
X"e7d40851",
X"d2e63f83",
X"e0800881",
X"ff067052",
X"55f3f73f",
X"74802e9d",
X"388155a1",
X"39748025",
X"943883e7",
X"d40851ff",
X"b1b13f80",
X"51f3db3f",
X"84396287",
X"387a802e",
X"f9b73880",
X"557483e0",
X"800c953d",
X"0d04fe3d",
X"0df4873f",
X"83e08008",
X"802e8638",
X"8051818a",
X"39f48c3f",
X"83e08008",
X"80fe38f4",
X"ac3f83e0",
X"8008802e",
X"b9388151",
X"f1e93f80",
X"51f3c23f",
X"eedd3f80",
X"0b83e7c0",
X"0cf8df3f",
X"83e08008",
X"53ff0b83",
X"e7c00cf0",
X"c93f7280",
X"cb3883e7",
X"bc3351f3",
X"9c3f7251",
X"f1b93f80",
X"c039f3d4",
X"3f83e080",
X"08802eb5",
X"388151f1",
X"a63f8051",
X"f2ff3fee",
X"9a3fad84",
X"0b83e390",
X"0c83e7c4",
X"0851d3f7",
X"3fff0b83",
X"e7c00cf0",
X"853f83e7",
X"c4085280",
X"5185f73f",
X"8151f4c6",
X"3f843d0d",
X"04fb3d0d",
X"800b83e7",
X"bc349080",
X"80528684",
X"808051ff",
X"b3ea3f83",
X"e0800881",
X"973889dc",
X"3f80fc80",
X"51ffb8a9",
X"3f83e080",
X"08559c80",
X"0a5480c0",
X"805380f7",
X"d45283e0",
X"800851f6",
X"ac3f83e7",
X"d8085380",
X"f7e45274",
X"51ffb2f2",
X"3f83e080",
X"088438f6",
X"ba3f83e7",
X"dc085380",
X"f7f05274",
X"51ffb2da",
X"3f83e080",
X"08b63887",
X"3dfc0554",
X"84808053",
X"86a88080",
X"5283e7dc",
X"0851ffb0",
X"e53f83e0",
X"80089338",
X"75848080",
X"2e098106",
X"8938810b",
X"83e7bc34",
X"8739800b",
X"83e7bc34",
X"83e7bc33",
X"51f1a63f",
X"8151f392",
X"3f938d3f",
X"8151f38a",
X"3f8151fd",
X"a13ffa39",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"0280f7fc",
X"0b83e38c",
X"0c80f880",
X"0b83e384",
X"0c80f884",
X"0b83e394",
X"0c83e08c",
X"08fc050c",
X"800b83e7",
X"c40b83e0",
X"8c08f805",
X"0c83e08c",
X"08f4050c",
X"ffb0f53f",
X"83e08008",
X"8605fc06",
X"83e08c08",
X"f0050c02",
X"83e08c08",
X"f0050831",
X"0d833d70",
X"83e08c08",
X"f8050870",
X"840583e0",
X"8c08f805",
X"0c0c51ff",
X"adbd3f83",
X"e08c08f4",
X"05088105",
X"83e08c08",
X"f4050c83",
X"e08c08f4",
X"0508872e",
X"098106ff",
X"ab388694",
X"808051ea",
X"d33fff0b",
X"83e7c00c",
X"800b83e7",
X"e40c84d8",
X"c00b83e7",
X"e00c8151",
X"edfd3f81",
X"51eea23f",
X"8051ee9d",
X"3f8151ee",
X"c33f8251",
X"eeeb3f80",
X"51ef933f",
X"8051efbd",
X"3f80d0af",
X"528051df",
X"b73ffce1",
X"3f83e08c",
X"08fc0508",
X"0d800b83",
X"e0800c87",
X"3d0d83e0",
X"8c0c0480",
X"3d0d81ff",
X"51800b83",
X"e7f41234",
X"ff115170",
X"f438823d",
X"0d04ff3d",
X"0d737033",
X"53518111",
X"33713471",
X"81123483",
X"3d0d04fb",
X"3d0d7779",
X"56568070",
X"71555552",
X"717525ac",
X"38721670",
X"33701470",
X"81ff0655",
X"51515171",
X"74278938",
X"81127081",
X"ff065351",
X"71811470",
X"83ffff06",
X"55525474",
X"7324d638",
X"7183e080",
X"0c873d0d",
X"04fb3d0d",
X"7756d781",
X"3f83e080",
X"08802ef6",
X"3883ea90",
X"08860570",
X"81ff0652",
X"53d5833f",
X"810b9088",
X"d4349088",
X"d4337081",
X"ff065153",
X"728b38fa",
X"813f8351",
X"eef13fea",
X"39805574",
X"1675822b",
X"54549088",
X"c0133374",
X"34811555",
X"74852e09",
X"8106e838",
X"810b9088",
X"d4347533",
X"83e7f434",
X"81163383",
X"e7f53482",
X"163383e7",
X"f6348316",
X"3383e7f7",
X"34845283",
X"e7f451fe",
X"ba3f83e0",
X"800881ff",
X"06841733",
X"57537276",
X"2e098106",
X"8c38d5aa",
X"3f83e080",
X"08802e9c",
X"3883ea90",
X"08a82e09",
X"81068b38",
X"83eaa808",
X"83ea900c",
X"8739a80b",
X"83ea900c",
X"80e451ed",
X"ea3f873d",
X"0d04f43d",
X"0d7e6059",
X"55805d80",
X"75822b71",
X"83ea9412",
X"0c83eaac",
X"175b5b57",
X"76793477",
X"772e83b7",
X"38765277",
X"51ffac86",
X"3f8e3dfc",
X"05549053",
X"83e9fc52",
X"7751ffab",
X"c13f7c56",
X"75902e09",
X"81068393",
X"3883e9fc",
X"51fd933f",
X"83e9fe51",
X"fd8c3f83",
X"ea8051fd",
X"853f7683",
X"ea8c0c77",
X"51ffa98d",
X"3f80f5fc",
X"5283e080",
X"0851cba6",
X"3f83e080",
X"08812e09",
X"810680d4",
X"387683ea",
X"a40c820b",
X"83e9fc34",
X"ff960b83",
X"e9fd3477",
X"51ffabd3",
X"3f83e080",
X"085583e0",
X"80087725",
X"883883e0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83e9fe34",
X"7483e9ff",
X"347683ea",
X"8034ff80",
X"0b83ea81",
X"34819039",
X"83e9fc33",
X"83e9fd33",
X"71882b07",
X"565b7483",
X"ffff2e09",
X"810680e8",
X"38fe800b",
X"83eaa40c",
X"810b83ea",
X"8c0cff0b",
X"83e9fc34",
X"ff0b83e9",
X"fd347751",
X"ffaae03f",
X"83e08008",
X"83eab00c",
X"83e08008",
X"5583e080",
X"08802588",
X"3883e080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"e9fe3474",
X"83e9ff34",
X"7683ea80",
X"34ff800b",
X"83ea8134",
X"810b83ea",
X"8b34a539",
X"7485962e",
X"09810680",
X"fe387583",
X"eaa40c77",
X"51ffaa94",
X"3f83ea8b",
X"3383e080",
X"08075574",
X"83ea8b34",
X"83ea8b33",
X"81065574",
X"802e8338",
X"845783ea",
X"803383ea",
X"81337188",
X"2b07565c",
X"7481802e",
X"098106a1",
X"3883e9fe",
X"3383e9ff",
X"3371882b",
X"07565bad",
X"80752787",
X"38768207",
X"579c3976",
X"81075796",
X"39748280",
X"2e098106",
X"87387683",
X"07578739",
X"7481ff26",
X"8a387783",
X"ea941b0c",
X"7679348e",
X"3d0d0480",
X"3d0d7284",
X"2983ea94",
X"05700883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"7083e7ec",
X"0c708429",
X"80fbc005",
X"700883ea",
X"a80c5151",
X"823d0d04",
X"fe3d0d81",
X"51de3f80",
X"0b83e9f8",
X"0c800b83",
X"e9f40cff",
X"0b83e7f0",
X"0ca80b83",
X"ea900cae",
X"51cfab3f",
X"800b83ea",
X"94545280",
X"73708405",
X"550c8112",
X"5271842e",
X"098106ef",
X"38843d0d",
X"04fe3d0d",
X"74028405",
X"96052253",
X"5371802e",
X"96387270",
X"81055433",
X"51cfb63f",
X"ff127083",
X"ffff0651",
X"52e73984",
X"3d0d04fe",
X"3d0d0292",
X"05225382",
X"ac51e8df",
X"3f80c351",
X"cf933f81",
X"9651e8d3",
X"3f725283",
X"e7f451ff",
X"b43f7252",
X"83e7f451",
X"f8d13f83",
X"e0800881",
X"ff0651ce",
X"f03f843d",
X"0d04ffb1",
X"3d0d80d1",
X"3df80551",
X"f8fb3f83",
X"e9f80881",
X"0583e9f8",
X"0c80cf3d",
X"33cf1170",
X"81ff0651",
X"56567483",
X"2688e638",
X"758f06ff",
X"05567583",
X"e7f0082e",
X"9b387583",
X"26963875",
X"83e7f00c",
X"75842983",
X"ea940570",
X"08535575",
X"51f9fb3f",
X"80762488",
X"c2387584",
X"2983ea94",
X"05557408",
X"802e88b3",
X"3883e7f0",
X"08842983",
X"ea940570",
X"08028805",
X"82b90533",
X"525b5574",
X"80d22e84",
X"b0387480",
X"d2249038",
X"74bf2e9c",
X"387480d0",
X"2e81d538",
X"87f23974",
X"80d32e80",
X"d3387480",
X"d72e81c4",
X"3887e139",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"055656cd",
X"ec3f80c1",
X"51cda63f",
X"f6cd3f83",
X"eaab3383",
X"e7f43481",
X"5283e7f4",
X"51cec73f",
X"8151fde7",
X"3f748b38",
X"83eaa808",
X"83ea900c",
X"8739a80b",
X"83ea900c",
X"cdb73f80",
X"c151ccf1",
X"3ff6983f",
X"900b83ea",
X"8b338106",
X"56567480",
X"2e833898",
X"5683ea80",
X"3383ea81",
X"3371882b",
X"07565974",
X"81802e09",
X"81069c38",
X"83e9fe33",
X"83e9ff33",
X"71882b07",
X"5657ad80",
X"75278c38",
X"75818007",
X"56853975",
X"a0075675",
X"83e7f434",
X"ff0b83e7",
X"f534e00b",
X"83e7f634",
X"800b83e7",
X"f7348452",
X"83e7f451",
X"cdbc3f84",
X"51869b39",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"055659cc",
X"ac3f7951",
X"ffa4c13f",
X"83e08008",
X"802e8a38",
X"80ce51cb",
X"d83f85f1",
X"3980c151",
X"cbcf3fcc",
X"c43fcaf9",
X"3f83eaa4",
X"08588375",
X"259b3883",
X"ea803383",
X"ea813371",
X"882b07fc",
X"1771297a",
X"05838005",
X"5a51578d",
X"39748180",
X"2918ff80",
X"05588180",
X"57805676",
X"762e9238",
X"cbab3f83",
X"e0800883",
X"e7f41734",
X"811656eb",
X"39cb9a3f",
X"83e08008",
X"81ff0677",
X"5383e7f4",
X"5256f4c3",
X"3f83e080",
X"0881ff06",
X"5575752e",
X"09810681",
X"95389451",
X"e49d3fcb",
X"943f80c1",
X"51cace3f",
X"cbc33f77",
X"527951ff",
X"a2d43f80",
X"5e80d13d",
X"fdf40554",
X"765383e7",
X"f4527951",
X"ffa0e13f",
X"0282b905",
X"33558159",
X"7480d72e",
X"09810680",
X"c5387752",
X"7951ffa2",
X"a53f80d1",
X"3dfdf005",
X"5476538f",
X"3d70537a",
X"5258ffa1",
X"dd3f8056",
X"76762ea2",
X"38751883",
X"e7f41733",
X"71337072",
X"32703070",
X"80257030",
X"7f06811d",
X"5d5f5151",
X"51525b55",
X"db3982ac",
X"51e3983f",
X"78802e86",
X"3880c351",
X"843980ce",
X"51c9c23f",
X"cab73fc8",
X"ec3f83d8",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055955",
X"80705d59",
X"80e451e2",
X"e23fc9d9",
X"3f80c151",
X"c9933f83",
X"ea8c0879",
X"2e82d638",
X"83eab008",
X"80fc0555",
X"80fd5274",
X"5185c13f",
X"83e08008",
X"5b778224",
X"b238ff18",
X"70872b83",
X"ffff8006",
X"80fa8c05",
X"83e7f459",
X"57558180",
X"55757081",
X"05573377",
X"70810559",
X"34ff1570",
X"81ff0651",
X"5574ea38",
X"82853977",
X"82e82e81",
X"a3387782",
X"e92e0981",
X"0681aa38",
X"78587787",
X"32703070",
X"72078025",
X"7a8a3270",
X"30707207",
X"80257307",
X"53545a51",
X"57557580",
X"2e973878",
X"78269238",
X"a00b83e7",
X"f41a3481",
X"197081ff",
X"065a55eb",
X"39811870",
X"81ff0659",
X"558a7827",
X"ffbc388f",
X"5883e7ef",
X"183383e7",
X"f41934ff",
X"187081ff",
X"06595577",
X"8426ea38",
X"9058800b",
X"83e7f419",
X"34811870",
X"81ff0670",
X"982b5259",
X"55748025",
X"e93880c6",
X"557a858f",
X"24843880",
X"c2557483",
X"e7f43480",
X"f10b83e7",
X"f734810b",
X"83e7f834",
X"7a83e7f5",
X"347a882c",
X"557483e7",
X"f63480cb",
X"3982f078",
X"2580c438",
X"7780fd29",
X"fd97d305",
X"527951ff",
X"9f803f80",
X"d13dfdec",
X"055480fd",
X"5383e7f4",
X"527951ff",
X"9eb83f7b",
X"81195956",
X"7580fc24",
X"83387858",
X"77882c55",
X"7483e8f1",
X"347783e8",
X"f2347583",
X"e8f33481",
X"805980cc",
X"3983eaa4",
X"08578378",
X"259b3883",
X"ea803383",
X"ea813371",
X"882b07fc",
X"1a712979",
X"05838005",
X"5951598d",
X"39778180",
X"2917ff80",
X"05578180",
X"59765279",
X"51ff9e8e",
X"3f80d13d",
X"fdec0554",
X"785383e7",
X"f4527951",
X"ff9dc73f",
X"7851f6bf",
X"3fc6da3f",
X"c58f3f8b",
X"3983e9f4",
X"08810583",
X"e9f40c80",
X"d13d0d04",
X"f6e03ffc",
X"39fc3d0d",
X"76787184",
X"2983ea94",
X"05700851",
X"53535370",
X"9e3880ce",
X"723480cf",
X"0b811334",
X"80ce0b82",
X"133480c5",
X"0b831334",
X"70841334",
X"80e73983",
X"eaac1333",
X"5480d272",
X"3473822a",
X"70810651",
X"5180cf53",
X"70843880",
X"d7537281",
X"1334a00b",
X"82133473",
X"83065170",
X"812e9e38",
X"70812488",
X"3870802e",
X"8f389f39",
X"70822e92",
X"3870832e",
X"92389339",
X"80d8558e",
X"3980d355",
X"893980cd",
X"55843980",
X"c4557483",
X"133480c4",
X"0b841334",
X"800b8513",
X"34863d0d",
X"0483e7ec",
X"0883e080",
X"0c04803d",
X"0d83e7ec",
X"08842980",
X"fbe00570",
X"0883e080",
X"0c51823d",
X"0d04fc3d",
X"0d767853",
X"54815380",
X"55873971",
X"10731054",
X"52737226",
X"5172802e",
X"a7387080",
X"2e863871",
X"8025e838",
X"72802e98",
X"38717426",
X"89387372",
X"31757407",
X"56547281",
X"2a72812a",
X"5353e539",
X"73517883",
X"38745170",
X"83e0800c",
X"863d0d04",
X"fe3d0d80",
X"53755274",
X"51ffa33f",
X"843d0d04",
X"fe3d0d81",
X"53755274",
X"51ff933f",
X"843d0d04",
X"fb3d0d77",
X"79555580",
X"56747625",
X"86387430",
X"55815673",
X"80258838",
X"73307681",
X"32575480",
X"53735274",
X"51fee73f",
X"83e08008",
X"5475802e",
X"873883e0",
X"80083054",
X"7383e080",
X"0c873d0d",
X"04fa3d0d",
X"787a5755",
X"80577477",
X"25863874",
X"30558157",
X"759f2c54",
X"81537574",
X"32743152",
X"7451feaa",
X"3f83e080",
X"08547680",
X"2e873883",
X"e0800830",
X"547383e0",
X"800c883d",
X"0d04fd3d",
X"0d755480",
X"740c800b",
X"84150c80",
X"0b88150c",
X"800b8c15",
X"0c87a680",
X"337081ff",
X"065151db",
X"a93f7081",
X"2a813271",
X"81327181",
X"06718106",
X"3184170c",
X"53537083",
X"2a813271",
X"822a8132",
X"71810671",
X"81063176",
X"0c525287",
X"a0903370",
X"09810688",
X"160c5183",
X"e0800880",
X"2e80c238",
X"83e08008",
X"812a7081",
X"0683e080",
X"08810631",
X"84160c51",
X"83e08008",
X"832a83e0",
X"8008822a",
X"71810671",
X"81063176",
X"0c525283",
X"e0800884",
X"2a810688",
X"150c83e0",
X"8008852a",
X"81068c15",
X"0c853d0d",
X"04fe3d0d",
X"74765452",
X"7151fece",
X"3f72812e",
X"a2388173",
X"268d3872",
X"822ea838",
X"72832e9c",
X"38e63971",
X"08e23884",
X"1208dd38",
X"881208d8",
X"38a53988",
X"1208812e",
X"9e389139",
X"88120881",
X"2e953871",
X"08913884",
X"12088c38",
X"8c120881",
X"2e098106",
X"ffb23884",
X"3d0d0400",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002b19",
X"00002b5a",
X"00002b7c",
X"00002b9e",
X"00002bc4",
X"00002bc4",
X"00002bc4",
X"00002bc4",
X"00002c35",
X"00002c86",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"43505520",
X"54757262",
X"6f3a2564",
X"78000000",
X"44726976",
X"65205475",
X"72626f3a",
X"25730000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"66726565",
X"7a65722e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"5374616e",
X"64617264",
X"00000000",
X"46617374",
X"28362900",
X"46617374",
X"28352900",
X"46617374",
X"28342900",
X"46617374",
X"28332900",
X"46617374",
X"28322900",
X"46617374",
X"28312900",
X"46617374",
X"28302900",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00003b28",
X"00003b2c",
X"00003b34",
X"00003b40",
X"00003b4c",
X"00003b58",
X"00003b64",
X"00003b68",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00000028",
X"00000006",
X"00000005",
X"00000004",
X"00000003",
X"00000002",
X"00000001",
X"00000000",
X"00003c08",
X"00003c14",
X"00003c1c",
X"00003c24",
X"00003c2c",
X"00003c34",
X"00003c3c",
X"00003c44",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
