
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f8",
X"c4738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80fb",
X"980c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f2",
X"f22d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580f186",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"96e80480",
X"3d0d80fc",
X"dc087008",
X"810683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d80fc",
X"dc087008",
X"70fe0676",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80fcdc08",
X"70087081",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80fcdc08",
X"700870fd",
X"06761007",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"fcdc0870",
X"0870822c",
X"bf0683e0",
X"800c5151",
X"823d0d04",
X"ff3d0d80",
X"fcdc0870",
X"0870fe83",
X"0676822b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80fcdc08",
X"70087088",
X"2c870683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80fcdc08",
X"700870f1",
X"ff067688",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d80fcdc",
X"08700870",
X"8b2cbf06",
X"83e0800c",
X"5151823d",
X"0d04ff3d",
X"0d80fcdc",
X"08700870",
X"f88fff06",
X"768b2b07",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"fcec0870",
X"0870882c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fcec0870",
X"0870892c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fcec0870",
X"08708a2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fcec0870",
X"08708b2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"fd3d0d75",
X"81e62987",
X"2a80fccc",
X"0854730c",
X"853d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d848080",
X"53805288",
X"800a51ff",
X"b33f8180",
X"80538052",
X"82800a51",
X"c63f843d",
X"0d04803d",
X"0d8151fc",
X"ce3f7280",
X"2e8338d2",
X"3f8151fc",
X"f03f8051",
X"fceb3f80",
X"51fcb83f",
X"823d0d04",
X"fd3d0d75",
X"52805480",
X"ff722588",
X"38810bff",
X"80135354",
X"ffbf1251",
X"70992686",
X"38e01252",
X"9e39ff9f",
X"12519971",
X"279538d0",
X"12e01370",
X"54545189",
X"71278838",
X"8f732783",
X"38805273",
X"802e8538",
X"81801252",
X"7181ff06",
X"83e0800c",
X"853d0d04",
X"803d0d86",
X"b8c05180",
X"71708105",
X"53347086",
X"c0c02e09",
X"8106f038",
X"823d0d04",
X"fe3d0d02",
X"97053351",
X"ff863f83",
X"e0800881",
X"ff0683e0",
X"9c085452",
X"8073249b",
X"3883e0b8",
X"08137283",
X"e0bc0807",
X"53537173",
X"3483e09c",
X"08810583",
X"e09c0c84",
X"3d0d04fa",
X"3d0d8280",
X"0a1b5580",
X"57883dfc",
X"05547953",
X"74527851",
X"b4f73f88",
X"3d0d04fe",
X"3d0d83e0",
X"b0085274",
X"51bbd93f",
X"83e08008",
X"8c387653",
X"755283e0",
X"b00851c7",
X"3f843d0d",
X"04fe3d0d",
X"83e0b008",
X"53755274",
X"51b6993f",
X"83e08008",
X"8d387753",
X"765283e0",
X"b00851ff",
X"a23f843d",
X"0d04fe3d",
X"0d83e0b4",
X"0851b58d",
X"3f83e080",
X"08818080",
X"2e098106",
X"8738b180",
X"80539a39",
X"83e0b408",
X"51b4f23f",
X"83e08008",
X"80d0802e",
X"09810692",
X"38b1b080",
X"5383e080",
X"085283e0",
X"b40851fe",
X"da3f843d",
X"0d04803d",
X"0dface3f",
X"83e08008",
X"842980fb",
X"a0057008",
X"83e0800c",
X"51823d0d",
X"04ee3d0d",
X"80438042",
X"80418070",
X"5a5bfdd4",
X"3f800b83",
X"e09c0c80",
X"0b83e0bc",
X"0c0b0b80",
X"f9e051af",
X"dd3f8180",
X"0b83e0bc",
X"0c0b0b80",
X"f9e451af",
X"cd3f80d0",
X"0b83e09c",
X"0c783070",
X"7a078025",
X"70872b83",
X"e0bc0c51",
X"55f9b93f",
X"83e08008",
X"520b0b80",
X"f9ec51af",
X"a53f80f8",
X"0b83e09c",
X"0c788132",
X"70307072",
X"07802570",
X"872b83e0",
X"bc0c5156",
X"56feeb3f",
X"83e08008",
X"520b0b80",
X"f9f851ae",
X"f93f81a0",
X"0b83e09c",
X"0c788232",
X"70307072",
X"07802570",
X"872b83e0",
X"bc0c5156",
X"83e0b408",
X"5256b094",
X"3f83e080",
X"08520b0b",
X"80fa8051",
X"aec83f81",
X"f00b83e0",
X"9c0c810b",
X"83e0a05b",
X"5883e09c",
X"0882197a",
X"32703070",
X"72078025",
X"70872b83",
X"e0bc0c51",
X"578e3d70",
X"55ff1b54",
X"575757a4",
X"a63f7970",
X"84055b08",
X"51afc93f",
X"745483e0",
X"80085377",
X"520b0b80",
X"fa8851ad",
X"f93fa817",
X"83e09c0c",
X"81185877",
X"852e0981",
X"06ffae38",
X"83900b83",
X"e09c0c78",
X"87327030",
X"70720780",
X"2570872b",
X"83e0bc0c",
X"51560b0b",
X"80fa9852",
X"56adc33f",
X"83e00b83",
X"e09c0c78",
X"88327030",
X"70720780",
X"2570872b",
X"83e0bc0c",
X"51560b0b",
X"80faac52",
X"56ad9f3f",
X"868da051",
X"f9923f80",
X"52913d70",
X"52558ba5",
X"3f835274",
X"518b9e3f",
X"61195978",
X"80258538",
X"80599039",
X"88792585",
X"38885987",
X"39788826",
X"82ae3878",
X"822b5580",
X"f8d41508",
X"04f6e53f",
X"83e08008",
X"61575575",
X"812e0981",
X"06893883",
X"e0800810",
X"55903975",
X"ff2e0981",
X"06883883",
X"e0800881",
X"2c559075",
X"25853890",
X"55883974",
X"80248338",
X"81557451",
X"f6c23f81",
X"e339f6d5",
X"3f83e080",
X"08610555",
X"74802585",
X"38805588",
X"39877525",
X"83388755",
X"7451f6d1",
X"3f81c139",
X"60873862",
X"802e81b8",
X"38a0970b",
X"83e0d00c",
X"83e0b408",
X"518ca93f",
X"fb803f81",
X"a3396056",
X"80762598",
X"389fb60b",
X"83e0d00c",
X"83e09415",
X"70085255",
X"8c8a3f74",
X"08529139",
X"75802591",
X"3883e094",
X"150851ad",
X"853f8052",
X"fd1951b8",
X"3962802e",
X"80ea3883",
X"e0941570",
X"0883e0a0",
X"08720c83",
X"e0a00cfd",
X"1a705351",
X"5596dc3f",
X"83e08008",
X"56805196",
X"d23f83e0",
X"80085274",
X"5192f13f",
X"75528051",
X"92ea3fb4",
X"3962802e",
X"af38a097",
X"0b83e0d0",
X"0c83e0b0",
X"08518ba0",
X"3f83e0b0",
X"0851ac94",
X"3f9c800a",
X"5380c080",
X"5283e080",
X"0851f99b",
X"3f81558c",
X"39628738",
X"7a802efa",
X"c5388055",
X"7483e080",
X"0c943d0d",
X"04fe3d0d",
X"f5c23f83",
X"e0800880",
X"2e863880",
X"5180f639",
X"f5ca3f83",
X"e0800880",
X"ea38f5f0",
X"3f83e080",
X"08802eaa",
X"388151f3",
X"c23f839b",
X"3f800b83",
X"e09c0cf9",
X"f43f83e0",
X"800853ff",
X"0b83e09c",
X"0c85ee3f",
X"72bd3872",
X"51f3a03f",
X"bb39f5a4",
X"3f83e080",
X"08802eb0",
X"388151f3",
X"8e3f82e7",
X"3f9fb60b",
X"83e0d00c",
X"83e0a008",
X"5189fd3f",
X"ff0b83e0",
X"9c0c85b9",
X"3f83e0a0",
X"08528051",
X"919e3f81",
X"51f68f3f",
X"843d0d04",
X"83e08c08",
X"0283e08c",
X"0cfa3d0d",
X"800b83e0",
X"a00b83e0",
X"8c08fc05",
X"0c83e08c",
X"08f8050c",
X"add03f83",
X"e0800886",
X"05fc0683",
X"e08c08f4",
X"050c0283",
X"e08c08f4",
X"0508310d",
X"853d7083",
X"e08c08fc",
X"05087084",
X"0583e08c",
X"08fc050c",
X"0c51aa9a",
X"3f83e08c",
X"08f80508",
X"810583e0",
X"8c08f805",
X"0c83e08c",
X"08f80508",
X"862e0981",
X"06ffad38",
X"84a88080",
X"5181aa3f",
X"ff0b83e0",
X"9c0c800b",
X"83e0bc0c",
X"86b8c00b",
X"83e0b80c",
X"8151f1cb",
X"3f8151f1",
X"f43f8051",
X"f1ef3f81",
X"51f2993f",
X"8151f2f6",
X"3f8251f2",
X"c03f8e84",
X"528051a7",
X"de3f8480",
X"805284a4",
X"808051ad",
X"b93f83e0",
X"800880d3",
X"3893b53f",
X"80fea451",
X"b1f83f83",
X"e0800883",
X"e0b40854",
X"0b0b80fa",
X"b45383e0",
X"80085283",
X"e08c08f4",
X"050caccc",
X"3f83e080",
X"088438f6",
X"c13fb080",
X"805480c0",
X"80530b0b",
X"80fac052",
X"83e08c08",
X"f4050851",
X"f6833f81",
X"51f3f33f",
X"9d8d3f81",
X"51f3eb3f",
X"fccf3ffc",
X"397183e0",
X"c40c8880",
X"800b83e0",
X"c00c8480",
X"800b83e0",
X"c80c04f0",
X"3d0d80fb",
X"d4085473",
X"3383e0cc",
X"3483a080",
X"5683e0c4",
X"081683e0",
X"c0081756",
X"54743374",
X"3483e0c8",
X"08165480",
X"74348116",
X"567583a0",
X"a02e0981",
X"06db3883",
X"a4805683",
X"e0c40816",
X"83e0c008",
X"17565474",
X"33743483",
X"e0c80816",
X"54807434",
X"81165675",
X"83a4a02e",
X"098106db",
X"3883a880",
X"5683e0c4",
X"081683e0",
X"c0081756",
X"54743374",
X"3483e0c8",
X"08165480",
X"74348116",
X"567583a8",
X"902e0981",
X"06db3880",
X"fbd40854",
X"ff743480",
X"5683e0c4",
X"081683e0",
X"c8081755",
X"55733375",
X"34811656",
X"7583a080",
X"2e098106",
X"e43883b0",
X"805683e0",
X"c4081683",
X"e0c80817",
X"55557333",
X"75348116",
X"56758480",
X"802e0981",
X"06e438f2",
X"ef3f893d",
X"58a25380",
X"f8f85277",
X"5180dc9f",
X"3f80578c",
X"805683e0",
X"c8081677",
X"19555573",
X"33753481",
X"16811858",
X"5676a22e",
X"098106e6",
X"3880fbf8",
X"08548674",
X"3480fbfc",
X"08548074",
X"3480fbf4",
X"08548074",
X"3480fbe4",
X"0854af74",
X"3480fbf0",
X"0854bf74",
X"3480fbec",
X"08548074",
X"3480fbe8",
X"08549f74",
X"3480fbe0",
X"08548074",
X"3480fbcc",
X"0854e074",
X"3480fbc4",
X"08547674",
X"3480fbc0",
X"08548374",
X"3480fbc8",
X"08548274",
X"34923d0d",
X"04fe3d0d",
X"805383e0",
X"c8081383",
X"e0c40814",
X"52527033",
X"72348113",
X"537283a0",
X"802e0981",
X"06e43883",
X"b0805383",
X"e0c80813",
X"83e0c408",
X"14525270",
X"33723481",
X"13537284",
X"80802e09",
X"8106e438",
X"83a08053",
X"83e0c808",
X"1383e0c4",
X"08145252",
X"70337234",
X"81135372",
X"83a0a02e",
X"098106e4",
X"3883a480",
X"5383e0c8",
X"081383e0",
X"c4081452",
X"52703372",
X"34811353",
X"7283a4a0",
X"2e098106",
X"e43883a8",
X"805383e0",
X"c8081383",
X"e0c40814",
X"52527033",
X"72348113",
X"537283a8",
X"902e0981",
X"06e43880",
X"fbd40851",
X"83e0cc33",
X"7134843d",
X"0d04fd3d",
X"0d755480",
X"740c800b",
X"84150c80",
X"0b88150c",
X"80fbd808",
X"70337081",
X"ff067081",
X"2a813271",
X"81327181",
X"06718106",
X"31841a0c",
X"56567083",
X"2a813271",
X"822a8132",
X"71810671",
X"81063179",
X"0c525551",
X"515180fb",
X"d0087033",
X"70098106",
X"88170c51",
X"51853d0d",
X"04fe3d0d",
X"74765452",
X"7151ff9a",
X"3f72812e",
X"a2388173",
X"268d3872",
X"822eab38",
X"72832e9f",
X"38e63971",
X"08e23884",
X"1208dd38",
X"881208d8",
X"38a03988",
X"1208812e",
X"098106cc",
X"38943988",
X"1208812e",
X"8d387108",
X"89388412",
X"08802eff",
X"b738843d",
X"0d04fc3d",
X"0d767052",
X"5580c6f6",
X"3f83e080",
X"0815ff05",
X"5473752e",
X"8e387333",
X"5372ae2e",
X"8638ff14",
X"54ef3977",
X"52811451",
X"80c68d3f",
X"83e08008",
X"307083e0",
X"80080780",
X"2583e080",
X"0c53863d",
X"0d04fc3d",
X"0d767052",
X"55abe13f",
X"83e08008",
X"54815383",
X"e0800880",
X"c1387451",
X"aba43f83",
X"e0800880",
X"fadc5383",
X"e0800852",
X"53ff8f3f",
X"83e08008",
X"a13880fa",
X"e0527251",
X"ff803f83",
X"e0800892",
X"3880fae4",
X"527251fe",
X"f13f83e0",
X"8008802e",
X"83388154",
X"73537283",
X"e0800c86",
X"3d0d04fd",
X"3d0d7570",
X"5254ab80",
X"3f815383",
X"e0800897",
X"387351aa",
X"c93f80fa",
X"e85283e0",
X"800851fe",
X"b93f83e0",
X"80085372",
X"83e0800c",
X"853d0d04",
X"e03d0da3",
X"3d087052",
X"5ea0f13f",
X"83e08008",
X"33943d56",
X"54739438",
X"80feb452",
X"745184b3",
X"397d5278",
X"51a3f33f",
X"84be397d",
X"51a0d93f",
X"83e08008",
X"527451a0",
X"893f83e0",
X"d0085293",
X"3d70525d",
X"a6e33f83",
X"e0800859",
X"800b83e0",
X"8008555b",
X"83e08008",
X"7b2e9438",
X"811b7452",
X"5ba9e43f",
X"83e08008",
X"5483e080",
X"08ee3880",
X"5aff7a43",
X"7a427a41",
X"5f790970",
X"9f2c7b06",
X"5b547a7a",
X"248438ff",
X"1b5af61a",
X"7009709f",
X"2c72067b",
X"ff125a5a",
X"52555580",
X"75259538",
X"7651a9a3",
X"3f83e080",
X"0876ff18",
X"58555773",
X"8024ed38",
X"747f2e86",
X"38ebe53f",
X"745f78ff",
X"1b70585d",
X"58807a25",
X"95387751",
X"a8f93f83",
X"e0800876",
X"ff185855",
X"58738024",
X"ed38800b",
X"83e09c0c",
X"800b83e0",
X"bc0c80fa",
X"ec519dce",
X"3f81800b",
X"83e0bc0c",
X"80faf451",
X"9dc03fa8",
X"0b83e09c",
X"0c76802e",
X"80e43883",
X"e09c0877",
X"79327030",
X"70720780",
X"2570872b",
X"83e0bc0c",
X"51567853",
X"5656a8b0",
X"3f83e080",
X"08802e88",
X"3880fafc",
X"519d873f",
X"7651a7f2",
X"3f83e080",
X"085280fa",
X"94519cf6",
X"3f7651a7",
X"fa3f83e0",
X"800883e0",
X"9c085557",
X"75742586",
X"38a81656",
X"f7397583",
X"e09c0c86",
X"f07624ff",
X"98388798",
X"0b83e09c",
X"0c77802e",
X"b1387751",
X"a7b03f83",
X"e0800878",
X"5255a7d0",
X"3f80fb84",
X"5483e080",
X"088d3887",
X"39807634",
X"fda03980",
X"fb805474",
X"53735280",
X"fad0519c",
X"953f8054",
X"80fb8c51",
X"9c8c3f81",
X"145473a8",
X"2e098106",
X"ef38868d",
X"a051e7f4",
X"3f805290",
X"3d705254",
X"fa873f83",
X"527351fa",
X"803f6180",
X"2e80ff38",
X"7b5473ff",
X"2e963878",
X"802e8180",
X"387851a6",
X"da3f83e0",
X"8008ff15",
X"5559e739",
X"78802e80",
X"eb387851",
X"a6d63f83",
X"e0800880",
X"2efc9638",
X"7851a69e",
X"3f83e080",
X"085280fa",
X"d851bfcb",
X"3f83e080",
X"08a5387c",
X"5180c182",
X"3f83e080",
X"085574ff",
X"16565480",
X"7425fc82",
X"38741d70",
X"33555673",
X"af2efed1",
X"38e83978",
X"51a5dd3f",
X"83e08008",
X"527c5180",
X"c0b83ffb",
X"e1397f88",
X"29601005",
X"7a056105",
X"5afc9239",
X"a23d0d04",
X"803d0d81",
X"ff51800b",
X"83e0dc12",
X"34ff1151",
X"70f43882",
X"3d0d04ff",
X"3d0d7370",
X"33535181",
X"11337134",
X"71811234",
X"833d0d04",
X"fb3d0d77",
X"79565680",
X"70715555",
X"52717525",
X"ac387216",
X"70337014",
X"7081ff06",
X"55515151",
X"71742789",
X"38811270",
X"81ff0653",
X"51718114",
X"7083ffff",
X"06555254",
X"747324d6",
X"387183e0",
X"800c873d",
X"0d04fd3d",
X"0d755494",
X"8f3f83e0",
X"8008802e",
X"f63883e2",
X"f8088605",
X"7081ff06",
X"525391e8",
X"3f8439ef",
X"903f93f0",
X"3f83e080",
X"08812ef3",
X"3892cb3f",
X"83e08008",
X"743492c2",
X"3f83e080",
X"08811534",
X"92b83f83",
X"e0800882",
X"153492ae",
X"3f83e080",
X"08831534",
X"92a43f83",
X"e0800884",
X"15348439",
X"eecf3f93",
X"af3f83e0",
X"8008802e",
X"f3387333",
X"83e0dc34",
X"81143383",
X"e0dd3482",
X"143383e0",
X"de348314",
X"3383e0df",
X"34845283",
X"e0dc51fe",
X"a73f83e0",
X"800881ff",
X"06841533",
X"55537274",
X"2e098106",
X"8c3892a0",
X"3f83e080",
X"08802e9a",
X"3883e2f8",
X"08a82e09",
X"81068938",
X"860b83e2",
X"f80c8739",
X"a80b83e2",
X"f80c80e4",
X"51e4893f",
X"853d0d04",
X"f43d0d7e",
X"60595580",
X"5d807582",
X"2b7183e2",
X"fc120c83",
X"e390175b",
X"5b577679",
X"3477772e",
X"83b13876",
X"5277519b",
X"e13f8e3d",
X"fc055490",
X"5383e2e4",
X"5277519b",
X"983f7c56",
X"75902e09",
X"8106838f",
X"3883e2e4",
X"51fd843f",
X"83e2e651",
X"fcfd3f83",
X"e2e851fc",
X"f63f7683",
X"e2f40c77",
X"5198e53f",
X"80fae052",
X"83e08008",
X"51f6873f",
X"83e08008",
X"812e0981",
X"0680d338",
X"7683e38c",
X"0c820b83",
X"e2e434ff",
X"960b83e2",
X"e5347751",
X"9bab3f83",
X"e0800855",
X"83e08008",
X"77258838",
X"83e08008",
X"8f055574",
X"842c7083",
X"ffff0670",
X"882a5851",
X"557583e2",
X"e6347483",
X"e2e73476",
X"83e2e834",
X"ff800b83",
X"e2e93481",
X"8f3983e2",
X"e43383e2",
X"e5337188",
X"2b07565b",
X"7483ffff",
X"2e098106",
X"80e738fe",
X"800b83e3",
X"8c0c810b",
X"83e2f40c",
X"ff0b83e2",
X"e434ff0b",
X"83e2e534",
X"77519ab9",
X"3f83e080",
X"0883e394",
X"0c83e080",
X"085583e0",
X"80088025",
X"883883e0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83e2e634",
X"7483e2e7",
X"347683e2",
X"e834ff80",
X"0b83e2e9",
X"34810b83",
X"e2f334a4",
X"39748596",
X"2e098106",
X"80fd3875",
X"83e38c0c",
X"775199ee",
X"3f83e2f3",
X"3383e080",
X"08075574",
X"83e2f334",
X"83e2f333",
X"81065574",
X"802e8338",
X"845783e2",
X"e83383e2",
X"e9337188",
X"2b07565c",
X"7481802e",
X"098106a1",
X"3883e2e6",
X"3383e2e7",
X"3371882b",
X"07565bad",
X"80752787",
X"38768207",
X"579c3976",
X"81075796",
X"39748280",
X"2e098106",
X"87387683",
X"07578739",
X"7481ff26",
X"8a387783",
X"e2fc1b0c",
X"7679348e",
X"3d0d0480",
X"3d0d7284",
X"2983e2fc",
X"05700883",
X"e0800c51",
X"823d0d04",
X"fe3d0d80",
X"0b83e2e0",
X"0c800b83",
X"e2dc0cff",
X"0b83e0d8",
X"0ca80b83",
X"e2f80cae",
X"518ca53f",
X"800b83e2",
X"fc545280",
X"73708405",
X"550c8112",
X"5271842e",
X"098106ef",
X"38843d0d",
X"04fe3d0d",
X"74028405",
X"96052253",
X"5371802e",
X"96387270",
X"81055433",
X"518cc43f",
X"ff127083",
X"ffff0651",
X"52e73984",
X"3d0d04fe",
X"3d0d0292",
X"05225382",
X"ac51dfa4",
X"3f80c351",
X"8ca13f81",
X"9651df98",
X"3f725283",
X"e0dc51ff",
X"b43f7252",
X"83e0dc51",
X"f8e63f83",
X"e0800881",
X"ff06518b",
X"fe3f843d",
X"0d04ffb1",
X"3d0d80d1",
X"3df80551",
X"f9903f83",
X"e2e00881",
X"0583e2e0",
X"0c80cf3d",
X"33cf1170",
X"81ff0651",
X"56567483",
X"2688cd38",
X"758f06ff",
X"05567583",
X"e0d8082e",
X"9b387583",
X"26963875",
X"83e0d80c",
X"75842983",
X"e2fc0570",
X"08535575",
X"51faa13f",
X"80762488",
X"a9387584",
X"2983e2fc",
X"05557408",
X"802e889a",
X"3883e0d8",
X"08842983",
X"e2fc0570",
X"08028805",
X"82b90533",
X"525b5574",
X"80d22e84",
X"9a387480",
X"d2249038",
X"74bf2e9c",
X"387480d0",
X"2e81d138",
X"87d93974",
X"80d32e80",
X"cf387480",
X"d72e81c0",
X"3887c839",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"0556568b",
X"803f80c1",
X"518ab43f",
X"f6e23f86",
X"0b83e0dc",
X"34815283",
X"e0dc518b",
X"ef3f8151",
X"fde93f74",
X"8938860b",
X"83e2f80c",
X"8739a80b",
X"83e2f80c",
X"8acf3f80",
X"c1518a83",
X"3ff6b13f",
X"900b83e2",
X"f3338106",
X"56567480",
X"2e833898",
X"5683e2e8",
X"3383e2e9",
X"3371882b",
X"07565974",
X"81802e09",
X"81069c38",
X"83e2e633",
X"83e2e733",
X"71882b07",
X"5657ad80",
X"75278c38",
X"75818007",
X"56853975",
X"a0075675",
X"83e0dc34",
X"ff0b83e0",
X"dd34e00b",
X"83e0de34",
X"800b83e0",
X"df348452",
X"83e0dc51",
X"8ae63f84",
X"51868639",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"05565989",
X"c43f7951",
X"94c03f83",
X"e0800880",
X"2e8a3880",
X"ce5188eb",
X"3f85dd39",
X"80c15188",
X"e23f89ea",
X"3f87ee3f",
X"83e38c08",
X"58837525",
X"9b3883e2",
X"e83383e2",
X"e9337188",
X"2b07fc17",
X"71297a05",
X"8380055a",
X"51578d39",
X"74818029",
X"18ff8005",
X"58818057",
X"80567676",
X"2e923888",
X"c13f83e0",
X"800883e0",
X"dc173481",
X"1656eb39",
X"88b03f83",
X"e0800881",
X"ff067753",
X"83e0dc52",
X"56f4dd3f",
X"83e08008",
X"81ff0655",
X"75752e09",
X"81068184",
X"3888b23f",
X"80c15187",
X"e63f88ee",
X"3f775279",
X"5192df3f",
X"805e80d1",
X"3dfdf405",
X"54765383",
X"e0dc5279",
X"5190e83f",
X"0282b905",
X"33558158",
X"7480d72e",
X"098106bc",
X"3880d13d",
X"fdf00554",
X"76538f3d",
X"70537a52",
X"5991ee3f",
X"80567676",
X"2ea23875",
X"1983e0dc",
X"17337133",
X"70723270",
X"30708025",
X"70307e06",
X"811d5d5e",
X"51515152",
X"5b55db39",
X"82ac51d9",
X"f33f7780",
X"2e863880",
X"c3518439",
X"80ce5186",
X"e63f87ee",
X"3f85f23f",
X"83d53902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"59558070",
X"5d598789",
X"3f80c151",
X"86bd3f83",
X"e2f40879",
X"2e82db38",
X"83e39408",
X"80fc0555",
X"80fd5274",
X"51bdc13f",
X"83e08008",
X"5b778224",
X"b238ff18",
X"70872b83",
X"ffff8006",
X"80fcf005",
X"83e0dc59",
X"57558180",
X"55757081",
X"05573377",
X"70810559",
X"34ff1570",
X"81ff0651",
X"5574ea38",
X"828a3977",
X"82e82e81",
X"aa387782",
X"e92e0981",
X"0681b138",
X"80fb8851",
X"8cd43f78",
X"58778732",
X"70307072",
X"0780257a",
X"8a327030",
X"70720780",
X"25730753",
X"545a5157",
X"5575802e",
X"97387878",
X"269238a0",
X"0b83e0dc",
X"1a348119",
X"7081ff06",
X"5a55eb39",
X"81187081",
X"ff065955",
X"8a7827ff",
X"bc388f58",
X"83e0d718",
X"3383e0dc",
X"1934ff18",
X"7081ff06",
X"59557784",
X"26ea3890",
X"58800b83",
X"e0dc1934",
X"81187081",
X"ff067098",
X"2b525955",
X"748025e9",
X"3880c655",
X"7a858f24",
X"843880c2",
X"557483e0",
X"dc3480f1",
X"0b83e0df",
X"34810b83",
X"e0e0347a",
X"83e0dd34",
X"7a882c55",
X"7483e0de",
X"3480c939",
X"82f07825",
X"80c23877",
X"80fd29fd",
X"97d30552",
X"79518f96",
X"3f80d13d",
X"fdec0554",
X"80fd5383",
X"e0dc5279",
X"518eca3f",
X"7b811959",
X"567580fc",
X"24833878",
X"5877882c",
X"557483e1",
X"d9347783",
X"e1da3475",
X"83e1db34",
X"81805980",
X"ca3983e3",
X"8c085783",
X"78259b38",
X"83e2e833",
X"83e2e933",
X"71882b07",
X"fc1a7129",
X"79058380",
X"05595159",
X"8d397781",
X"802917ff",
X"80055781",
X"80597652",
X"79518ea6",
X"3f80d13d",
X"fdec0554",
X"785383e0",
X"dc527951",
X"8ddb3f78",
X"51f6d83f",
X"84943f82",
X"983f8b39",
X"83e2dc08",
X"810583e2",
X"dc0c80d1",
X"3d0d04f6",
X"f93fdfc5",
X"3ff939fc",
X"3d0d7678",
X"71842983",
X"e2fc0570",
X"08515353",
X"53709e38",
X"80ce7234",
X"80cf0b81",
X"133480ce",
X"0b821334",
X"80c50b83",
X"13347084",
X"133480e7",
X"3983e390",
X"13335480",
X"d2723473",
X"822a7081",
X"06515180",
X"cf537084",
X"3880d753",
X"72811334",
X"a00b8213",
X"34738306",
X"5170812e",
X"9e387081",
X"24883870",
X"802e8f38",
X"9f397082",
X"2e923870",
X"832e9238",
X"933980d8",
X"558e3980",
X"d3558939",
X"80cd5584",
X"3980c455",
X"74831334",
X"80c40b84",
X"1334800b",
X"85133486",
X"3d0d04fe",
X"3d0d80fc",
X"88087033",
X"7081ff06",
X"70842a81",
X"32810655",
X"51525371",
X"802e8c38",
X"a8733480",
X"fc880851",
X"b8713471",
X"83e0800c",
X"843d0d04",
X"fe3d0d80",
X"fc880870",
X"337081ff",
X"0670852a",
X"81328106",
X"55515253",
X"71802e8c",
X"38987334",
X"80fc8808",
X"51b87134",
X"7183e080",
X"0c843d0d",
X"04803d0d",
X"80fc8408",
X"51937134",
X"80fc9008",
X"51ff7134",
X"823d0d04",
X"fe3d0d02",
X"93053380",
X"fc840853",
X"53807234",
X"8a51d3c0",
X"3fd33f80",
X"fc940852",
X"80f87234",
X"80fcac08",
X"52807234",
X"fa1380fc",
X"b4085353",
X"72723480",
X"fc9c0852",
X"80723480",
X"fca40852",
X"72723480",
X"fc880852",
X"80723480",
X"fc880852",
X"b8723484",
X"3d0d04ff",
X"3d0d028f",
X"053380fc",
X"8c085252",
X"717134fe",
X"9e3f83e0",
X"8008802e",
X"f638833d",
X"0d04803d",
X"0d8439dc",
X"b03ffeb8",
X"3f83e080",
X"08802ef3",
X"3880fc8c",
X"08703370",
X"81ff0683",
X"e0800c51",
X"51823d0d",
X"04803d0d",
X"80fc8408",
X"51a37134",
X"80fc9008",
X"51ff7134",
X"80fc8808",
X"51a87134",
X"80fc8808",
X"51b87134",
X"823d0d04",
X"803d0d80",
X"fc840870",
X"337081c0",
X"06703070",
X"802583e0",
X"800c5151",
X"5151823d",
X"0d04ff3d",
X"0d80fc88",
X"08703370",
X"81ff0670",
X"832a8132",
X"70810651",
X"51515252",
X"70802ee5",
X"38b07234",
X"80fc8808",
X"51b87134",
X"833d0d04",
X"803d0d80",
X"fcc00870",
X"08810683",
X"e0800c51",
X"823d0d04",
X"fd3d0d75",
X"77545480",
X"73259438",
X"73708105",
X"55335280",
X"fb905185",
X"9d3fff13",
X"53e93985",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"b5923f83",
X"e080087a",
X"27ee3874",
X"802e80dd",
X"38745275",
X"51b4fd3f",
X"83e08008",
X"75537652",
X"54b5a43f",
X"83e08008",
X"7a537552",
X"56b4e53f",
X"83e08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"e08008c5",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9f",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fc813f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd53f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbb13f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83e0900c",
X"7183e094",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383e090",
X"085283e0",
X"940851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"80c0a653",
X"51fc983f",
X"8052873d",
X"51d03f86",
X"3d0d04fd",
X"3d0d7570",
X"5254a58e",
X"3f83e080",
X"08145372",
X"742e9238",
X"ff137033",
X"535371af",
X"2e098106",
X"ee388113",
X"537283e0",
X"800c853d",
X"0d04fd3d",
X"0d757770",
X"535454c7",
X"3f83e080",
X"08732ea1",
X"3883e080",
X"08733152",
X"ff125271",
X"ff2e8f38",
X"72708105",
X"54337470",
X"81055634",
X"eb39ff14",
X"54807434",
X"853d0d04",
X"803d0d72",
X"51ff903f",
X"823d0d04",
X"7183e080",
X"0c04803d",
X"0d725180",
X"7134810b",
X"bc120c80",
X"0b80c012",
X"0c823d0d",
X"04800b83",
X"e5bc0824",
X"8a38a5f8",
X"3fff0b83",
X"e5bc0c80",
X"0b83e080",
X"0c04ff3d",
X"0d735283",
X"e3980872",
X"2e8d38d9",
X"3f715197",
X"853f7183",
X"e3980c83",
X"3d0d04f4",
X"3d0d7e60",
X"625c5a55",
X"8154bc15",
X"08819138",
X"7451cf3f",
X"7958807a",
X"2580f738",
X"83e5ec08",
X"70892a57",
X"83ff0678",
X"84807231",
X"56565773",
X"78258338",
X"73557583",
X"e5bc082e",
X"8438ff89",
X"3f83e5bc",
X"088025a6",
X"3875892b",
X"5199f13f",
X"83e5ec08",
X"8f3dfc11",
X"555c5481",
X"52f81b51",
X"97d63f76",
X"1483e5ec",
X"0c7583e5",
X"bc0c7453",
X"76527851",
X"a4a93f83",
X"e0800883",
X"e5ec0816",
X"83e5ec0c",
X"78763176",
X"1b5b5956",
X"778024ff",
X"8b38617a",
X"710c5475",
X"5475802e",
X"83388154",
X"7383e080",
X"0c8e3d0d",
X"04fc3d0d",
X"fe9b3f76",
X"51feaf3f",
X"863dfc05",
X"5302a205",
X"22527751",
X"96f63f79",
X"863d2271",
X"0c5483e0",
X"80085483",
X"e0800880",
X"2e833881",
X"547383e0",
X"800c863d",
X"0d04fd3d",
X"0d7683e5",
X"bc085353",
X"80722489",
X"3871732e",
X"8438fdd1",
X"3f7551fd",
X"e53f7251",
X"98be3f73",
X"5273802e",
X"83388152",
X"7183e080",
X"0c853d0d",
X"04803d0d",
X"7280c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d72bc11",
X"0883e080",
X"0c51823d",
X"0d0480c4",
X"0b83e080",
X"0c04fd3d",
X"0d757771",
X"54705355",
X"53a0e73f",
X"82c81308",
X"bc150c82",
X"c0130880",
X"c0150cfc",
X"ec3f7351",
X"94983f73",
X"83e3980c",
X"83e08008",
X"5383e080",
X"08802e83",
X"38815372",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"775553fc",
X"c03f7280",
X"2ea538bc",
X"13085273",
X"519ff13f",
X"83e08008",
X"8f387752",
X"7251ff9a",
X"3f83e080",
X"08538a39",
X"82cc1308",
X"53d83981",
X"537283e0",
X"800c853d",
X"0d04fe3d",
X"0dff0b83",
X"e5bc0c74",
X"83e39c0c",
X"7583e5b8",
X"0ca0de3f",
X"83e08008",
X"81ff0652",
X"81537199",
X"3883e5d4",
X"518f903f",
X"83e08008",
X"5283e080",
X"08802e83",
X"38725271",
X"537283e0",
X"800c843d",
X"0d04fa3d",
X"0d787a82",
X"c4120882",
X"c4120870",
X"72245956",
X"56575773",
X"732e0981",
X"06913880",
X"c0165280",
X"c017519d",
X"e23f83e0",
X"80085574",
X"83e0800c",
X"883d0d04",
X"f63d0d7c",
X"5b807b71",
X"5c54577a",
X"772e8c38",
X"811a82cc",
X"1408545a",
X"72f63880",
X"5980d939",
X"7a548157",
X"80707b7b",
X"315a5755",
X"ff185374",
X"732580c1",
X"3882cc14",
X"08527351",
X"ff8c3f80",
X"0b83e080",
X"0825a138",
X"82cc1408",
X"82cc1108",
X"82cc160c",
X"7482cc12",
X"0c537580",
X"2e863872",
X"82cc170c",
X"72548057",
X"7382cc15",
X"08811757",
X"5556ffb8",
X"39811959",
X"800bff1b",
X"54547873",
X"25833881",
X"54768132",
X"70750651",
X"5372ff90",
X"388c3d0d",
X"04f73d0d",
X"7b7d5a5a",
X"82d05283",
X"e5b80851",
X"a89e3f83",
X"e0800857",
X"f9e33f79",
X"5283e5c0",
X"5196c73f",
X"83e08008",
X"53805483",
X"e0800874",
X"2e098106",
X"82833883",
X"e39c080b",
X"0b80fad8",
X"53705255",
X"9da03f0b",
X"0b80fad8",
X"5280c015",
X"519d933f",
X"74bc160c",
X"7282c016",
X"0c810b82",
X"c4160c81",
X"0b82c816",
X"0cff1773",
X"57578197",
X"3983e3a8",
X"3370822a",
X"70810651",
X"54547281",
X"86387381",
X"2a810658",
X"7780fc38",
X"76802e81",
X"903882d0",
X"15ff1875",
X"842a8106",
X"82c4130c",
X"83e3a833",
X"810682c8",
X"130c7b54",
X"71535856",
X"9cb43f75",
X"519ccb3f",
X"83e08008",
X"1653af73",
X"70810555",
X"3472bc17",
X"0c83e3a9",
X"5272519c",
X"953f83e3",
X"a00882c0",
X"170c83e3",
X"b6528390",
X"15519c82",
X"3f7782cc",
X"170c7880",
X"2e8d3875",
X"51782d83",
X"e0800880",
X"2e8d3874",
X"802e8638",
X"7582cc16",
X"0c755583",
X"e3a05283",
X"e5c05195",
X"e73f83e0",
X"80088a38",
X"83e3a933",
X"5372fed1",
X"38800b82",
X"cc170c78",
X"802e8938",
X"83e39c08",
X"51fcb93f",
X"83e39c08",
X"547383e0",
X"800c8b3d",
X"0d04ff3d",
X"0d805273",
X"51fdb63f",
X"833d0d04",
X"f03d0d62",
X"705254f6",
X"923f83e0",
X"80087453",
X"873d7053",
X"5555f6b2",
X"3ff7923f",
X"7351d33f",
X"63537452",
X"83e08008",
X"51fab93f",
X"923d0d04",
X"7183e080",
X"0c0480c0",
X"1283e080",
X"0c04803d",
X"0d7282c0",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"cc110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"82c41108",
X"83e0800c",
X"51823d0d",
X"04f63d0d",
X"7c83e098",
X"08595981",
X"792782a9",
X"38788819",
X"082782a1",
X"38773356",
X"75822e81",
X"9b387582",
X"24893875",
X"812e8d38",
X"828b3975",
X"832e81b7",
X"38828239",
X"7883ffff",
X"0670812a",
X"117083ff",
X"ff067083",
X"ff067189",
X"2a903d5f",
X"525a5151",
X"557683ff",
X"2e8e3882",
X"5476538c",
X"18081552",
X"7951a939",
X"75547653",
X"8c180815",
X"5279519a",
X"d83f83e0",
X"800881bd",
X"38755483",
X"e0800853",
X"8c180815",
X"8105528c",
X"3dfd0551",
X"9abb3f83",
X"e0800881",
X"a03802a9",
X"05338c3d",
X"3371882b",
X"077a8106",
X"71842a53",
X"57585674",
X"8638769f",
X"ff065675",
X"55818039",
X"75547810",
X"83fe0653",
X"78882a8c",
X"19080552",
X"8c3dfc05",
X"5199fa3f",
X"83e08008",
X"80df3802",
X"a905338c",
X"3d337188",
X"2b075657",
X"80d13984",
X"5478822b",
X"83fc0653",
X"78872a8c",
X"19080552",
X"8c3dfc05",
X"5199ca3f",
X"83e08008",
X"b03802ab",
X"05330284",
X"05aa0533",
X"71982b71",
X"902b0702",
X"8c05a905",
X"3370882b",
X"7207903d",
X"337180ff",
X"fffe8006",
X"07515253",
X"57585683",
X"39815574",
X"83e0800c",
X"8c3d0d04",
X"fb3d0d83",
X"e09808fe",
X"19881208",
X"fe055556",
X"54805674",
X"73278d38",
X"82143375",
X"71299416",
X"08055753",
X"7583e080",
X"0c873d0d",
X"04fc3d0d",
X"7683e098",
X"08555580",
X"75238815",
X"08537281",
X"2e883888",
X"14087326",
X"85388152",
X"b2397290",
X"38733352",
X"71832e09",
X"81068538",
X"90140853",
X"728c160c",
X"72802e8d",
X"387251ff",
X"933f83e0",
X"80085285",
X"39901408",
X"52719016",
X"0c805271",
X"83e0800c",
X"863d0d04",
X"fa3d0d78",
X"83e09808",
X"71228105",
X"7083ffff",
X"06575457",
X"5573802e",
X"88389015",
X"08537286",
X"38835280",
X"e739738f",
X"06527180",
X"da388113",
X"90160c8c",
X"15085372",
X"9038830b",
X"84172257",
X"52737627",
X"80c638bf",
X"39821633",
X"ff057484",
X"2a065271",
X"b2387251",
X"fbdb3f81",
X"527183e0",
X"800827a8",
X"38835283",
X"e0800888",
X"1708279c",
X"3883e080",
X"088c160c",
X"83e08008",
X"51fdf93f",
X"83e08008",
X"90160c73",
X"75238052",
X"7183e080",
X"0c883d0d",
X"04f23d0d",
X"60626458",
X"5d5b7533",
X"5574a02e",
X"09810688",
X"38811670",
X"4456ef39",
X"62703356",
X"5674af2e",
X"09810684",
X"38811643",
X"800b881c",
X"0c627033",
X"515574a0",
X"2691387a",
X"51fdd23f",
X"83e08008",
X"56807c34",
X"83a83993",
X"3d841c08",
X"70585a5f",
X"8a55a076",
X"70810558",
X"34ff1555",
X"74ff2e09",
X"8106ef38",
X"8070595d",
X"887f085f",
X"5a7c811e",
X"7081ff06",
X"60137033",
X"70af3270",
X"30a07327",
X"71802507",
X"5151525b",
X"535f5755",
X"7480d838",
X"76ae2e09",
X"81068338",
X"8155777a",
X"27750755",
X"74802e9f",
X"38798832",
X"703078ae",
X"32703070",
X"73079f2a",
X"53515751",
X"5675ac38",
X"88588b5a",
X"ffab39ff",
X"9f175574",
X"99268938",
X"e0177081",
X"ff065855",
X"77811970",
X"81ff0672",
X"1c535a57",
X"55767534",
X"ff87397c",
X"1e7f0c80",
X"5576a026",
X"83388155",
X"748b1a34",
X"7a51fc91",
X"3f83e080",
X"0880f538",
X"a0547a22",
X"70852b83",
X"e0065455",
X"901b0852",
X"7b5194d1",
X"3f83e080",
X"085783e0",
X"80088182",
X"387b3355",
X"74802e80",
X"f5388b1c",
X"3370832a",
X"70810651",
X"565674b4",
X"388b7c84",
X"1d0883e0",
X"8008595b",
X"5b58ff18",
X"5877ff2e",
X"9a387970",
X"81055b33",
X"79708105",
X"5b337171",
X"31525656",
X"75802ee2",
X"38863975",
X"802ebc38",
X"7a51fbf4",
X"3fff8639",
X"83e08008",
X"5683e080",
X"08802ea9",
X"3883e080",
X"08832e09",
X"810680de",
X"38841b08",
X"8b113351",
X"557480d2",
X"38845680",
X"cd398356",
X"ec398156",
X"80c43976",
X"56841b08",
X"8b113351",
X"5574b738",
X"8b1c3370",
X"842a7081",
X"06515657",
X"74802ed5",
X"38951c33",
X"941d3371",
X"982b7190",
X"2b079b1f",
X"337f9a05",
X"3371882b",
X"0772077f",
X"88050c5a",
X"585658fc",
X"da397583",
X"e0800c90",
X"3d0d04f8",
X"3d0d7a7c",
X"59578254",
X"83fe5377",
X"52765192",
X"e03f8356",
X"83e08008",
X"80ec3881",
X"17337733",
X"71882b07",
X"56568256",
X"7482d4d5",
X"2e098106",
X"80d43875",
X"54b65377",
X"52765192",
X"b43f83e0",
X"80089838",
X"81173377",
X"3371882b",
X"0783e080",
X"08525656",
X"748182c6",
X"2eac3882",
X"5480d253",
X"77527651",
X"928b3f83",
X"e0800898",
X"38811733",
X"77337188",
X"2b0783e0",
X"80085256",
X"56748182",
X"c62e8338",
X"81567583",
X"e0800c8a",
X"3d0d04ec",
X"3d0d6659",
X"800b83e0",
X"980c7856",
X"78802e83",
X"e83891a5",
X"3f83e080",
X"08810655",
X"82567483",
X"d8387475",
X"538e3d70",
X"535858fe",
X"c23f83e0",
X"800881ff",
X"06567581",
X"2e098106",
X"80d43890",
X"5483be53",
X"74527651",
X"91973f83",
X"e0800880",
X"c9388e3d",
X"33557480",
X"2e80c938",
X"02bb0533",
X"028405ba",
X"05337198",
X"2b71902b",
X"07028c05",
X"b9053370",
X"882b7207",
X"943d3371",
X"0770587c",
X"5754525d",
X"575956fd",
X"e63f83e0",
X"800881ff",
X"06567583",
X"2e098106",
X"86388156",
X"82db3975",
X"802e8638",
X"875682d1",
X"39a4548d",
X"53775276",
X"5190ae3f",
X"815683e0",
X"800882bd",
X"3802ba05",
X"33028405",
X"b9053371",
X"882b0758",
X"5c76ab38",
X"0280ca05",
X"33028405",
X"80c90533",
X"71982b71",
X"902b0796",
X"3d337088",
X"2b720702",
X"940580c7",
X"05337107",
X"54525d57",
X"585602b3",
X"05337771",
X"29028805",
X"b2053302",
X"8c05b105",
X"3371882b",
X"07701c70",
X"8c1f0c5e",
X"5957585c",
X"8d3d3382",
X"1a3402b5",
X"05338f3d",
X"3371882b",
X"07595b77",
X"841a2302",
X"b7053302",
X"8405b605",
X"3371882b",
X"07565b74",
X"ab380280",
X"c6053302",
X"840580c5",
X"05337198",
X"2b71902b",
X"07953d33",
X"70882b72",
X"07029405",
X"80c30533",
X"71075152",
X"53575d5b",
X"74763177",
X"3178842a",
X"8f3d3354",
X"71713153",
X"56569880",
X"3f83e080",
X"08820570",
X"881b0c70",
X"9ff62681",
X"05575583",
X"fff67527",
X"83388356",
X"75793475",
X"832e0981",
X"06af3802",
X"80d20533",
X"02840580",
X"d1053371",
X"982b7190",
X"2b07983d",
X"3370882b",
X"72070294",
X"0580cf05",
X"33710790",
X"1f0c525d",
X"57595686",
X"39761a90",
X"1a0c8419",
X"228c1a08",
X"1871842a",
X"05941b0c",
X"5c800b81",
X"1a347883",
X"e0980c80",
X"567583e0",
X"800c963d",
X"0d04e93d",
X"0d83e098",
X"08568654",
X"75802e81",
X"a638800b",
X"81173499",
X"3de01146",
X"6a54c011",
X"53ec0551",
X"f6cf3f83",
X"e0800854",
X"83e08008",
X"81853889",
X"3d335473",
X"802e9338",
X"02ab0533",
X"70842a70",
X"81065155",
X"5573802e",
X"86388354",
X"80e53902",
X"b505338f",
X"3d337198",
X"2b71902b",
X"07028c05",
X"bb053302",
X"9005ba05",
X"3371882b",
X"077207a0",
X"1b0c0290",
X"05bf0533",
X"029405be",
X"05337198",
X"2b71902b",
X"07029c05",
X"bd053370",
X"882b7207",
X"993d3371",
X"077f9c05",
X"0c5283e0",
X"8008981f",
X"0c565a52",
X"52535759",
X"57810b81",
X"173483e0",
X"80085473",
X"83e0800c",
X"993d0d04",
X"f53d0d7d",
X"60028805",
X"ba052272",
X"83e09808",
X"5b5d5a5c",
X"5c807b23",
X"86567680",
X"2e81e038",
X"81173381",
X"06558556",
X"74802e81",
X"d2389c17",
X"08981808",
X"31557478",
X"27873874",
X"83ffff06",
X"5877802e",
X"81ae3898",
X"17087083",
X"ff065656",
X"7480ca38",
X"821733ff",
X"0576892a",
X"067081ff",
X"065a5578",
X"a0387587",
X"38a01708",
X"558d39a4",
X"170851ef",
X"e03f83e0",
X"80085581",
X"752780f8",
X"3874a418",
X"0ca41708",
X"51f28d3f",
X"83e08008",
X"802e80e4",
X"3883e080",
X"0819a818",
X"0c981708",
X"83ff0684",
X"80713170",
X"83ffff06",
X"58515577",
X"76278338",
X"77567554",
X"98170883",
X"ff0653a8",
X"17085279",
X"557b8338",
X"7b557451",
X"8ad33f83",
X"e08008a4",
X"38981708",
X"1698180c",
X"751a7877",
X"317083ff",
X"ff067d22",
X"7905525a",
X"565a747b",
X"23fece39",
X"80568839",
X"800b8118",
X"34815675",
X"83e0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83e09808",
X"55568655",
X"73802e81",
X"dc388114",
X"33810653",
X"85557280",
X"2e81ce38",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"a9388214",
X"3370892b",
X"56537680",
X"2eb53874",
X"52ff1651",
X"92ee3f83",
X"e08008ff",
X"18765470",
X"53585392",
X"df3f83e0",
X"80087326",
X"96387430",
X"70780670",
X"98170c77",
X"7131a417",
X"08525851",
X"538939a0",
X"140870a4",
X"160c5374",
X"7627b438",
X"7251edc1",
X"3f83e080",
X"0853810b",
X"83e08008",
X"2780cb38",
X"83e08008",
X"88150827",
X"80c03883",
X"e08008a4",
X"150c9814",
X"08159815",
X"0c757531",
X"56c93998",
X"14081670",
X"98160c73",
X"5256efc8",
X"3f83e080",
X"08802e96",
X"38821433",
X"ff057689",
X"2a0683e0",
X"800805a8",
X"150c8055",
X"8839800b",
X"81153481",
X"557483e0",
X"800c883d",
X"0d04ee3d",
X"0d645686",
X"5583e098",
X"08802e80",
X"f638943d",
X"f4118418",
X"0c6654d4",
X"05527551",
X"f1973f83",
X"e0800855",
X"83e08008",
X"80cf3889",
X"3d335473",
X"802ebc38",
X"02ab0533",
X"70842a70",
X"81065155",
X"55845573",
X"802ebc38",
X"02b50533",
X"8f3d3371",
X"982b7190",
X"2b07028c",
X"05bb0533",
X"029005ba",
X"05337188",
X"2b077207",
X"881b0c53",
X"57595775",
X"51eed23f",
X"83e08008",
X"5574832e",
X"09810683",
X"38845574",
X"83e0800c",
X"943d0d04",
X"e43d0d6e",
X"a13d0840",
X"5d865683",
X"e0980880",
X"2e849b38",
X"9e3df405",
X"841e0c7e",
X"98387c51",
X"ee973f83",
X"e0800856",
X"84843981",
X"41828039",
X"834181fb",
X"39933d7f",
X"96054159",
X"807f8295",
X"055f5675",
X"6081ff05",
X"34834190",
X"1d08762e",
X"81dd38a0",
X"547c2270",
X"852b83e0",
X"06545890",
X"1d085278",
X"5186ae3f",
X"83e08008",
X"4183e080",
X"08ffb838",
X"78335c7b",
X"802effb4",
X"388b1933",
X"70bf0671",
X"81065243",
X"5574802e",
X"80e8387b",
X"81bf0655",
X"748f2480",
X"dd389a19",
X"33557480",
X"d5389c19",
X"33557480",
X"2e80cb38",
X"f31e7058",
X"5e815675",
X"8b2e0981",
X"0685388e",
X"568b3975",
X"9a2e0981",
X"0683389c",
X"56751970",
X"70810552",
X"33713381",
X"1a821a5f",
X"5b525b55",
X"74863879",
X"77348539",
X"80df7734",
X"777b5757",
X"7aa02e09",
X"8106c038",
X"81567b81",
X"e5327030",
X"709f2a51",
X"51557bae",
X"2e933874",
X"802e8e38",
X"61832a70",
X"81065155",
X"74802e97",
X"387c51ec",
X"f73f83e0",
X"80084183",
X"e0800887",
X"38901d08",
X"fea53880",
X"60347580",
X"2e88387d",
X"527f5183",
X"b13f6080",
X"2e863880",
X"0b901e0c",
X"60566083",
X"2e098106",
X"8838800b",
X"901e0c85",
X"396081d2",
X"38891f57",
X"901d0880",
X"2e81a838",
X"80567519",
X"70335155",
X"74a02ea0",
X"3874852e",
X"09810684",
X"3881e555",
X"74777081",
X"05593481",
X"167081ff",
X"06575587",
X"7627d738",
X"88193355",
X"74a02ea9",
X"38ae7770",
X"81055934",
X"88567519",
X"70335155",
X"74a02e95",
X"38747770",
X"81055934",
X"81167081",
X"ff065755",
X"8a7627e2",
X"388b1933",
X"7f880534",
X"9f19339e",
X"1a337198",
X"2b71902b",
X"079d1c33",
X"70882b72",
X"079c1e33",
X"7107640c",
X"52991d33",
X"981e3371",
X"882b0753",
X"51535759",
X"56747f84",
X"05239719",
X"33961a33",
X"71882b07",
X"5656747f",
X"86052380",
X"77347c51",
X"eafe3f83",
X"e0800856",
X"83e08008",
X"832e0981",
X"06883880",
X"0b901e0c",
X"8056961f",
X"3355748a",
X"38891f52",
X"961f5181",
X"b13f7583",
X"e0800c9e",
X"3d0d04fd",
X"3d0d7577",
X"53547333",
X"51708938",
X"71335170",
X"802ea138",
X"73337233",
X"52537271",
X"278538ff",
X"51943970",
X"73278538",
X"81518b39",
X"81148113",
X"5354d339",
X"80517083",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"54547233",
X"7081ff06",
X"52527080",
X"2ea33871",
X"81ff0681",
X"14ffbf12",
X"53545270",
X"99268938",
X"a0127081",
X"ff065351",
X"71747081",
X"055634d2",
X"39807434",
X"853d0d04",
X"ffbd3d0d",
X"80c63d08",
X"52a53d70",
X"5254ffb3",
X"3f80c73d",
X"0852853d",
X"705253ff",
X"a63f7252",
X"7351fedf",
X"3f80c53d",
X"0d04fe3d",
X"0d747653",
X"53717081",
X"05533351",
X"70737081",
X"05553470",
X"f038843d",
X"0d04fe3d",
X"0d745280",
X"72335253",
X"70732e8d",
X"38811281",
X"14713353",
X"545270f5",
X"387283e0",
X"800c843d",
X"0d04fc3d",
X"0d765574",
X"83e68008",
X"2eaf3880",
X"53745187",
X"cd3f83e0",
X"800881ff",
X"06ff1470",
X"81ff0672",
X"30709f2a",
X"51525553",
X"5472802e",
X"843871dd",
X"3873fe38",
X"7483e680",
X"0c863d0d",
X"04ff3d0d",
X"ff0b83e6",
X"800c84af",
X"3f815187",
X"913f83e0",
X"800881ff",
X"065271ee",
X"3881d63f",
X"7183e080",
X"0c833d0d",
X"04fc3d0d",
X"76028405",
X"a2052202",
X"8805a605",
X"227a5455",
X"5555ff82",
X"3f72802e",
X"a03883e6",
X"94143375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552dd",
X"39800b83",
X"e0800c86",
X"3d0d04fc",
X"3d0d7678",
X"7a115653",
X"55805371",
X"742e9338",
X"72155170",
X"3383e694",
X"13348112",
X"81145452",
X"ea39800b",
X"83e0800c",
X"863d0d04",
X"fd3d0d90",
X"5483e680",
X"08518780",
X"3f83e080",
X"0881ff06",
X"ff157130",
X"71307073",
X"079f2a72",
X"9f2a0652",
X"55525553",
X"72db3885",
X"3d0d04ff",
X"3d0d83e6",
X"8c081083",
X"e6840807",
X"80fcc408",
X"52710c83",
X"3d0d0480",
X"0b83e68c",
X"0ce13f04",
X"810b83e6",
X"8c0cd83f",
X"04ed3f04",
X"7183e688",
X"0c04803d",
X"0d8051f4",
X"3f810b83",
X"e68c0c81",
X"0b83e684",
X"0cffb83f",
X"823d0d04",
X"803d0d72",
X"30707407",
X"802583e6",
X"840c51ff",
X"a23f823d",
X"0d04fe3d",
X"0d029305",
X"3380fcc8",
X"0854730c",
X"80fcc408",
X"52710870",
X"81065151",
X"70f73872",
X"087081ff",
X"0683e080",
X"0c51843d",
X"0d04803d",
X"0d81ff51",
X"cd3f83e0",
X"800881ff",
X"0683e080",
X"0c823d0d",
X"04ff3d0d",
X"74902b74",
X"0780fcb8",
X"0852710c",
X"833d0d04",
X"04fb3d0d",
X"78028405",
X"9f053370",
X"982b5557",
X"55728025",
X"9b387580",
X"ff065680",
X"5280f751",
X"e03f83e0",
X"800881ff",
X"06547381",
X"2680ff38",
X"8051fee0",
X"3fff9f3f",
X"8151fed8",
X"3fff973f",
X"7551fee6",
X"3f74982a",
X"51fedf3f",
X"74902a70",
X"81ff0652",
X"53fed33f",
X"74882a70",
X"81ff0652",
X"53fec73f",
X"7481ff06",
X"51febf3f",
X"81557580",
X"c02e0981",
X"06863881",
X"95558d39",
X"7580c82e",
X"09810684",
X"38818755",
X"7451fe9e",
X"3f8a55fe",
X"c53f83e0",
X"800881ff",
X"0670982b",
X"54547280",
X"258c38ff",
X"157081ff",
X"06565374",
X"e2387383",
X"e0800c87",
X"3d0d04fa",
X"3d0dfdbe",
X"3f8051fd",
X"d33f8a54",
X"fe903fff",
X"147081ff",
X"06555373",
X"f3387374",
X"535580c0",
X"51fea63f",
X"83e08008",
X"81ff0654",
X"73812e09",
X"810682a1",
X"3883aa52",
X"80c851fe",
X"8c3f83e0",
X"800881ff",
X"06537281",
X"2e098106",
X"81a93874",
X"54873d74",
X"115456fd",
X"c53f83e0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e5",
X"38029a05",
X"33537281",
X"2e098106",
X"81db3802",
X"9b053353",
X"80ce9054",
X"7281aa2e",
X"8e3881c9",
X"3980e451",
X"ff9fdd3f",
X"ff145473",
X"802e81b9",
X"38820a52",
X"81e951fd",
X"a43f83e0",
X"800881ff",
X"065372dd",
X"38725280",
X"fa51fd91",
X"3f83e080",
X"0881ff06",
X"53728191",
X"38725473",
X"1653fcd2",
X"3f83e080",
X"08733481",
X"147081ff",
X"06555383",
X"7427e838",
X"873d3370",
X"862a7081",
X"06515454",
X"8c557280",
X"e4388455",
X"80df3974",
X"5281e951",
X"fccb3f83",
X"e0800881",
X"ff065382",
X"5581e956",
X"81732786",
X"38735580",
X"c15680ce",
X"90548b39",
X"80e451ff",
X"9ece3fff",
X"14547380",
X"2ea93880",
X"527551fc",
X"983f83e0",
X"800881ff",
X"065372e0",
X"38848052",
X"80d051fc",
X"843f83e0",
X"800881ff",
X"06537280",
X"2e833880",
X"557483e6",
X"90348051",
X"fafe3ffb",
X"bd3f883d",
X"0d04fb3d",
X"0d775480",
X"0b83e690",
X"3370832a",
X"70810651",
X"55575572",
X"752e0981",
X"06853873",
X"892b5473",
X"5280d151",
X"fbbb3f83",
X"e0800881",
X"ff065372",
X"bd3882b8",
X"c054fafe",
X"3f83e080",
X"0881ff06",
X"537281ff",
X"2e098106",
X"8938ff14",
X"5473e738",
X"9f397281",
X"fe2e0981",
X"06963883",
X"ea945283",
X"e69451fa",
X"e83fface",
X"3ffacb3f",
X"83398155",
X"8051fa80",
X"3ffabf3f",
X"7481ff06",
X"83e0800c",
X"873d0d04",
X"fb3d0d77",
X"83e69456",
X"548151f9",
X"e33f83e6",
X"90337083",
X"2a708106",
X"51545672",
X"85387389",
X"2b547352",
X"80d851fa",
X"b43f83e0",
X"800881ff",
X"06537280",
X"e53881ff",
X"51f9cb3f",
X"81fe51f9",
X"c53f8480",
X"53747081",
X"05563351",
X"f9b83fff",
X"137083ff",
X"ff065153",
X"72eb3872",
X"51f9a73f",
X"7251f9a2",
X"3ff9cb3f",
X"83e08008",
X"9f0653a7",
X"88547285",
X"2e8d389a",
X"3980e451",
X"ff9c853f",
X"ff1454f9",
X"ad3f83e0",
X"800881ff",
X"2e843873",
X"e8388051",
X"f8da3ff9",
X"993f800b",
X"83e0800c",
X"873d0d04",
X"83e08c08",
X"0283e08c",
X"0cfd3d0d",
X"805383e0",
X"8c088c05",
X"085283e0",
X"8c088805",
X"085183d4",
X"3f83e080",
X"087083e0",
X"800c5485",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"fd3d0d81",
X"5383e08c",
X"088c0508",
X"5283e08c",
X"08880508",
X"5183a13f",
X"83e08008",
X"7083e080",
X"0c54853d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cf9",
X"3d0d800b",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"05088025",
X"b93883e0",
X"8c088805",
X"083083e0",
X"8c088805",
X"0c800b83",
X"e08c08f4",
X"050c83e0",
X"8c08fc05",
X"088a3881",
X"0b83e08c",
X"08f4050c",
X"83e08c08",
X"f4050883",
X"e08c08fc",
X"050c83e0",
X"8c088c05",
X"088025b9",
X"3883e08c",
X"088c0508",
X"3083e08c",
X"088c050c",
X"800b83e0",
X"8c08f005",
X"0c83e08c",
X"08fc0508",
X"8a38810b",
X"83e08c08",
X"f0050c83",
X"e08c08f0",
X"050883e0",
X"8c08fc05",
X"0c805383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"05085181",
X"df3f83e0",
X"80087083",
X"e08c08f8",
X"050c5483",
X"e08c08fc",
X"0508802e",
X"903883e0",
X"8c08f805",
X"083083e0",
X"8c08f805",
X"0c83e08c",
X"08f80508",
X"7083e080",
X"0c54893d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cfb",
X"3d0d800b",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"05088025",
X"993883e0",
X"8c088805",
X"083083e0",
X"8c088805",
X"0c810b83",
X"e08c08fc",
X"050c83e0",
X"8c088c05",
X"08802590",
X"3883e08c",
X"088c0508",
X"3083e08c",
X"088c050c",
X"815383e0",
X"8c088c05",
X"085283e0",
X"8c088805",
X"0851bd3f",
X"83e08008",
X"7083e08c",
X"08f8050c",
X"5483e08c",
X"08fc0508",
X"802e9038",
X"83e08c08",
X"f8050830",
X"83e08c08",
X"f8050c83",
X"e08c08f8",
X"05087083",
X"e0800c54",
X"873d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cfd3d0d",
X"810b83e0",
X"8c08fc05",
X"0c800b83",
X"e08c08f8",
X"050c83e0",
X"8c088c05",
X"0883e08c",
X"08880508",
X"27b93883",
X"e08c08fc",
X"0508802e",
X"ae38800b",
X"83e08c08",
X"8c050824",
X"a23883e0",
X"8c088c05",
X"081083e0",
X"8c088c05",
X"0c83e08c",
X"08fc0508",
X"1083e08c",
X"08fc050c",
X"ffb83983",
X"e08c08fc",
X"0508802e",
X"80e13883",
X"e08c088c",
X"050883e0",
X"8c088805",
X"0826ad38",
X"83e08c08",
X"88050883",
X"e08c088c",
X"05083183",
X"e08c0888",
X"050c83e0",
X"8c08f805",
X"0883e08c",
X"08fc0508",
X"0783e08c",
X"08f8050c",
X"83e08c08",
X"fc050881",
X"2a83e08c",
X"08fc050c",
X"83e08c08",
X"8c050881",
X"2a83e08c",
X"088c050c",
X"ff953983",
X"e08c0890",
X"0508802e",
X"933883e0",
X"8c088805",
X"087083e0",
X"8c08f405",
X"0c519139",
X"83e08c08",
X"f8050870",
X"83e08c08",
X"f4050c51",
X"83e08c08",
X"f4050883",
X"e0800c85",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"ff3d0d80",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"88050881",
X"06ff1170",
X"097083e0",
X"8c088c05",
X"080683e0",
X"8c08fc05",
X"081183e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"812a83e0",
X"8c088805",
X"0c83e08c",
X"088c0508",
X"1083e08c",
X"088c050c",
X"51515151",
X"83e08c08",
X"88050880",
X"2e8438ff",
X"ab3983e0",
X"8c08fc05",
X"087083e0",
X"800c5183",
X"3d0d83e0",
X"8c0c04fc",
X"3d0d7670",
X"797b5555",
X"55558f72",
X"278c3872",
X"75078306",
X"5170802e",
X"a938ff12",
X"5271ff2e",
X"98387270",
X"81055433",
X"74708105",
X"5634ff12",
X"5271ff2e",
X"098106ea",
X"387483e0",
X"800c863d",
X"0d047451",
X"72708405",
X"54087170",
X"8405530c",
X"72708405",
X"54087170",
X"8405530c",
X"72708405",
X"54087170",
X"8405530c",
X"72708405",
X"54087170",
X"8405530c",
X"f0125271",
X"8f26c938",
X"83722795",
X"38727084",
X"05540871",
X"70840553",
X"0cfc1252",
X"718326ed",
X"387054ff",
X"81390000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"000009a5",
X"000009e6",
X"00000a08",
X"00000a26",
X"00000a26",
X"00000a26",
X"00000a26",
X"00000a95",
X"00000ac5",
X"70704740",
X"9c704268",
X"9c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"43617274",
X"72696467",
X"6520386b",
X"2073696d",
X"706c6500",
X"45786974",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"25732025",
X"73000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"524f4d00",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"6e616d65",
X"20000000",
X"25303278",
X"00000000",
X"00000000",
X"00000000",
X"00003c9c",
X"00003ca0",
X"00003ca8",
X"00003cb4",
X"00003cc0",
X"00003ccc",
X"00003cd8",
X"00003cdc",
X"0001d20f",
X"0001d400",
X"0001d401",
X"0001d409",
X"0001d010",
X"0001d301",
X"0001d300",
X"0001d20a",
X"0001d01b",
X"0001d016",
X"0001d019",
X"0001d018",
X"0001d017",
X"0001d01a",
X"0001d403",
X"0001d402",
X"0001d40e",
X"0004007c",
X"00040078",
X"00040074",
X"00040068",
X"00040060",
X"0004005c",
X"00040058",
X"00040054",
X"00040050",
X"0004004c",
X"00040048",
X"00040044",
X"00040040",
X"00040034",
X"00040030",
X"0004002c",
X"00040028",
X"00040024",
X"00040020",
X"0004001c",
X"00040018",
X"00040014",
X"00040010",
X"0004000c",
X"00040008",
X"00040004",
X"00040000",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
