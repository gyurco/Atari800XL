
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81ea",
X"fc738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81f3",
X"e80c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757580f7",
X"932d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7580f6d2",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80e0e004",
X"fd3d0d75",
X"705254ae",
X"aa3f83c0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"c0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83c0",
X"8008732e",
X"a13883c0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183c0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83c2d008",
X"248a38b4",
X"fb3fff0b",
X"83c2d00c",
X"800b83c0",
X"800c04ff",
X"3d0d7352",
X"83c0ac08",
X"722e8d38",
X"d93f7151",
X"96a03f71",
X"83c0ac0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"55805681",
X"54bc1508",
X"762e0981",
X"06819138",
X"7451c83f",
X"7958757a",
X"2580f738",
X"83c38008",
X"70892a57",
X"83ff0678",
X"84807231",
X"56565773",
X"78258338",
X"73557583",
X"c2d0082e",
X"8438ff82",
X"3f83c2d0",
X"088025a6",
X"3875892b",
X"5198dc3f",
X"83c38008",
X"8f3dfc11",
X"555c5481",
X"52f81b51",
X"96c63f76",
X"1483c380",
X"0c7583c2",
X"d00c7453",
X"76527851",
X"b3a53f83",
X"c0800883",
X"c3800816",
X"83c3800c",
X"78763176",
X"1b5b5956",
X"778024ff",
X"8b38617a",
X"710c5475",
X"5475802e",
X"83388154",
X"7383c080",
X"0c8e3d0d",
X"04fc3d0d",
X"fe943f76",
X"51fea83f",
X"863dfc05",
X"53785277",
X"5195e93f",
X"7975710c",
X"5483c080",
X"085483c0",
X"8008802e",
X"83388154",
X"7383c080",
X"0c863d0d",
X"04fe3d0d",
X"7583c2d0",
X"08535380",
X"72248938",
X"71732e84",
X"38fdcf3f",
X"7451fde3",
X"3f725197",
X"ae3f83c0",
X"80085283",
X"c0800880",
X"2e833881",
X"527183c0",
X"800c843d",
X"0d04803d",
X"0d7280c0",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"3d0d72bc",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"c40b83c0",
X"800c04fd",
X"3d0d7577",
X"71547053",
X"5553a9fb",
X"3f82c813",
X"08bc150c",
X"82c01308",
X"80c0150c",
X"fce43f73",
X"5193ab3f",
X"7383c0ac",
X"0c83c080",
X"085383c0",
X"8008802e",
X"83388153",
X"7283c080",
X"0c853d0d",
X"04fd3d0d",
X"75775553",
X"fcb83f72",
X"802ea538",
X"bc130852",
X"7351a985",
X"3f83c080",
X"088f3877",
X"527251ff",
X"9a3f83c0",
X"8008538a",
X"3982cc13",
X"0853d839",
X"81537283",
X"c0800c85",
X"3d0d04fe",
X"3d0dff0b",
X"83c2d00c",
X"7483c0b0",
X"0c7583c2",
X"cc0cafd9",
X"3f83c080",
X"0881ff06",
X"52815371",
X"993883c2",
X"e8518e94",
X"3f83c080",
X"085283c0",
X"8008802e",
X"83387252",
X"71537283",
X"c0800c84",
X"3d0d04fa",
X"3d0d787a",
X"82c41208",
X"82c41208",
X"70722459",
X"56565757",
X"73732e09",
X"81069138",
X"80c01652",
X"80c01751",
X"a6f63f83",
X"c0800855",
X"7483c080",
X"0c883d0d",
X"04f63d0d",
X"7c5b807b",
X"715c5457",
X"7a772e8c",
X"38811a82",
X"cc140854",
X"5a72f638",
X"805980d9",
X"397a5481",
X"5780707b",
X"7b315a57",
X"55ff1853",
X"74732580",
X"c13882cc",
X"14085273",
X"51ff8c3f",
X"800b83c0",
X"800825a1",
X"3882cc14",
X"0882cc11",
X"0882cc16",
X"0c7482cc",
X"120c5375",
X"802e8638",
X"7282cc17",
X"0c725480",
X"577382cc",
X"15088117",
X"575556ff",
X"b8398119",
X"59800bff",
X"1b545478",
X"73258338",
X"81547681",
X"32707506",
X"515372ff",
X"90388c3d",
X"0d04f73d",
X"0d7b7d5a",
X"5a82d052",
X"83c2cc08",
X"5180e5ce",
X"3f83c080",
X"0857f9da",
X"3f795283",
X"c2d45195",
X"b73f83c0",
X"80085480",
X"5383c080",
X"08732e09",
X"81068283",
X"3883c0b0",
X"080b0b81",
X"f0985370",
X"5256a6b3",
X"3f0b0b81",
X"f0985280",
X"c01651a6",
X"a63f75bc",
X"170c7382",
X"c0170c81",
X"0b82c417",
X"0c810b82",
X"c8170c73",
X"82cc170c",
X"ff1782d0",
X"17555781",
X"913983c0",
X"bc337082",
X"2a708106",
X"51545572",
X"81803874",
X"812a8106",
X"587780f6",
X"3874842a",
X"810682c4",
X"150c83c0",
X"bc338106",
X"82c8150c",
X"79527351",
X"a5cd3f73",
X"51a5e43f",
X"83c08008",
X"1453af73",
X"70810555",
X"3472bc15",
X"0c83c0bd",
X"527251a5",
X"ae3f83c0",
X"b40882c0",
X"150c83c0",
X"ca5280c0",
X"1451a59b",
X"3f78802e",
X"8d387351",
X"782d83c0",
X"8008802e",
X"99387782",
X"cc150c75",
X"802e8638",
X"7382cc17",
X"0c7382d0",
X"15ff1959",
X"55567680",
X"2e9b3883",
X"c0b45283",
X"c2d45194",
X"ad3f83c0",
X"80088a38",
X"83c0bd33",
X"5372fed2",
X"3878802e",
X"893883c0",
X"b00851fc",
X"b83f83c0",
X"b0085372",
X"83c0800c",
X"8b3d0d04",
X"ff3d0d80",
X"527351fd",
X"b53f833d",
X"0d04f03d",
X"0d627052",
X"54f6893f",
X"83c08008",
X"7453873d",
X"70535555",
X"f6a93ff7",
X"893f7351",
X"d33f6353",
X"745283c0",
X"800851fa",
X"b83f923d",
X"0d047183",
X"c0800c04",
X"80c01283",
X"c0800c04",
X"803d0d72",
X"82c01108",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"7282cc11",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d7282c4",
X"110883c0",
X"800c5182",
X"3d0d04f9",
X"3d0d7983",
X"c0900857",
X"57817727",
X"81963876",
X"88170827",
X"818e3875",
X"33557482",
X"2e893874",
X"832eb338",
X"80fe3974",
X"54761083",
X"fe065376",
X"882a8c17",
X"08055289",
X"3dfc0551",
X"aa873f83",
X"c0800880",
X"df38029d",
X"0533893d",
X"3371882b",
X"07565680",
X"d1398454",
X"76822b83",
X"fc065376",
X"872a8c17",
X"08055289",
X"3dfc0551",
X"a9d73f83",
X"c08008b0",
X"38029f05",
X"33028405",
X"9e053371",
X"982b7190",
X"2b07028c",
X"059d0533",
X"70882b72",
X"078d3d33",
X"7180ffff",
X"fe800607",
X"51525357",
X"58568339",
X"81557483",
X"c0800c89",
X"3d0d04fb",
X"3d0d83c0",
X"9008fe19",
X"881208fe",
X"05555654",
X"80567473",
X"278d3882",
X"14337571",
X"29941608",
X"05575375",
X"83c0800c",
X"873d0d04",
X"fc3d0d76",
X"52800b83",
X"c0900870",
X"33515253",
X"70832e09",
X"81069138",
X"95123394",
X"13337198",
X"2b71902b",
X"07555551",
X"9b12339a",
X"13337188",
X"2b077407",
X"83c0800c",
X"55863d0d",
X"04fc3d0d",
X"7683c090",
X"08555580",
X"75238815",
X"08537281",
X"2e883888",
X"14087326",
X"85388152",
X"b2397290",
X"38733352",
X"71832e09",
X"81068538",
X"90140853",
X"728c160c",
X"72802e8d",
X"387251fe",
X"d63f83c0",
X"80085285",
X"39901408",
X"52719016",
X"0c805271",
X"83c0800c",
X"863d0d04",
X"fa3d0d78",
X"83c09008",
X"71228105",
X"7083ffff",
X"06575457",
X"5573802e",
X"88389015",
X"08537286",
X"38835280",
X"e739738f",
X"06527180",
X"da388113",
X"90160c8c",
X"15085372",
X"9038830b",
X"84172257",
X"52737627",
X"80c638bf",
X"39821633",
X"ff057484",
X"2a065271",
X"b2387251",
X"fcb13f81",
X"527183c0",
X"800827a8",
X"38835283",
X"c0800888",
X"1708279c",
X"3883c080",
X"088c160c",
X"83c08008",
X"51fdbc3f",
X"83c08008",
X"90160c73",
X"75238052",
X"7183c080",
X"0c883d0d",
X"04f23d0d",
X"60626458",
X"5e5b7533",
X"5574a02e",
X"09810688",
X"38811670",
X"4456ef39",
X"62703356",
X"5674af2e",
X"09810684",
X"38811643",
X"800b881c",
X"0c627033",
X"5155749f",
X"2691387a",
X"51fdd23f",
X"83c08008",
X"56807d34",
X"83813993",
X"3d841c08",
X"7058595f",
X"8a55a076",
X"70810558",
X"34ff1555",
X"74ff2e09",
X"8106ef38",
X"80705a5c",
X"887f085f",
X"5a7b811d",
X"7081ff06",
X"60137033",
X"70af3270",
X"30a07327",
X"71802507",
X"5151525b",
X"535e5755",
X"7480e738",
X"76ae2e09",
X"81068338",
X"8155787a",
X"27750755",
X"74802e9f",
X"38798832",
X"703078ae",
X"32703070",
X"73079f2a",
X"53515751",
X"5675bb38",
X"88598b5a",
X"ffab3976",
X"982b5574",
X"80258738",
X"81ea8c17",
X"3357ff9f",
X"17557499",
X"268938e0",
X"177081ff",
X"06585578",
X"811a7081",
X"ff06721b",
X"535b5755",
X"767534fe",
X"f8397b1e",
X"7f0c8055",
X"76a02683",
X"38815574",
X"8b19347a",
X"51fc823f",
X"83c08008",
X"80f538a0",
X"547a2270",
X"852b83e0",
X"06545590",
X"1b08527c",
X"51a4923f",
X"83c08008",
X"5783c080",
X"08818138",
X"7c335574",
X"802e80f4",
X"388b1d33",
X"70832a70",
X"81065156",
X"5674b438",
X"8b7d841d",
X"0883c080",
X"08595b5b",
X"58ff1858",
X"77ff2e9a",
X"38797081",
X"055b3379",
X"7081055b",
X"33717131",
X"52565675",
X"802ee238",
X"86397580",
X"2e96387a",
X"51fbe53f",
X"ff863983",
X"c0800856",
X"83c08008",
X"b6388339",
X"7656841b",
X"088b1133",
X"515574a7",
X"388b1d33",
X"70842a70",
X"81065156",
X"56748938",
X"83569439",
X"81569039",
X"7c51fa94",
X"3f83c080",
X"08881c0c",
X"fd813975",
X"83c0800c",
X"903d0d04",
X"f83d0d7a",
X"7c595782",
X"5483fe53",
X"77527651",
X"a2d73f83",
X"5683c080",
X"0880ec38",
X"81173377",
X"3371882b",
X"07565682",
X"567482d4",
X"d52e0981",
X"0680d438",
X"7554b653",
X"77527651",
X"a2ab3f83",
X"c0800898",
X"38811733",
X"77337188",
X"2b0783c0",
X"80085256",
X"56748182",
X"c62eac38",
X"825480d2",
X"53775276",
X"51a2823f",
X"83c08008",
X"98388117",
X"33773371",
X"882b0783",
X"c0800852",
X"56567481",
X"82c62e83",
X"38815675",
X"83c0800c",
X"8a3d0d04",
X"eb3d0d67",
X"5a800b83",
X"c0900ca1",
X"a43f83c0",
X"80088106",
X"55825674",
X"83ef3874",
X"75538f3d",
X"70535759",
X"feca3f83",
X"c0800881",
X"ff065776",
X"812e0981",
X"0680d438",
X"905483be",
X"53745275",
X"51a1963f",
X"83c08008",
X"80c9388f",
X"3d335574",
X"802e80c9",
X"3802bf05",
X"33028405",
X"be053371",
X"982b7190",
X"2b07028c",
X"05bd0533",
X"70882b72",
X"07953d33",
X"71077058",
X"7b575e52",
X"5e575957",
X"fdee3f83",
X"c0800881",
X"ff065776",
X"832e0981",
X"06863881",
X"5682f239",
X"76802e86",
X"38865682",
X"e839a454",
X"8d537852",
X"7551a0ad",
X"3f815683",
X"c0800882",
X"d43802be",
X"05330284",
X"05bd0533",
X"71882b07",
X"595d77ab",
X"380280ce",
X"05330284",
X"0580cd05",
X"3371982b",
X"71902b07",
X"973d3370",
X"882b7207",
X"02940580",
X"cb053371",
X"0754525e",
X"57595602",
X"b7053378",
X"71290288",
X"05b60533",
X"028c05b5",
X"05337188",
X"2b07701d",
X"707f8c05",
X"0c5f5957",
X"595d8e3d",
X"33821b34",
X"02b90533",
X"903d3371",
X"882b075a",
X"5c78841b",
X"2302bb05",
X"33028405",
X"ba053371",
X"882b0756",
X"5c74ab38",
X"0280ca05",
X"33028405",
X"80c90533",
X"71982b71",
X"902b0796",
X"3d337088",
X"2b720702",
X"940580c7",
X"05337107",
X"51525357",
X"5e5c7476",
X"31783179",
X"842a903d",
X"33547171",
X"31535656",
X"80d6b33f",
X"83c08008",
X"82057088",
X"1c0c83c0",
X"8008e08a",
X"05565674",
X"83dffe26",
X"83388257",
X"83fff676",
X"27853883",
X"57893986",
X"5676802e",
X"80db3876",
X"7a347683",
X"2e098106",
X"b0380280",
X"d6053302",
X"840580d5",
X"05337198",
X"2b71902b",
X"07993d33",
X"70882b72",
X"07029405",
X"80d30533",
X"71077f90",
X"050c525e",
X"57585686",
X"39771b90",
X"1b0c841a",
X"228c1b08",
X"1971842a",
X"05941c0c",
X"5d800b81",
X"1b347983",
X"c0900c80",
X"567583c0",
X"800c973d",
X"0d04e93d",
X"0d83c090",
X"08568554",
X"75802e81",
X"8238800b",
X"81173499",
X"3de01146",
X"6a548a3d",
X"705458ec",
X"0551f6e5",
X"3f83c080",
X"085483c0",
X"800880df",
X"38893d33",
X"5473802e",
X"913802ab",
X"05337084",
X"2a810651",
X"5574802e",
X"86388354",
X"80c13976",
X"51f4893f",
X"83c08008",
X"a0170c02",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"9c1c0c52",
X"78981b0c",
X"53565957",
X"810b8117",
X"34745473",
X"83c0800c",
X"993d0d04",
X"f53d0d7d",
X"7f617283",
X"c090085a",
X"5d5d595c",
X"807b0c85",
X"5775802e",
X"81e03881",
X"16338106",
X"55845774",
X"802e81d2",
X"38913974",
X"81173486",
X"39800b81",
X"17348157",
X"81c0399c",
X"16089817",
X"08315574",
X"78278338",
X"74587780",
X"2e81a938",
X"98160870",
X"83ff0656",
X"577480cf",
X"38821633",
X"ff057789",
X"2a067081",
X"ff065a55",
X"78a03876",
X"8738a016",
X"08558d39",
X"a4160851",
X"f0e93f83",
X"c0800855",
X"817527ff",
X"a83874a4",
X"170ca416",
X"0851f283",
X"3f83c080",
X"085583c0",
X"8008802e",
X"ff893883",
X"c0800819",
X"a8170c98",
X"160883ff",
X"06848071",
X"31515577",
X"75278338",
X"77557483",
X"ffff0654",
X"98160883",
X"ff0653a8",
X"16085279",
X"577b8338",
X"7b577651",
X"9ad33f83",
X"c08008fe",
X"d0389816",
X"08159817",
X"0c741a78",
X"76317c08",
X"177d0c59",
X"5afed339",
X"80577683",
X"c0800c8d",
X"3d0d04fa",
X"3d0d7883",
X"c0900855",
X"56855573",
X"802e81e3",
X"38811433",
X"81065384",
X"5572802e",
X"81d5389c",
X"14085372",
X"76278338",
X"72569814",
X"0857800b",
X"98150c75",
X"802e81b9",
X"38821433",
X"70892b56",
X"5376802e",
X"b7387452",
X"ff165180",
X"d1b43f83",
X"c08008ff",
X"18765470",
X"53585380",
X"d1a43f83",
X"c0800873",
X"26963874",
X"30707806",
X"7098170c",
X"777131a4",
X"17085258",
X"51538939",
X"a0140870",
X"a4160c53",
X"747627b9",
X"387251ee",
X"d63f83c0",
X"80085381",
X"0b83c080",
X"08278b38",
X"88140883",
X"c0800826",
X"8838800b",
X"811534b0",
X"3983c080",
X"08a4150c",
X"98140815",
X"98150c75",
X"753156c4",
X"39981408",
X"16709816",
X"0c735256",
X"efc53f83",
X"c080088c",
X"3883c080",
X"08811534",
X"81559439",
X"821433ff",
X"0576892a",
X"0683c080",
X"0805a815",
X"0c805574",
X"83c0800c",
X"883d0d04",
X"ef3d0d63",
X"56855583",
X"c0900880",
X"2e80d238",
X"933df405",
X"84170c64",
X"53883d70",
X"53765257",
X"f1cf3f83",
X"c0800855",
X"83c08008",
X"b438883d",
X"33547380",
X"2ea13802",
X"a7053370",
X"842a7081",
X"06515555",
X"83557380",
X"2e973876",
X"51eef53f",
X"83c08008",
X"88170c75",
X"51efa63f",
X"83c08008",
X"557483c0",
X"800c933d",
X"0d04e43d",
X"0d6ea13d",
X"08405e85",
X"5683c090",
X"08802e84",
X"85389e3d",
X"f405841f",
X"0c7e9838",
X"7d51eef5",
X"3f83c080",
X"085683ee",
X"39814181",
X"f6398341",
X"81f13993",
X"3d7f9605",
X"4159807f",
X"8295055e",
X"56756081",
X"ff053483",
X"41901e08",
X"762e81d3",
X"38a0547d",
X"2270852b",
X"83e00654",
X"58901e08",
X"52785196",
X"dc3f83c0",
X"80084183",
X"c08008ff",
X"b8387833",
X"5c7b802e",
X"ffb4388b",
X"193370bf",
X"06718106",
X"52435574",
X"802e80de",
X"387b81bf",
X"0655748f",
X"2480d338",
X"9a193355",
X"7480cb38",
X"f31d7058",
X"5d815675",
X"8b2e0981",
X"0685388e",
X"568b3975",
X"9a2e0981",
X"0683389c",
X"56751970",
X"70810552",
X"33713381",
X"1a821a5f",
X"5b525b55",
X"74863879",
X"77348539",
X"80df7734",
X"777b5757",
X"7aa02e09",
X"8106c038",
X"81567b81",
X"e5327030",
X"709f2a51",
X"51557bae",
X"2e933874",
X"802e8e38",
X"61832a70",
X"81065155",
X"74802e97",
X"387d51ed",
X"df3f83c0",
X"80084183",
X"c0800887",
X"38901e08",
X"feaf3880",
X"60347580",
X"2e88387c",
X"527f518e",
X"823f6080",
X"2e863880",
X"0b901f0c",
X"60566083",
X"2e853860",
X"81d03889",
X"1f57901e",
X"08802e81",
X"a8388056",
X"75197033",
X"515574a0",
X"2ea03874",
X"852e0981",
X"06843881",
X"e5557477",
X"70810559",
X"34811670",
X"81ff0657",
X"55877627",
X"d7388819",
X"335574a0",
X"2ea938ae",
X"77708105",
X"59348856",
X"75197033",
X"515574a0",
X"2e953874",
X"77708105",
X"59348116",
X"7081ff06",
X"57558a76",
X"27e2388b",
X"19337f88",
X"05349f19",
X"339e1a33",
X"71982b71",
X"902b079d",
X"1c337088",
X"2b72079c",
X"1e337107",
X"640c5299",
X"1d33981e",
X"3371882b",
X"07535153",
X"57595674",
X"7f840523",
X"97193396",
X"1a337188",
X"2b075656",
X"747f8605",
X"23807734",
X"7d51ebf0",
X"3f83c080",
X"08833270",
X"30707207",
X"9f2c83c0",
X"80080652",
X"5656961f",
X"3355748a",
X"38891f52",
X"961f518c",
X"8e3f7583",
X"c0800c9e",
X"3d0d04f4",
X"3d0d7e8f",
X"3dec1156",
X"56589053",
X"f0155277",
X"51e0d23f",
X"83c08008",
X"80d63878",
X"902e0981",
X"0680cd38",
X"02ab0533",
X"81f3f00b",
X"81f3f033",
X"5758568c",
X"3974762e",
X"8a388417",
X"70335657",
X"74f33876",
X"33705755",
X"74802eac",
X"38821722",
X"708a2b90",
X"3dec0556",
X"70555656",
X"96800a52",
X"7751e081",
X"3f83c080",
X"08863878",
X"752e8538",
X"80568539",
X"81173356",
X"7583c080",
X"0c8e3d0d",
X"04fc3d0d",
X"76705255",
X"8b953f83",
X"c0800815",
X"ff055473",
X"752e8e38",
X"73335372",
X"ae2e8638",
X"ff1454ef",
X"39775281",
X"14518aad",
X"3f83c080",
X"08307083",
X"c0800807",
X"802583c0",
X"800c5386",
X"3d0d04fc",
X"3d0d7670",
X"5255e6ee",
X"3f83c080",
X"08548153",
X"83c08008",
X"80c13874",
X"51e6b13f",
X"83c08008",
X"81f0a853",
X"83c08008",
X"5253ff91",
X"3f83c080",
X"08a13881",
X"f0ac5272",
X"51ff823f",
X"83c08008",
X"923881f0",
X"b0527251",
X"fef33f83",
X"c0800880",
X"2e833881",
X"54735372",
X"83c0800c",
X"863d0d04",
X"fd3d0d75",
X"705254e6",
X"8d3f8153",
X"83c08008",
X"98387351",
X"e5d63f83",
X"c3980852",
X"83c08008",
X"51feba3f",
X"83c08008",
X"537283c0",
X"800c853d",
X"0d04df3d",
X"0da43d08",
X"70525edb",
X"f43f83c0",
X"80083395",
X"3d565473",
X"963881f7",
X"c0527451",
X"898d3f9a",
X"397d5278",
X"51defc3f",
X"84d0397d",
X"51dbda3f",
X"83c08008",
X"527451db",
X"8a3f8043",
X"80428041",
X"804083c3",
X"a0085294",
X"3d70525d",
X"e1e43f83",
X"c0800859",
X"800b83c0",
X"8008555b",
X"83c08008",
X"7b2e9438",
X"811b7452",
X"5be4e63f",
X"83c08008",
X"5483c080",
X"08ee3880",
X"5aff5f79",
X"09709f2c",
X"7b065b54",
X"7a7a2484",
X"38ff1b5a",
X"f61a7009",
X"709f2c72",
X"067bff12",
X"5a5a5255",
X"55807525",
X"95387651",
X"e4ab3f83",
X"c0800876",
X"ff185855",
X"57738024",
X"ed38747f",
X"2e8638a1",
X"b53f745f",
X"78ff1b70",
X"585d5880",
X"7a259538",
X"7751e481",
X"3f83c080",
X"0876ff18",
X"58555873",
X"8024ed38",
X"800b83c7",
X"d00c800b",
X"83c8980c",
X"81f0b451",
X"8d8c3f81",
X"800b83c8",
X"980c81f0",
X"bc518cfe",
X"3fa80b83",
X"c7d00c76",
X"802e80e4",
X"3883c7d0",
X"08777932",
X"70307072",
X"07802570",
X"872b83c8",
X"980c5156",
X"78535656",
X"e3b83f83",
X"c0800880",
X"2e883881",
X"f0c4518c",
X"c53f7651",
X"e2fa3f83",
X"c0800852",
X"81f2a451",
X"8cb43f76",
X"51e3823f",
X"83c08008",
X"83c7d008",
X"55577574",
X"258638a8",
X"1656f739",
X"7583c7d0",
X"0c86f076",
X"24ff9838",
X"87980b83",
X"c7d00c77",
X"802eb138",
X"7751e2b8",
X"3f83c080",
X"08785255",
X"e2d83f81",
X"f0cc5483",
X"c080088d",
X"38873980",
X"763481d0",
X"3981f0c8",
X"54745373",
X"5281f09c",
X"518bd33f",
X"805481f0",
X"a4518bca",
X"3f811454",
X"73a82e09",
X"8106ef38",
X"868da051",
X"9da83f80",
X"52903d70",
X"525780c7",
X"a93f8352",
X"765180c7",
X"a13f6281",
X"8f386180",
X"2e80fb38",
X"7b5473ff",
X"2e963878",
X"802e818a",
X"387851e1",
X"dc3f83c0",
X"8008ff15",
X"5559e739",
X"78802e80",
X"f5387851",
X"e1d83f83",
X"c0800880",
X"2efc8e38",
X"7851e1a0",
X"3f83c080",
X"085281f0",
X"985183e0",
X"3f83c080",
X"08a3387c",
X"5185983f",
X"83c08008",
X"5574ff16",
X"56548074",
X"25ae3874",
X"1d703355",
X"5673af2e",
X"fecd38e9",
X"397851e0",
X"e13f83c0",
X"8008527c",
X"5184d03f",
X"8f397f88",
X"29601005",
X"7a056105",
X"5afc9039",
X"62802efb",
X"d1388052",
X"765180c6",
X"813fa33d",
X"0d04803d",
X"0d9088b8",
X"337081ff",
X"0670842a",
X"81327081",
X"06515151",
X"5170802e",
X"8d38a80b",
X"9088b834",
X"b80b9088",
X"b8347083",
X"c0800c82",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067085",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d3898",
X"0b9088b8",
X"34b80b90",
X"88b83470",
X"83c0800c",
X"823d0d04",
X"930b9088",
X"bc34ff0b",
X"9088a834",
X"04ff3d0d",
X"028f0533",
X"52800b90",
X"88bc348a",
X"519aef3f",
X"df3f80f8",
X"0b9088a0",
X"34800b90",
X"888834fa",
X"12527190",
X"88803480",
X"0b908898",
X"34719088",
X"90349088",
X"b8528072",
X"34b87234",
X"833d0d04",
X"803d0d02",
X"8b053351",
X"709088b4",
X"34febf3f",
X"83c08008",
X"802ef638",
X"823d0d04",
X"803d0d84",
X"39a8de3f",
X"fed93f83",
X"c0800880",
X"2ef33890",
X"88b43370",
X"81ff0683",
X"c0800c51",
X"823d0d04",
X"803d0da3",
X"0b9088bc",
X"34ff0b90",
X"88a83490",
X"88b851a8",
X"7134b871",
X"34823d0d",
X"04803d0d",
X"9088bc33",
X"70982b70",
X"802583c0",
X"800c5151",
X"823d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"832a8132",
X"70810651",
X"51515170",
X"802ee838",
X"b00b9088",
X"b834b80b",
X"9088b834",
X"823d0d04",
X"803d0d90",
X"80ac0881",
X"0683c080",
X"0c823d0d",
X"04fd3d0d",
X"75775454",
X"80732594",
X"38737081",
X"05553352",
X"81f0d051",
X"87843fff",
X"1353e939",
X"853d0d04",
X"fd3d0d75",
X"77535473",
X"33517089",
X"38713351",
X"70802ea1",
X"38733372",
X"33525372",
X"71278538",
X"ff519439",
X"70732785",
X"3881518b",
X"39811481",
X"135354d3",
X"39805170",
X"83c0800c",
X"853d0d04",
X"fd3d0d75",
X"77545472",
X"337081ff",
X"06525270",
X"802ea338",
X"7181ff06",
X"8114ffbf",
X"12535452",
X"70992689",
X"38a01270",
X"81ff0653",
X"51717470",
X"81055634",
X"d2398074",
X"34853d0d",
X"04ffbd3d",
X"0d80c63d",
X"0852a53d",
X"705254ff",
X"b33f80c7",
X"3d085285",
X"3d705253",
X"ffa63f72",
X"527351fe",
X"df3f80c5",
X"3d0d04fe",
X"3d0d7476",
X"53537170",
X"81055333",
X"51707370",
X"81055534",
X"70f03884",
X"3d0d04fe",
X"3d0d7452",
X"80723352",
X"5370732e",
X"8d388112",
X"81147133",
X"53545270",
X"f5387283",
X"c0800c84",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"be8c3f83",
X"c080087a",
X"27ee3874",
X"802e80dd",
X"38745275",
X"51bdf73f",
X"83c08008",
X"75537652",
X"54bdfb3f",
X"83c08008",
X"7a537552",
X"56bddf3f",
X"83c08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"c08008c5",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9f",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fc813f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd53f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbb13f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83c0940c",
X"7183c098",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383c094",
X"085283c0",
X"980851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"bdbe5351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fc3d",
X"0d765574",
X"83c3ac08",
X"2eaf3880",
X"53745187",
X"c13f83c0",
X"800881ff",
X"06ff1470",
X"81ff0672",
X"30709f2a",
X"51525553",
X"5472802e",
X"843871dd",
X"3873fe38",
X"7483c3ac",
X"0c863d0d",
X"04ff3d0d",
X"ff0b83c3",
X"ac0c84a5",
X"3f815187",
X"853f83c0",
X"800881ff",
X"065271ee",
X"3881d33f",
X"7183c080",
X"0c833d0d",
X"04fc3d0d",
X"76028405",
X"a2052202",
X"8805a605",
X"227a5455",
X"5555ff82",
X"3f72802e",
X"a03883c3",
X"c0143375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552dd",
X"39800b83",
X"c0800c86",
X"3d0d04fc",
X"3d0d7678",
X"7a115653",
X"55805371",
X"742e9338",
X"72155170",
X"3383c3c0",
X"13348112",
X"81145452",
X"ea39800b",
X"83c0800c",
X"863d0d04",
X"fd3d0d90",
X"5483c3ac",
X"085186f4",
X"3f83c080",
X"0881ff06",
X"ff157130",
X"71307073",
X"079f2a72",
X"9f2a0652",
X"55525553",
X"72db3885",
X"3d0d0480",
X"3d0d83c3",
X"b8081083",
X"c3b00807",
X"9080a80c",
X"823d0d04",
X"800b83c3",
X"b80ce43f",
X"04810b83",
X"c3b80cdb",
X"3f04ed3f",
X"047183c3",
X"b40c0480",
X"3d0d8051",
X"f43f810b",
X"83c3b80c",
X"810b83c3",
X"b00cffbb",
X"3f823d0d",
X"04803d0d",
X"72307074",
X"07802583",
X"c3b00c51",
X"ffa53f82",
X"3d0d0480",
X"3d0d028b",
X"05339080",
X"a40c9080",
X"a8087081",
X"06515170",
X"f5389080",
X"a4087081",
X"ff0683c0",
X"800c5182",
X"3d0d0480",
X"3d0d81ff",
X"51d13f83",
X"c0800881",
X"ff0683c0",
X"800c823d",
X"0d04803d",
X"0d73902b",
X"73079080",
X"b40c823d",
X"0d0404fb",
X"3d0d7802",
X"84059f05",
X"3370982b",
X"55575572",
X"80259b38",
X"7580ff06",
X"56805280",
X"f751e03f",
X"83c08008",
X"81ff0654",
X"73812680",
X"ff388051",
X"fee73fff",
X"a23f8151",
X"fedf3fff",
X"9a3f7551",
X"feed3f74",
X"982a51fe",
X"e63f7490",
X"2a7081ff",
X"065253fe",
X"da3f7488",
X"2a7081ff",
X"065253fe",
X"ce3f7481",
X"ff0651fe",
X"c63f8155",
X"7580c02e",
X"09810686",
X"38819555",
X"8d397580",
X"c82e0981",
X"06843881",
X"87557451",
X"fea53f8a",
X"55fec83f",
X"83c08008",
X"81ff0670",
X"982b5454",
X"7280258c",
X"38ff1570",
X"81ff0656",
X"5374e238",
X"7383c080",
X"0c873d0d",
X"04fa3d0d",
X"fdc53f80",
X"51fdda3f",
X"8a54fe93",
X"3fff1470",
X"81ff0655",
X"5373f338",
X"73745355",
X"80c051fe",
X"a63f83c0",
X"800881ff",
X"06547381",
X"2e098106",
X"829f3883",
X"aa5280c8",
X"51fe8c3f",
X"83c08008",
X"81ff0653",
X"72812e09",
X"810681a8",
X"38745487",
X"3d741154",
X"56fdc83f",
X"83c08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e53802",
X"9a053353",
X"72812e09",
X"810681d9",
X"38029b05",
X"335380ce",
X"90547281",
X"aa2e8d38",
X"81c73980",
X"e4518b9a",
X"3fff1454",
X"73802e81",
X"b838820a",
X"5281e951",
X"fda53f83",
X"c0800881",
X"ff065372",
X"de387252",
X"80fa51fd",
X"923f83c0",
X"800881ff",
X"06537281",
X"90387254",
X"731653fc",
X"d63f83c0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e8",
X"38873d33",
X"70862a70",
X"81065154",
X"548c5572",
X"80e33884",
X"5580de39",
X"745281e9",
X"51fccc3f",
X"83c08008",
X"81ff0653",
X"825581e9",
X"56817327",
X"86387355",
X"80c15680",
X"ce90548a",
X"3980e451",
X"8a8c3fff",
X"14547380",
X"2ea93880",
X"527551fc",
X"9a3f83c0",
X"800881ff",
X"065372e1",
X"38848052",
X"80d051fc",
X"863f83c0",
X"800881ff",
X"06537280",
X"2e833880",
X"557483c3",
X"bc348051",
X"fb873ffb",
X"c23f883d",
X"0d04fb3d",
X"0d775480",
X"0b83c3bc",
X"3370832a",
X"70810651",
X"55575572",
X"752e0981",
X"06853873",
X"892b5473",
X"5280d151",
X"fbbd3f83",
X"c0800881",
X"ff065372",
X"bd3882b8",
X"c054fb83",
X"3f83c080",
X"0881ff06",
X"537281ff",
X"2e098106",
X"8938ff14",
X"5473e738",
X"9f397281",
X"fe2e0981",
X"06963883",
X"c7c05283",
X"c3c051fa",
X"ed3ffad3",
X"3ffad03f",
X"83398155",
X"8051fa89",
X"3ffac43f",
X"7481ff06",
X"83c0800c",
X"873d0d04",
X"fb3d0d77",
X"83c3c056",
X"548151f9",
X"ec3f83c3",
X"bc337083",
X"2a708106",
X"51545672",
X"85387389",
X"2b547352",
X"80d851fa",
X"b63f83c0",
X"800881ff",
X"06537280",
X"e43881ff",
X"51f9d43f",
X"81fe51f9",
X"ce3f8480",
X"53747081",
X"05563351",
X"f9c13fff",
X"137083ff",
X"ff065153",
X"72eb3872",
X"51f9b03f",
X"7251f9ab",
X"3ff9d03f",
X"83c08008",
X"9f0653a7",
X"88547285",
X"2e8c3899",
X"3980e451",
X"87c43fff",
X"1454f9b3",
X"3f83c080",
X"0881ff2e",
X"843873e9",
X"388051f8",
X"e43ff99f",
X"3f800b83",
X"c0800c87",
X"3d0d0471",
X"83c7c40c",
X"8880800b",
X"83c7c00c",
X"8480800b",
X"83c7c80c",
X"04fd3d0d",
X"77701755",
X"7705ff1a",
X"535371ff",
X"2e943873",
X"70810555",
X"33517073",
X"70810555",
X"34ff1252",
X"e939853d",
X"0d04fb3d",
X"0d87a681",
X"0b83c7c4",
X"08565675",
X"3383a680",
X"1634a054",
X"83a08053",
X"83c7c408",
X"5283c7c0",
X"0851ffb1",
X"3fa05483",
X"a4805383",
X"c7c40852",
X"83c7c008",
X"51ff9e3f",
X"905483a8",
X"805383c7",
X"c4085283",
X"c7c00851",
X"ff8b3fa0",
X"53805283",
X"c7c80883",
X"a0800551",
X"86953fa0",
X"53805283",
X"c7c80883",
X"a4800551",
X"86853f90",
X"53805283",
X"c7c80883",
X"a8800551",
X"85f53fff",
X"763483a0",
X"80548053",
X"83c7c408",
X"5283c7c8",
X"0851fec5",
X"3f80d080",
X"5483b080",
X"5383c7c4",
X"085283c7",
X"c80851fe",
X"b03f87ba",
X"3fa25480",
X"5383c7c8",
X"088c8005",
X"5281f4e4",
X"51fe9a3f",
X"860b87a8",
X"8334800b",
X"87a88234",
X"800b87a0",
X"9a34af0b",
X"87a09634",
X"bf0b87a0",
X"9734800b",
X"87a09834",
X"9f0b87a0",
X"9934800b",
X"87a09b34",
X"e00b87a8",
X"8934a20b",
X"87a88034",
X"830b87a4",
X"8f34820b",
X"87a88134",
X"873d0d04",
X"fc3d0d83",
X"a0805480",
X"5383c7c8",
X"085283c7",
X"c40851fd",
X"b83f80d0",
X"805483b0",
X"805383c7",
X"c8085283",
X"c7c40851",
X"fda33fa0",
X"5483a080",
X"5383c7c8",
X"085283c7",
X"c40851fd",
X"903fa054",
X"83a48053",
X"83c7c808",
X"5283c7c4",
X"0851fcfd",
X"3f905483",
X"a8805383",
X"c7c80852",
X"83c7c408",
X"51fcea3f",
X"83c7c408",
X"5583a680",
X"153387a6",
X"8134863d",
X"0d04fa3d",
X"0d787052",
X"55c1e33f",
X"83ffff0b",
X"83c08008",
X"25a93874",
X"51c1e43f",
X"83c08008",
X"9e3883c0",
X"80085788",
X"3dfc0554",
X"84808053",
X"83c7c408",
X"527451ff",
X"bf963fff",
X"bedc3f88",
X"3d0d04fa",
X"3d0d7870",
X"5255c1a2",
X"3f83ffff",
X"0b83c080",
X"08259638",
X"8057883d",
X"fc055484",
X"80805383",
X"c7c40852",
X"7451c095",
X"3f883d0d",
X"04803d0d",
X"90809008",
X"810683c0",
X"800c823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087081",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fd0676",
X"1007720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870822c",
X"bf0683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe830676",
X"822b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087088",
X"2c870683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f1ff06",
X"76882b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"912cbf06",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fc87",
X"ffff0676",
X"912b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087099",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70ffbf0a",
X"0676992b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90808008",
X"70882c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"0870892c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708a",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8b2c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708c2cbf",
X"0683c080",
X"0c51823d",
X"0d04fe3d",
X"0d7481e6",
X"29872a90",
X"80a00c84",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70810554",
X"34ff1151",
X"f039843d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"8405540c",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"84808053",
X"80528880",
X"0a51ffb3",
X"3f818080",
X"53805282",
X"800a51c6",
X"3f843d0d",
X"04803d0d",
X"8151fcaa",
X"3f72802e",
X"90388051",
X"fdfe3fcd",
X"3f83c7cc",
X"3351fdf4",
X"3f8151fc",
X"bb3f8051",
X"fcb63f80",
X"51fc873f",
X"823d0d04",
X"fd3d0d75",
X"52805480",
X"ff722588",
X"38810bff",
X"80135354",
X"ffbf1251",
X"70992686",
X"38e01252",
X"b039ff9f",
X"12519971",
X"27a738d0",
X"12e01354",
X"51708926",
X"85387252",
X"9839728f",
X"26853872",
X"528f3971",
X"ba2e0981",
X"0685389a",
X"52833980",
X"5273802e",
X"85388180",
X"12527181",
X"ff0683c0",
X"800c853d",
X"0d04803d",
X"0d84d8c0",
X"51807170",
X"81055334",
X"7084e0c0",
X"2e098106",
X"f038823d",
X"0d04fe3d",
X"0d029705",
X"3351fef4",
X"3f83c080",
X"0881ff06",
X"83c7d008",
X"54528073",
X"249b3883",
X"c8940813",
X"7283c898",
X"08075353",
X"71733483",
X"c7d00881",
X"0583c7d0",
X"0c843d0d",
X"04fa3d0d",
X"82800a1b",
X"55805788",
X"3dfc0554",
X"79537452",
X"7851ffba",
X"ac3f883d",
X"0d04fe3d",
X"0d83c7e8",
X"08527451",
X"c1903f83",
X"c080088c",
X"38765375",
X"5283c7e8",
X"0851c63f",
X"843d0d04",
X"fe3d0d83",
X"c7e80853",
X"75527451",
X"ffbbce3f",
X"83c08008",
X"8d387753",
X"765283c7",
X"e80851ff",
X"a03f843d",
X"0d04f73d",
X"0daaaa3f",
X"83c08008",
X"81ff06ff",
X"05577683",
X"38815780",
X"feec3f83",
X"c0800883",
X"c0800856",
X"5a871533",
X"5473802e",
X"80df3874",
X"0881ecb8",
X"2e098106",
X"80d33880",
X"0b911633",
X"55597379",
X"2e80c638",
X"74569a16",
X"33547383",
X"2e098106",
X"a438a416",
X"70335558",
X"80527351",
X"a8943f80",
X"53805273",
X"51a8b43f",
X"81145476",
X"74258338",
X"80547378",
X"34811980",
X"d8179117",
X"33565759",
X"78742e09",
X"8106ffbe",
X"3881c415",
X"98c01b55",
X"5574742e",
X"098106ff",
X"88388b3d",
X"0d04f63d",
X"0d80fdde",
X"3f83c080",
X"087d83c0",
X"80085859",
X"5b7783c7",
X"d00c8716",
X"33557480",
X"2e81a738",
X"75085473",
X"81eff02e",
X"09810693",
X"38901633",
X"53871633",
X"5281f0d8",
X"51e8f33f",
X"81883973",
X"81ecb82e",
X"09810680",
X"fd387452",
X"81f0ec51",
X"e8dc3f80",
X"70911833",
X"565b5973",
X"792e80e6",
X"38a41657",
X"f6173355",
X"79802e91",
X"38ff1554",
X"73822689",
X"38a81870",
X"83c7d00c",
X"5874812e",
X"09810687",
X"3881f0f4",
X"518d3974",
X"822e0981",
X"068a3881",
X"f0fc51e8",
X"953f9539",
X"74832e09",
X"81068f38",
X"76338105",
X"5281f188",
X"51e7ff3f",
X"815a8119",
X"80d81891",
X"18335658",
X"5978742e",
X"098106ff",
X"9f38a818",
X"81c41798",
X"c01d5657",
X"5875742e",
X"098106fe",
X"b8388c3d",
X"0d04fe3d",
X"0d83c7e8",
X"0851ffb7",
X"c13f83c0",
X"80088180",
X"802e0981",
X"06883883",
X"c1808053",
X"9c3983c7",
X"e80851ff",
X"b7a43f83",
X"c0800880",
X"d0802e09",
X"81069338",
X"83c1b080",
X"5383c080",
X"085283c7",
X"e80851fb",
X"d43f843d",
X"0d04803d",
X"0df6fc3f",
X"83c08008",
X"842981f5",
X"88057008",
X"83c0800c",
X"51823d0d",
X"04ed3d0d",
X"80448043",
X"80428041",
X"80705a5b",
X"facc3f80",
X"0b83c7d0",
X"0c800b83",
X"c8980c81",
X"f1dc51e6",
X"c53f8180",
X"0b83c898",
X"0c81f1e0",
X"51e6b73f",
X"80d00b83",
X"c7d00c78",
X"30707a07",
X"80257087",
X"2b83c898",
X"0c5155f5",
X"ed3f83c0",
X"80085281",
X"f1e851e6",
X"913f80f8",
X"0b83c7d0",
X"0c788132",
X"70307072",
X"07802570",
X"872b83c8",
X"980c5156",
X"569e9d3f",
X"83c08008",
X"5281f1f8",
X"51e5e73f",
X"81a00b83",
X"c7d00c78",
X"82327030",
X"70720780",
X"2570872b",
X"83c8980c",
X"515656fe",
X"c53f83c0",
X"80085281",
X"f28851e5",
X"bd3f81c8",
X"0b83c7d0",
X"0c788332",
X"70307072",
X"07802570",
X"872b83c8",
X"980c5156",
X"83c7e808",
X"5256ffb2",
X"983f83c0",
X"80085281",
X"f29051e5",
X"8d3f8298",
X"0b83c7d0",
X"0c810b83",
X"c7d45b58",
X"83c7d008",
X"83197a32",
X"70307072",
X"07802570",
X"872b83c8",
X"980c5157",
X"8e3d7055",
X"ff1b5457",
X"57579bdf",
X"3f797084",
X"055b0851",
X"ffb1ce3f",
X"745483c0",
X"80085377",
X"5281f298",
X"51e4bf3f",
X"a81783c7",
X"d00c8118",
X"5877852e",
X"098106ff",
X"af3883b8",
X"0b83c7d0",
X"0c788832",
X"70307072",
X"07802570",
X"872b83c8",
X"980c5156",
X"56f4b93f",
X"81f2a855",
X"83c08008",
X"802e8f38",
X"83c7e408",
X"51ffb0f9",
X"3f83c080",
X"08557452",
X"81f2b051",
X"e3ec3f83",
X"e00b83c7",
X"d00c7889",
X"32703070",
X"72078025",
X"70872b83",
X"c8980c51",
X"5681f2bc",
X"5256e3ca",
X"3f84b00b",
X"83c7d00c",
X"788a3270",
X"30707207",
X"80257087",
X"2b83c898",
X"0c515681",
X"f2d45256",
X"e3a83f80",
X"0b83c898",
X"0c858051",
X"f9ec3f86",
X"8da051f5",
X"853f8052",
X"913d7052",
X"559f873f",
X"83527451",
X"9f803f63",
X"557483a6",
X"38611959",
X"78802585",
X"38745990",
X"398a7925",
X"85388a59",
X"8739788a",
X"26838538",
X"78822b55",
X"81ec8c15",
X"0804f2a6",
X"3f83c080",
X"08615755",
X"75812e09",
X"81068938",
X"83c08008",
X"10559039",
X"75ff2e09",
X"81068838",
X"83c08008",
X"812c5590",
X"75258538",
X"90558839",
X"74802483",
X"38815574",
X"51f2803f",
X"82ba399a",
X"b63f83c0",
X"80086105",
X"55748025",
X"85388055",
X"88398775",
X"25833887",
X"5574518e",
X"983f8298",
X"39f1f03f",
X"83c08008",
X"61055574",
X"80258538",
X"80558839",
X"86752583",
X"38865574",
X"51f1e93f",
X"81f63960",
X"87386280",
X"2e81ed38",
X"83c39c08",
X"83c3980c",
X"adec0b83",
X"c3a00c83",
X"c7e80851",
X"d2b43ff9",
X"e13f81d0",
X"39605680",
X"76259838",
X"ad8b0b83",
X"c3a00c83",
X"c7c41570",
X"085255d2",
X"953f7408",
X"52923975",
X"80259238",
X"83c7c415",
X"0851ffae",
X"923f8052",
X"fc1951b8",
X"3962802e",
X"81963883",
X"c7c41570",
X"0883c7d4",
X"08720c83",
X"c7d40cfc",
X"1a705351",
X"558ce53f",
X"83c08008",
X"5680518c",
X"db3f83c0",
X"80085274",
X"5188f43f",
X"75528051",
X"88ed3f80",
X"df396055",
X"807525b6",
X"3883c3a8",
X"0883c398",
X"0cadec0b",
X"83c3a00c",
X"83c7e408",
X"51d19f3f",
X"83c7e408",
X"51cec03f",
X"83c08008",
X"81ff0670",
X"5255f0c9",
X"3f74802e",
X"a7388155",
X"ab397480",
X"259e3883",
X"c7e40851",
X"ffad843f",
X"8051f0ad",
X"3f8e3962",
X"802e8938",
X"f5943f84",
X"39628738",
X"7a802ef8",
X"ff388055",
X"7483c080",
X"0c953d0d",
X"04fe3d0d",
X"83c88451",
X"8183c43f",
X"83c7f451",
X"8183bc3f",
X"f0bf3f83",
X"c0800880",
X"2e863880",
X"51818a39",
X"f0c43f83",
X"c0800880",
X"fe38f0e4",
X"3f83c080",
X"08802eb9",
X"388151ee",
X"a13f8051",
X"effa3fea",
X"993f800b",
X"83c7d00c",
X"f8973f83",
X"c0800853",
X"ff0b83c7",
X"d00cec8c",
X"3f7280cb",
X"3883c7cc",
X"3351efd4",
X"3f7251ed",
X"f13f80c0",
X"39f08c3f",
X"83c08008",
X"802eb538",
X"8151edde",
X"3f8051ef",
X"b73fe9d6",
X"3fad8b0b",
X"83c3a00c",
X"83c7d408",
X"51cfb73f",
X"ff0b83c7",
X"d00cebc8",
X"3f83c7d4",
X"08528051",
X"86d13f81",
X"51f0fe3f",
X"843d0d04",
X"fb3d0d80",
X"5283c884",
X"5180f2cb",
X"3f815283",
X"c7f45180",
X"f2c13f80",
X"0b83c7cc",
X"34908080",
X"52868480",
X"8051ffaf",
X"963f83c0",
X"800881a0",
X"3883c7f0",
X"08518188",
X"f73f8a99",
X"3f81f7a8",
X"51ffb3cc",
X"3f83c080",
X"08559c80",
X"0a5480c0",
X"805381f2",
X"dc5283c0",
X"800851f2",
X"c73f83c7",
X"e8085381",
X"f2ec5274",
X"51ffae95",
X"3f83c080",
X"088438f5",
X"d53f83c7",
X"ec085381",
X"f2f85274",
X"51ffadfd",
X"3f83c080",
X"08b63887",
X"3dfc0554",
X"84808053",
X"86a88080",
X"5283c7ec",
X"0851ffac",
X"883f83c0",
X"80089338",
X"75848080",
X"2e098106",
X"8938810b",
X"83c7cc34",
X"8739800b",
X"83c7cc34",
X"83c7cc33",
X"51edc13f",
X"8151efad",
X"3f93cb3f",
X"8151efa5",
X"3f8151fc",
X"f43ffa39",
X"83c08c08",
X"0283c08c",
X"0cfb3d0d",
X"0281f384",
X"0b83c39c",
X"0c81f388",
X"0b83c394",
X"0c81f38c",
X"0b83c3a8",
X"0c81f390",
X"0b83c3a4",
X"0c83c08c",
X"08fc050c",
X"800b83c7",
X"d40b83c0",
X"8c08f805",
X"0c83c08c",
X"08f4050c",
X"ffac903f",
X"83c08008",
X"8605fc06",
X"83c08c08",
X"f0050c02",
X"83c08c08",
X"f0050831",
X"0d833d70",
X"83c08c08",
X"f8050870",
X"840583c0",
X"8c08f805",
X"0c0c51ff",
X"a8d13f83",
X"c08c08f4",
X"05088105",
X"83c08c08",
X"f4050c83",
X"c08c08f4",
X"0508882e",
X"098106ff",
X"ab388694",
X"808051e5",
X"ea3fff0b",
X"83c7d00c",
X"800b83c8",
X"980c84d8",
X"c00b83c8",
X"940c8151",
X"ea903f81",
X"51eab53f",
X"8051eab0",
X"3f8151ea",
X"d63f8251",
X"eafe3f80",
X"51eba63f",
X"8051ebd0",
X"3f80d1ae",
X"528051da",
X"ce3ffcbc",
X"3f83c08c",
X"08fc0508",
X"0d800b83",
X"c0800c87",
X"3d0d83c0",
X"8c0c0480",
X"3d0d81ff",
X"51800b83",
X"c8a81234",
X"ff115170",
X"f438823d",
X"0d04ff3d",
X"0d737033",
X"53518111",
X"33713471",
X"81123483",
X"3d0d04ff",
X"3d0d83ca",
X"c408a82e",
X"0981068b",
X"3883cadc",
X"0883cac4",
X"0c8739a8",
X"0b83cac4",
X"0c83cac4",
X"08860570",
X"81ff0652",
X"52d0d63f",
X"833d0d04",
X"fb3d0d77",
X"79565680",
X"70715555",
X"52717525",
X"ac387216",
X"70337014",
X"7081ff06",
X"55515151",
X"71742789",
X"38811270",
X"81ff0653",
X"51718114",
X"7083ffff",
X"06555254",
X"747324d6",
X"387183c0",
X"800c873d",
X"0d04fb3d",
X"0d775689",
X"39f9c63f",
X"8351eafe",
X"3fd1dd3f",
X"83c08008",
X"802eee38",
X"83cac408",
X"86057081",
X"ff065253",
X"cfe33f81",
X"0b9088d4",
X"34f99e3f",
X"8351ead6",
X"3f9088d4",
X"337081ff",
X"06555373",
X"802eea38",
X"73862a70",
X"81065153",
X"72ffbe38",
X"73982b53",
X"80732480",
X"de38d0cd",
X"3f83c080",
X"085583c0",
X"800880cf",
X"38741675",
X"822b5454",
X"9088c013",
X"33743481",
X"15557485",
X"2e098106",
X"e8387533",
X"83c8a834",
X"81163383",
X"c8a93482",
X"163383c8",
X"aa348316",
X"3383c8ab",
X"34845283",
X"c8a851fe",
X"933f83c0",
X"800881ff",
X"06841733",
X"55537274",
X"2e8738fd",
X"ce3ffed1",
X"3980e451",
X"e9c83f87",
X"3d0d04f4",
X"3d0d7e60",
X"5955805d",
X"8075822b",
X"7183cac8",
X"120c83ca",
X"e0175b5b",
X"57767934",
X"77772e83",
X"b7387652",
X"7751ffa6",
X"ec3f8e3d",
X"fc055490",
X"5383cab0",
X"527751ff",
X"a6a73f7c",
X"5675902e",
X"09810683",
X"933883ca",
X"b051fcde",
X"3f83cab2",
X"51fcd73f",
X"83cab451",
X"fcd03f76",
X"83cac00c",
X"7751ffa3",
X"ec3f81f0",
X"ac5283c0",
X"800851c6",
X"8c3f83c0",
X"8008812e",
X"09810680",
X"d4387683",
X"cad80c82",
X"0b83cab0",
X"34ff960b",
X"83cab134",
X"7751ffa6",
X"b93f83c0",
X"80085583",
X"c0800877",
X"25883883",
X"c080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583cab2",
X"347483ca",
X"b3347683",
X"cab434ff",
X"800b83ca",
X"b5348190",
X"3983cab0",
X"3383cab1",
X"3371882b",
X"07565b74",
X"83ffff2e",
X"09810680",
X"e838fe80",
X"0b83cad8",
X"0c810b83",
X"cac00cff",
X"0b83cab0",
X"34ff0b83",
X"cab13477",
X"51ffa5c6",
X"3f83c080",
X"0883cae4",
X"0c83c080",
X"085583c0",
X"80088025",
X"883883c0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83cab234",
X"7483cab3",
X"347683ca",
X"b434ff80",
X"0b83cab5",
X"34810b83",
X"cabf34a5",
X"39748596",
X"2e098106",
X"80fe3875",
X"83cad80c",
X"7751ffa4",
X"fa3f83ca",
X"bf3383c0",
X"80080755",
X"7483cabf",
X"3483cabf",
X"33810655",
X"74802e83",
X"38845783",
X"cab43383",
X"cab53371",
X"882b0756",
X"5c748180",
X"2e098106",
X"a13883ca",
X"b23383ca",
X"b3337188",
X"2b07565b",
X"ad807527",
X"87387682",
X"07579c39",
X"76810757",
X"96397482",
X"802e0981",
X"06873876",
X"83075787",
X"397481ff",
X"268a3877",
X"83cac81b",
X"0c767934",
X"8e3d0d04",
X"803d0d72",
X"842983ca",
X"c8057008",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"727083c8",
X"a00c7084",
X"2981f6dc",
X"05700883",
X"cadc0c51",
X"51823d0d",
X"04fe3d0d",
X"8151de3f",
X"800b83ca",
X"ac0c800b",
X"83caa80c",
X"ff0b83c8",
X"a40ca80b",
X"83cac40c",
X"ae51ca91",
X"3f800b83",
X"cac85452",
X"80737084",
X"05550c81",
X"12527184",
X"2e098106",
X"ef38843d",
X"0d04fe3d",
X"0d740284",
X"05960522",
X"53537180",
X"2e963872",
X"70810554",
X"3351ca9c",
X"3fff1270",
X"83ffff06",
X"5152e739",
X"843d0d04",
X"fe3d0d02",
X"92052253",
X"82ac51e4",
X"bd3f80c3",
X"51c9f93f",
X"819651e4",
X"b13f7252",
X"83c8a851",
X"ffb43f72",
X"5283c8a8",
X"51f8cd3f",
X"83c08008",
X"81ff0651",
X"c9d63f84",
X"3d0d04ff",
X"b13d0d80",
X"d13df805",
X"51f8f73f",
X"83caac08",
X"810583ca",
X"ac0c80cf",
X"3d33cf11",
X"7081ff06",
X"51565674",
X"832688e7",
X"38758f06",
X"ff055675",
X"83c8a408",
X"2e9b3875",
X"83269638",
X"7583c8a4",
X"0c758429",
X"83cac805",
X"70085355",
X"7551f9fb",
X"3f807624",
X"88c33875",
X"842983ca",
X"c8055574",
X"08802e88",
X"b43883c8",
X"a4088429",
X"83cac805",
X"70080288",
X"0582b905",
X"33525b55",
X"7480d22e",
X"84b03874",
X"80d22490",
X"3874bf2e",
X"9c387480",
X"d02e81d5",
X"3887f239",
X"7480d32e",
X"80d33874",
X"80d72e81",
X"c43887e1",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055656",
X"c8d23f80",
X"c151c88c",
X"3ff6983f",
X"83cadf33",
X"83c8a834",
X"815283c8",
X"a851c9a9",
X"3f8151fd",
X"e73f748b",
X"3883cadc",
X"0883cac4",
X"0c8739a8",
X"0b83cac4",
X"0cc89d3f",
X"80c151c7",
X"d73ff5e3",
X"3f900b83",
X"cabf3381",
X"06565674",
X"802e8338",
X"985683ca",
X"b43383ca",
X"b5337188",
X"2b075659",
X"7481802e",
X"0981069c",
X"3883cab2",
X"3383cab3",
X"3371882b",
X"075657ad",
X"8075278c",
X"38758180",
X"07568539",
X"75a00756",
X"7583c8a8",
X"34ff0b83",
X"c8a934e0",
X"0b83c8aa",
X"34800b83",
X"c8ab3484",
X"5283c8a8",
X"51c89e3f",
X"8451869b",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055659",
X"c7923f79",
X"51ff9fa7",
X"3f83c080",
X"08802e8a",
X"3880ce51",
X"c6be3f85",
X"f13980c1",
X"51c6b53f",
X"c7a63fc5",
X"df3f83ca",
X"d8085883",
X"75259b38",
X"83cab433",
X"83cab533",
X"71882b07",
X"fc177129",
X"7a058380",
X"055a5157",
X"8d397481",
X"802918ff",
X"80055881",
X"80578056",
X"76762e92",
X"38c6913f",
X"83c08008",
X"83c8a817",
X"34811656",
X"eb39c680",
X"3f83c080",
X"0881ff06",
X"775383c8",
X"a85256f4",
X"bf3f83c0",
X"800881ff",
X"06557575",
X"2e098106",
X"81953894",
X"51dffb3f",
X"c5fa3f80",
X"c151c5b4",
X"3fc6a53f",
X"77527951",
X"ff9dba3f",
X"805e80d1",
X"3dfdf405",
X"54765383",
X"c8a85279",
X"51ff9bc0",
X"3f0282b9",
X"05335581",
X"597480d7",
X"2e098106",
X"80c53877",
X"527951ff",
X"9d8b3f80",
X"d13dfdf0",
X"05547653",
X"8f3d7053",
X"7a5258ff",
X"9cc33f80",
X"5676762e",
X"a2387518",
X"83c8a817",
X"33713370",
X"72327030",
X"70802570",
X"307f0681",
X"1d5d5f51",
X"5151525b",
X"55db3982",
X"ac51def6",
X"3f78802e",
X"863880c3",
X"51843980",
X"ce51c4a8",
X"3fc5993f",
X"c3d23f83",
X"d8390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290559",
X"5580705d",
X"5980e451",
X"dec03fc4",
X"bf3f80c1",
X"51c3f93f",
X"83cac008",
X"792e82d6",
X"3883cae4",
X"0880fc05",
X"5580fd52",
X"745185c2",
X"3f83c080",
X"085b7782",
X"24b238ff",
X"1870872b",
X"83ffff80",
X"0681f5a8",
X"0583c8a8",
X"59575581",
X"80557570",
X"81055733",
X"77708105",
X"5934ff15",
X"7081ff06",
X"515574ea",
X"38828539",
X"7782e82e",
X"81a33877",
X"82e92e09",
X"810681aa",
X"38785877",
X"87327030",
X"70720780",
X"257a8a32",
X"70307072",
X"07802573",
X"0753545a",
X"51575575",
X"802e9738",
X"78782692",
X"38a00b83",
X"c8a81a34",
X"81197081",
X"ff065a55",
X"eb398118",
X"7081ff06",
X"59558a78",
X"27ffbc38",
X"8f5883c8",
X"a3183383",
X"c8a81934",
X"ff187081",
X"ff065955",
X"778426ea",
X"38905880",
X"0b83c8a8",
X"19348118",
X"7081ff06",
X"70982b52",
X"59557480",
X"25e93880",
X"c6557a85",
X"8f248438",
X"80c25574",
X"83c8a834",
X"80f10b83",
X"c8ab3481",
X"0b83c8ac",
X"347a83c8",
X"a9347a88",
X"2c557483",
X"c8aa3480",
X"cb3982f0",
X"782580c4",
X"387780fd",
X"29fd97d3",
X"05527951",
X"ff99e63f",
X"80d13dfd",
X"ec055480",
X"fd5383c8",
X"a8527951",
X"ff999e3f",
X"7b811959",
X"567580fc",
X"24833878",
X"5877882c",
X"557483c9",
X"a5347783",
X"c9a63475",
X"83c9a734",
X"81805980",
X"cc3983ca",
X"d8085783",
X"78259b38",
X"83cab433",
X"83cab533",
X"71882b07",
X"fc1a7129",
X"79058380",
X"05595159",
X"8d397781",
X"802917ff",
X"80055781",
X"80597652",
X"7951ff98",
X"f43f80d1",
X"3dfdec05",
X"54785383",
X"c8a85279",
X"51ff98ad",
X"3f7851f6",
X"bf3fc1bc",
X"3fffbff4",
X"3f8b3983",
X"caa80881",
X"0583caa8",
X"0c80d13d",
X"0d04f6df",
X"3ffc39fc",
X"3d0d7678",
X"71842983",
X"cac80570",
X"08515353",
X"53709e38",
X"80ce7234",
X"80cf0b81",
X"133480ce",
X"0b821334",
X"80c50b83",
X"13347084",
X"133480e7",
X"3983cae0",
X"13335480",
X"d2723473",
X"822a7081",
X"06515180",
X"cf537084",
X"3880d753",
X"72811334",
X"a00b8213",
X"34738306",
X"5170812e",
X"9e387081",
X"24883870",
X"802e8f38",
X"9f397082",
X"2e923870",
X"832e9238",
X"933980d8",
X"558e3980",
X"d3558939",
X"80cd5584",
X"3980c455",
X"74831334",
X"80c40b84",
X"1334800b",
X"85133486",
X"3d0d0483",
X"c8a00883",
X"c0800c04",
X"803d0d83",
X"c8a00884",
X"2981f6fc",
X"05700883",
X"c0800c51",
X"823d0d04",
X"fc3d0d76",
X"78535481",
X"53805587",
X"39711073",
X"10545273",
X"72265172",
X"802ea738",
X"70802e86",
X"38718025",
X"e8387280",
X"2e983871",
X"74268938",
X"73723175",
X"74075654",
X"72812a72",
X"812a5353",
X"e5397351",
X"78833874",
X"517083c0",
X"800c863d",
X"0d04fe3d",
X"0d805375",
X"527451ff",
X"a33f843d",
X"0d04fe3d",
X"0d815375",
X"527451ff",
X"933f843d",
X"0d04fb3d",
X"0d777955",
X"55805674",
X"76258638",
X"74305581",
X"56738025",
X"88387330",
X"76813257",
X"54805373",
X"527451fe",
X"e73f83c0",
X"80085475",
X"802e8738",
X"83c08008",
X"30547383",
X"c0800c87",
X"3d0d04fa",
X"3d0d787a",
X"57558057",
X"74772586",
X"38743055",
X"8157759f",
X"2c548153",
X"75743274",
X"31527451",
X"feaa3f83",
X"c0800854",
X"76802e87",
X"3883c080",
X"08305473",
X"83c0800c",
X"883d0d04",
X"fc3d0d76",
X"5580750c",
X"800b8416",
X"0c800b88",
X"160c800b",
X"8c160c83",
X"c8845180",
X"e9b13f83",
X"c7f45180",
X"e9a93f87",
X"a6803370",
X"81ff0670",
X"71842a06",
X"515152d6",
X"f03f7181",
X"2a813272",
X"81327181",
X"06718106",
X"3184180c",
X"54547183",
X"2a813272",
X"822a8132",
X"70810672",
X"7131780c",
X"51535387",
X"a0903387",
X"a0913370",
X"81ff0670",
X"73068132",
X"81068819",
X"0c515353",
X"83c08008",
X"802e80c2",
X"3883c080",
X"08812a70",
X"810683c0",
X"80088106",
X"3184170c",
X"5283c080",
X"08832a83",
X"c0800882",
X"2a718106",
X"71810631",
X"770c5353",
X"83c08008",
X"842a8106",
X"88160c83",
X"c0800885",
X"2a81068c",
X"160c863d",
X"0d04fe3d",
X"0d747654",
X"527151fe",
X"ab3f7281",
X"2ea23881",
X"73268d38",
X"72822ea8",
X"3872832e",
X"9c38e639",
X"7108e238",
X"841208dd",
X"38881208",
X"d838a539",
X"88120881",
X"2e9e3891",
X"39881208",
X"812e9538",
X"71089138",
X"8412088c",
X"388c1208",
X"812e0981",
X"06ffb238",
X"843d0d04",
X"fb3d0d78",
X"0284059f",
X"05335556",
X"800b81ee",
X"a4565381",
X"732b7406",
X"5271802e",
X"83388152",
X"74708205",
X"56227073",
X"902b0790",
X"809c0c51",
X"81135372",
X"882e0981",
X"06d93880",
X"5383caec",
X"13335170",
X"81ff2eb2",
X"38701081",
X"ecc40570",
X"22555180",
X"73177033",
X"701081ec",
X"c4057022",
X"51515152",
X"5273712e",
X"91388112",
X"5271862e",
X"098106f1",
X"38739080",
X"9c0c8113",
X"5372862e",
X"098106ff",
X"b8388053",
X"72167033",
X"51517081",
X"ff2e9438",
X"701081ec",
X"c4057022",
X"70848080",
X"0790809c",
X"0c515181",
X"13537286",
X"2e098106",
X"d7388053",
X"72165170",
X"3383caec",
X"14348113",
X"5372862e",
X"098106ec",
X"38873d0d",
X"0404fe3d",
X"0d750284",
X"05930533",
X"81065252",
X"70883871",
X"9080940c",
X"8e397081",
X"2e098106",
X"86387190",
X"80980c84",
X"3d0d04fb",
X"3d0d7898",
X"2b70982c",
X"7b982b70",
X"982c0290",
X"059f0533",
X"810683cb",
X"88117033",
X"70982b70",
X"982c5158",
X"5c5a5651",
X"55515470",
X"742e0981",
X"06943883",
X"cae81233",
X"70982b70",
X"982c5152",
X"5670732e",
X"b1387375",
X"347283ca",
X"e8133483",
X"cae93383",
X"cb893371",
X"982b7190",
X"2b0783ca",
X"e8337088",
X"2b720783",
X"cb883371",
X"079080b8",
X"0c525953",
X"5452873d",
X"0d04fe3d",
X"0d748111",
X"33713371",
X"882b0783",
X"c0800c53",
X"51843d0d",
X"0483caf4",
X"3383c080",
X"0c04f53d",
X"0d02bb05",
X"33028405",
X"bf053302",
X"880580c3",
X"0533028c",
X"0580c605",
X"22665c5a",
X"5e5c567a",
X"557b5489",
X"53a1527d",
X"5180df84",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8d3d0d04",
X"83c08c08",
X"0283c08c",
X"0cf53d0d",
X"83c08c08",
X"88050883",
X"c08c088f",
X"053383c0",
X"8c089205",
X"22028c05",
X"73900583",
X"c08c08e8",
X"050c83c0",
X"8c08f805",
X"0c83c08c",
X"08f0050c",
X"83c08c08",
X"ec050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"f0050883",
X"c08c08e0",
X"050c83c0",
X"8c08fc05",
X"0c83c08c",
X"08f00508",
X"89278a38",
X"890b83c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"860587ff",
X"fc0683c0",
X"8c08e005",
X"0c0283c0",
X"8c08e005",
X"08310d85",
X"3d705583",
X"c08c08ec",
X"05085483",
X"c08c08f0",
X"05085383",
X"c08c08f4",
X"05085283",
X"c08c08e4",
X"050c80e8",
X"dd3f83c0",
X"800881ff",
X"0683c08c",
X"08e40508",
X"83c08c08",
X"ec050c83",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08802e8c",
X"3883c08c",
X"08f80508",
X"0d89c839",
X"83c08c08",
X"f0050880",
X"2e89a638",
X"83c08c08",
X"ec050881",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"842ea938",
X"840b83c0",
X"8c08e005",
X"082588c7",
X"3883c08c",
X"08e00508",
X"852e859b",
X"3883c08c",
X"08e00508",
X"a12e87ad",
X"3888ac39",
X"800b83c0",
X"8c08ec05",
X"08850533",
X"83c08c08",
X"e0050c83",
X"c08c08fc",
X"050c83c0",
X"8c08e005",
X"08832e09",
X"81068883",
X"3883c08c",
X"08e80508",
X"81053383",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08812687",
X"e638810b",
X"83c08c08",
X"e0050880",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08fc050c",
X"83c08c08",
X"ec050882",
X"053383c0",
X"8c08e005",
X"08870534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088b0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08e005",
X"088c0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088d0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08e005",
X"088e0523",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088a0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"08057094",
X"0508fcff",
X"ff067194",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08ec0508",
X"86053383",
X"c08c08e0",
X"050c83c0",
X"8c08f405",
X"0c83c08c",
X"08e00508",
X"83c08c08",
X"fc05082e",
X"098106b6",
X"3883c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08fc0508",
X"83c08c08",
X"e005088b",
X"053483c0",
X"8c08ec05",
X"08870533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508812e",
X"8f3883c0",
X"8c08e005",
X"08822eb7",
X"38848c39",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"820b83c0",
X"8c08e005",
X"088a0534",
X"83d93983",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c83",
X"c08c08fc",
X"050883c0",
X"8c08e005",
X"088a0534",
X"83a13983",
X"c08c08fc",
X"0508802e",
X"83953883",
X"c08c08ec",
X"05088305",
X"33830683",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08832e09",
X"810682f3",
X"3883c08c",
X"08ec0508",
X"82053370",
X"982b83c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"83c08c08",
X"e0050880",
X"2582cc38",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"83c08c08",
X"ec050886",
X"053383c0",
X"8c08e005",
X"0880d605",
X"3483c08c",
X"08e00508",
X"840583c0",
X"8c08ec05",
X"08820533",
X"8f0683c0",
X"8c08e405",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"e4050883",
X"c08c08e0",
X"05083483",
X"c08c08ec",
X"05088405",
X"3383c08c",
X"08e00508",
X"81053480",
X"0b83c08c",
X"08e00508",
X"82053483",
X"c08c08e0",
X"050808ff",
X"83ff0682",
X"800783c0",
X"8c08e005",
X"080c83c0",
X"8c08e805",
X"08810533",
X"810583c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"83c08c08",
X"e8050881",
X"05348183",
X"3983c08c",
X"08fc0508",
X"802e80f7",
X"3883c08c",
X"08ec0508",
X"86053383",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08a22e09",
X"810680d7",
X"3883c08c",
X"08ec0508",
X"88053383",
X"c08c08ec",
X"05088705",
X"33718280",
X"290583c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c52",
X"83c08c08",
X"e4050c83",
X"c08c08f4",
X"050c83c0",
X"8c08e405",
X"0883c08c",
X"08e00508",
X"88052383",
X"c08c08ec",
X"05083383",
X"c08c08f0",
X"05087131",
X"7083ffff",
X"0683c08c",
X"08f0050c",
X"83c08c08",
X"e0050c83",
X"c08c08ec",
X"05080583",
X"c08c08ec",
X"050cf6d0",
X"3983c08c",
X"08f80508",
X"0d83c08c",
X"08f00508",
X"83c08c08",
X"e0050c83",
X"c08c08f8",
X"05080d83",
X"c08c08e0",
X"050883c0",
X"800c8d3d",
X"0d83c08c",
X"0c0483c0",
X"8c080283",
X"c08c0ce7",
X"3d0d83c0",
X"8c088805",
X"08028405",
X"83c08c08",
X"e8050c83",
X"c08c08d4",
X"050c800b",
X"83cb9034",
X"83c08c08",
X"d4050890",
X"0583c08c",
X"08c4050c",
X"800b83c0",
X"8c08c405",
X"0834800b",
X"83c08c08",
X"c4050881",
X"0534800b",
X"83c08c08",
X"c8050c83",
X"c08c08c8",
X"050880d8",
X"2983c08c",
X"08c40508",
X"0583c08c",
X"08ffb805",
X"0c800b83",
X"c08c08ff",
X"b8050880",
X"d8050c83",
X"c08c08ff",
X"b8050884",
X"0583c08c",
X"08ffb805",
X"0c83c08c",
X"08c80508",
X"83c08c08",
X"ffb80508",
X"34880b83",
X"c08c08ff",
X"b8050881",
X"0534800b",
X"83c08c08",
X"ffb80508",
X"82053483",
X"c08c08ff",
X"b8050808",
X"ffa1ff06",
X"a0800783",
X"c08c08ff",
X"b805080c",
X"83c08c08",
X"c8050881",
X"057081ff",
X"0683c08c",
X"08c8050c",
X"83c08c08",
X"ffb8050c",
X"810b83c0",
X"8c08c805",
X"0827fedb",
X"3883c08c",
X"08ec0570",
X"5483c08c",
X"08cc050c",
X"925283c0",
X"8c08d405",
X"085180dc",
X"843f83c0",
X"800881ff",
X"067083c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffbc",
X"050891c6",
X"3883c08c",
X"08f40551",
X"f18c3f83",
X"c0800883",
X"ffff0683",
X"c08c08f6",
X"055283c0",
X"8c08e005",
X"0cf0f33f",
X"83c08008",
X"83ffff06",
X"83c08c08",
X"fd053383",
X"c08c08ff",
X"bc050883",
X"c08c08c8",
X"050c83c0",
X"8c08c005",
X"0c83c08c",
X"08dc050c",
X"83c08c08",
X"c8050883",
X"c08c08c0",
X"05082780",
X"fe3883c0",
X"8c08cc05",
X"085483c0",
X"8c08c805",
X"08538952",
X"83c08c08",
X"d4050851",
X"80db8b3f",
X"83c08008",
X"81ff0683",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"bc050883",
X"eb3883c0",
X"8c08ee05",
X"51eff33f",
X"83c08008",
X"83ffff06",
X"5383c08c",
X"08c80508",
X"5283c08c",
X"08d40508",
X"51f0b53f",
X"83c08c08",
X"c8050881",
X"057081ff",
X"0683c08c",
X"08c8050c",
X"83c08c08",
X"ffb8050c",
X"fef23983",
X"c08c08c4",
X"05088105",
X"3383c08c",
X"08c0050c",
X"83c08c08",
X"c0050883",
X"9e3883c0",
X"8c08c005",
X"0883c08c",
X"08ffb805",
X"0c83c08c",
X"08e00508",
X"88de2e09",
X"81068b38",
X"810b83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08dc05",
X"08858e2e",
X"09810682",
X"c5388170",
X"83c08c08",
X"ffb80508",
X"0683c08c",
X"08ffb805",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"ffb80508",
X"802e829e",
X"3883c08c",
X"08c80508",
X"83c08c08",
X"c4050881",
X"053483c0",
X"8c08c005",
X"0883c08c",
X"08c40508",
X"87053483",
X"c08c08c0",
X"050883c0",
X"8c08c405",
X"088b0534",
X"83c08c08",
X"c0050883",
X"c08c08c4",
X"05088c05",
X"34830b83",
X"c08c08c4",
X"05088d05",
X"3483c08c",
X"08c00508",
X"83c08c08",
X"c405088e",
X"0523830b",
X"83c08c08",
X"c405088a",
X"053483c0",
X"8c08c405",
X"08940508",
X"83808007",
X"83c08c08",
X"c4050894",
X"050c83ca",
X"f4337083",
X"c08c08c8",
X"05080583",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"b8050883",
X"caf43483",
X"c08c08ff",
X"bc050883",
X"c08c08c4",
X"05089405",
X"3483c08c",
X"08c80508",
X"83c08c08",
X"c4050880",
X"d6053483",
X"c08c08c8",
X"050883c0",
X"8c08c405",
X"08840534",
X"8e0b83c0",
X"8c08c405",
X"08850534",
X"83c08c08",
X"c0050883",
X"c08c08c4",
X"05088605",
X"3483c08c",
X"08c40508",
X"840508ff",
X"83ff0682",
X"800783c0",
X"8c08c405",
X"0884050c",
X"a23981db",
X"0b83c08c",
X"08ffb805",
X"0c8cc339",
X"83c08c08",
X"ffbc0508",
X"83c08c08",
X"ffb8050c",
X"8cb03983",
X"c08c08f1",
X"05335283",
X"c08c08d4",
X"05085180",
X"d7903f80",
X"0b83c08c",
X"08c40508",
X"81053383",
X"c08c08ff",
X"b8050c83",
X"c08c08c8",
X"050c83c0",
X"8c08c805",
X"0883c08c",
X"08ffb805",
X"08278acb",
X"3883c08c",
X"08c80508",
X"80d82970",
X"83c08c08",
X"c4050805",
X"70880570",
X"83053383",
X"c08c08ff",
X"b8050c83",
X"c08c08cc",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08d805",
X"0c83c08c",
X"08ffb805",
X"08888938",
X"83c08c08",
X"ffbc0508",
X"8d053383",
X"c08c08d0",
X"050c83c0",
X"8c08d005",
X"0887ed38",
X"83c08c08",
X"cc050822",
X"02840571",
X"860587ff",
X"fc0683c0",
X"8c08ffb8",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08c0050c",
X"0283c08c",
X"08ffb805",
X"08310d89",
X"3d705983",
X"c08c08c0",
X"05085883",
X"c08c08ff",
X"bc050887",
X"05335783",
X"c08c08ff",
X"b8050ca2",
X"5583c08c",
X"08d00508",
X"54865381",
X"815283c0",
X"8c08d405",
X"085180c9",
X"c33f83c0",
X"800881ff",
X"0683c08c",
X"08d0050c",
X"83c08c08",
X"d0050881",
X"c03883c0",
X"8c08ffbc",
X"05089605",
X"5383c08c",
X"08c00508",
X"5283c08c",
X"08ffb805",
X"0851acf7",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"802e8185",
X"3883c08c",
X"08ffbc05",
X"08940583",
X"c08c08ff",
X"bc050896",
X"05337086",
X"2a83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08c0050c",
X"83c08c08",
X"ffb80508",
X"832e0981",
X"0680c638",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"cc050882",
X"053483ca",
X"f4337081",
X"0583c08c",
X"08ffb805",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffb805",
X"0883caf4",
X"3483c08c",
X"08ffbc05",
X"0883c08c",
X"08c00508",
X"3483c08c",
X"08e40508",
X"0d83c08c",
X"08d00508",
X"81ff0683",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"bc0508fb",
X"e33883c0",
X"8c08d805",
X"0883c08c",
X"08c40508",
X"05880570",
X"82053351",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"832e0981",
X"0680e338",
X"83c08c08",
X"ffbc0508",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"81057081",
X"ff065183",
X"c08c08ff",
X"b8050c81",
X"0b83c08c",
X"08ffb805",
X"0827dd38",
X"800b83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"05088105",
X"7081ff06",
X"5183c08c",
X"08ffb805",
X"0c970b83",
X"c08c08ff",
X"b8050827",
X"dd3883c0",
X"8c08e005",
X"0880f932",
X"70307080",
X"25515183",
X"c08c08ff",
X"b8050c83",
X"c08c08dc",
X"0508912e",
X"09810680",
X"f93883c0",
X"8c08ffb8",
X"0508802e",
X"80ec3883",
X"c08c08c8",
X"050880e2",
X"38850b83",
X"c08c08c4",
X"0508a605",
X"34a00b83",
X"c08c08c4",
X"0508a705",
X"34850b83",
X"c08c08c4",
X"0508a805",
X"3480c00b",
X"83c08c08",
X"c40508a9",
X"0534860b",
X"83c08c08",
X"c40508aa",
X"0534900b",
X"83c08c08",
X"c40508ab",
X"0534860b",
X"83c08c08",
X"c40508ac",
X"0534a00b",
X"83c08c08",
X"c40508ad",
X"053483c0",
X"8c08e005",
X"0889d832",
X"70307080",
X"25515183",
X"c08c08ff",
X"b8050c83",
X"c08c08dc",
X"050883ed",
X"ec2e0981",
X"0680f638",
X"817083c0",
X"8c08ffb8",
X"05080683",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"b8050880",
X"2e80ce38",
X"83c08c08",
X"c8050880",
X"c438840b",
X"83c08c08",
X"c40508aa",
X"053480c0",
X"0b83c08c",
X"08c40508",
X"ab053484",
X"0b83c08c",
X"08c40508",
X"ac053490",
X"0b83c08c",
X"08c40508",
X"ad053483",
X"c08c08ff",
X"bc050883",
X"c08c08c4",
X"05088c05",
X"3483c08c",
X"08e00508",
X"80f93270",
X"30708025",
X"515183c0",
X"8c08ffb8",
X"050c83c0",
X"8c08dc05",
X"08862e09",
X"810680c3",
X"38817083",
X"c08c08ff",
X"b8050806",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb80508",
X"802e9c38",
X"83c08c08",
X"c8050893",
X"3883c08c",
X"08ffbc05",
X"0883c08c",
X"08c40508",
X"8d053483",
X"c08c08e0",
X"0508b4b4",
X"32703070",
X"80255151",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"dc050890",
X"892e0981",
X"06a23883",
X"c08c08ff",
X"b8050880",
X"2e963883",
X"c08c08c8",
X"05088d38",
X"820b83c0",
X"8c08c405",
X"088d0534",
X"83c08c08",
X"c8050880",
X"d82983c0",
X"8c08c405",
X"08057084",
X"05708305",
X"3383c08c",
X"08ffb805",
X"0c83c08c",
X"08cc050c",
X"83c08c08",
X"c0050c80",
X"58805783",
X"c08c08ff",
X"b8050856",
X"80558054",
X"8a53a152",
X"83c08c08",
X"d4050851",
X"80c1f53f",
X"83c08008",
X"81ff0670",
X"30709f2a",
X"5183c08c",
X"08ffb805",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffbc05",
X"08a02e8c",
X"3883c08c",
X"08ffb805",
X"08f5dd38",
X"83c08c08",
X"c005088b",
X"053383c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"0508802e",
X"b43883c0",
X"8c08cc05",
X"08830533",
X"83c08c08",
X"ffb8050c",
X"80588057",
X"83c08c08",
X"ffb80508",
X"56805580",
X"548b53a1",
X"5283c08c",
X"08d40508",
X"5180c0f0",
X"3f83c08c",
X"08c80508",
X"81057081",
X"ff0683c0",
X"8c08c405",
X"08810533",
X"5283c08c",
X"08c8050c",
X"83c08c08",
X"ffb8050c",
X"f5a43980",
X"0b83c08c",
X"08c8050c",
X"83c08c08",
X"c8050880",
X"d82983c0",
X"8c08d405",
X"0805709a",
X"053383c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb8",
X"0508822e",
X"098106a9",
X"3883cb90",
X"56815580",
X"5483c08c",
X"08ffb805",
X"085383c0",
X"8c08ffbc",
X"05089705",
X"335283c0",
X"8c08d405",
X"0851e0ae",
X"3f83c08c",
X"08c80508",
X"81057081",
X"ff0683c0",
X"8c08c805",
X"0c83c08c",
X"08ffb805",
X"0c810b83",
X"c08c08c8",
X"050827fe",
X"fb38810b",
X"83c08c08",
X"c4050834",
X"800b83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08e805",
X"080d83c0",
X"8c08ffb8",
X"050883c0",
X"800c9b3d",
X"0d83c08c",
X"0c04f43d",
X"0d901f59",
X"800b811a",
X"33555b7a",
X"742781ad",
X"387a80d8",
X"29198a11",
X"33555573",
X"832e0981",
X"06818838",
X"94153357",
X"80527651",
X"dde03f80",
X"53805276",
X"51de803f",
X"b3e43f83",
X"c080085c",
X"80587781",
X"c4291c87",
X"11335555",
X"73802e80",
X"c0387408",
X"81ecb82e",
X"098106b5",
X"3880755b",
X"567580d8",
X"291a9a11",
X"33555573",
X"832e0981",
X"069238a4",
X"15703355",
X"55767427",
X"8738ff14",
X"54737534",
X"81167081",
X"ff065754",
X"817627d1",
X"38811870",
X"81ff0659",
X"548f7827",
X"ffa43883",
X"caf433ff",
X"05547383",
X"caf43481",
X"1b7081ff",
X"06811b33",
X"5f5c547c",
X"7b26fed5",
X"38800b83",
X"c0800c8e",
X"3d0d0483",
X"c08c0802",
X"83c08c0c",
X"e63d0d83",
X"c08c0888",
X"05080284",
X"05719005",
X"70337083",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08cc",
X"050c83c0",
X"8c08dc05",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"ffa40508",
X"802e9f8c",
X"38800b83",
X"c08c08cc",
X"05088105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08d4050c",
X"83c08c08",
X"d4050883",
X"c08c08ff",
X"a4050825",
X"9ed43883",
X"c08c08d4",
X"050880d8",
X"2983c08c",
X"08cc0508",
X"05840570",
X"86053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"a4050880",
X"2e9de038",
X"b18a3f83",
X"c08c08ff",
X"bc050880",
X"d4050883",
X"c0800826",
X"9dc93802",
X"83c08c08",
X"ffbc0508",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08d8",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08fc05",
X"2383c08c",
X"08ffa405",
X"08860583",
X"fc0683c0",
X"8c08ffa4",
X"050c0283",
X"c08c08ff",
X"a4050831",
X"0d853d70",
X"5583c08c",
X"08fc0554",
X"83c08c08",
X"ffbc0508",
X"5383c08c",
X"08e00508",
X"5283c08c",
X"08c0050c",
X"b8e23f83",
X"c0800881",
X"ff0683c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"05089c92",
X"3883c08c",
X"08ffbc05",
X"08870533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e80d5",
X"3883c08c",
X"08ffbc05",
X"08860533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"822e0981",
X"06b33883",
X"c08c08fc",
X"052283c0",
X"8c08ffa4",
X"050c870b",
X"83c08c08",
X"ffa40508",
X"27973883",
X"c08c08c0",
X"05088205",
X"5283c08c",
X"08c00508",
X"3351d7b4",
X"3f83c08c",
X"08ffbc05",
X"08860533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"832e0981",
X"069afb38",
X"83c08c08",
X"ffbc0508",
X"920583c0",
X"8c08ffbc",
X"05088905",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08c4050c",
X"83c08c08",
X"ffa40508",
X"832eb638",
X"83c08c08",
X"c4050882",
X"053383c0",
X"8c08fc05",
X"2283c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa805",
X"0883c08c",
X"08ffac05",
X"08269a96",
X"38800b83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa40508",
X"832e0981",
X"0688c138",
X"83c08c08",
X"c0050833",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffb00508",
X"2e098106",
X"87fa3883",
X"c08c08c0",
X"05088105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08942e09",
X"810687d8",
X"3883c08c",
X"08c00508",
X"82053370",
X"810683c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffb0",
X"05082e8a",
X"38880b83",
X"c08c08e4",
X"050c83c0",
X"8c08ffa8",
X"0508812a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9138",
X"83c08c08",
X"e4050884",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"ffa80508",
X"822a7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"913883c0",
X"8c08e405",
X"08820783",
X"c08c08e4",
X"050c83c0",
X"8c08ffa8",
X"0508832a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9138",
X"83c08c08",
X"e4050881",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"c0050883",
X"05337098",
X"2b83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"08802591",
X"3883c08c",
X"08e40508",
X"900783c0",
X"8c08e405",
X"0c83c08c",
X"08ffa805",
X"0881ff06",
X"70852a70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050880",
X"2e913883",
X"c08c08e4",
X"0508a007",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"a8050884",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e92",
X"3883c08c",
X"08e40508",
X"80c00783",
X"c08c08e4",
X"050c83c0",
X"8c08ffa8",
X"0508862a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9238",
X"83c08c08",
X"e4050881",
X"800783c0",
X"8c08e405",
X"0c83c08c",
X"08ffa805",
X"08810683",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e923883",
X"c08c08e4",
X"05088280",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"ffa80508",
X"812a7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"923883c0",
X"8c08e405",
X"08848007",
X"83c08c08",
X"e4050c83",
X"c08c08c0",
X"05088405",
X"3370982b",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa40508",
X"80259238",
X"83c08c08",
X"e4050888",
X"800783c0",
X"8c08e405",
X"0c83c08c",
X"08c00508",
X"85053370",
X"982b83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"05088025",
X"923883c0",
X"8c08e405",
X"08908007",
X"83c08c08",
X"e4050c83",
X"c08c08c0",
X"05088205",
X"337081ff",
X"0670852a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa40508",
X"802e9238",
X"83c08c08",
X"e40508a0",
X"800783c0",
X"8c08e405",
X"0c83c08c",
X"08ffa805",
X"08842a70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e933883",
X"c08c08e4",
X"050880c0",
X"800783c0",
X"8c08e405",
X"0c83c08c",
X"08ffa805",
X"08862a70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e933883",
X"c08c08e4",
X"05088180",
X"800783c0",
X"8c08e405",
X"0c83c08c",
X"08ffac05",
X"08982b83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"25933883",
X"c08c08e4",
X"05088280",
X"800783c0",
X"8c08e405",
X"0c83c08c",
X"08c00508",
X"87053370",
X"982b83c0",
X"8c08c005",
X"08890533",
X"70982b70",
X"982c7398",
X"2c818005",
X"54515383",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a8050883",
X"c08c08f8",
X"052380ff",
X"0b83c08c",
X"08ffa405",
X"083183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08fa05",
X"2384d939",
X"800b83c0",
X"8c08e405",
X"0c81800b",
X"83c08c08",
X"f8052381",
X"800b83c0",
X"8c08fa05",
X"2384b939",
X"83c08c08",
X"ffb00508",
X"1083c08c",
X"0805f805",
X"83c08c08",
X"ffb00508",
X"842983c0",
X"8c08ffb0",
X"05081005",
X"83c08c08",
X"c4050805",
X"70840570",
X"3383c08c",
X"08c00508",
X"05703383",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b4050883",
X"c08c08ff",
X"b8050823",
X"83c08c08",
X"ffa80508",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050890",
X"2e098106",
X"be3883c0",
X"8c08ffa8",
X"05083383",
X"c08c08c0",
X"05080581",
X"05703370",
X"82802983",
X"c08c08ff",
X"b4050805",
X"515183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffb8",
X"05082383",
X"c08c08ff",
X"ac050886",
X"052283c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa8",
X"0508a238",
X"83c08c08",
X"ffac0508",
X"88052283",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050881",
X"ff2e80e5",
X"3883c08c",
X"08ffb805",
X"08227083",
X"c08c08ff",
X"a8050831",
X"70828029",
X"713183c0",
X"8c08ffac",
X"05088805",
X"227083c0",
X"8c08ffa8",
X"05083170",
X"73355383",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"ac050c51",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffb80508",
X"2383c08c",
X"08ffb005",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a4050c81",
X"0b83c08c",
X"08ffb005",
X"0827fce0",
X"38800b83",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"b0050810",
X"83c08c08",
X"c4050805",
X"70900570",
X"3383c08c",
X"08c00508",
X"05703372",
X"81053370",
X"72065153",
X"5183c08c",
X"08ffa805",
X"0c5183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"9b38900b",
X"83c08c08",
X"ffb00508",
X"2b83c08c",
X"08e40508",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"ffb00508",
X"81057081",
X"ff0683c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa4",
X"050c970b",
X"83c08c08",
X"ffb00508",
X"27fef438",
X"83c08c08",
X"f8052283",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a40508bf",
X"26913883",
X"c08c08e4",
X"05088207",
X"83c08c08",
X"e4050c81",
X"c00b83c0",
X"8c08ffa4",
X"05082791",
X"3883c08c",
X"08e40508",
X"810783c0",
X"8c08e405",
X"0c83c08c",
X"08fa0522",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"bf269138",
X"83c08c08",
X"e4050888",
X"0783c08c",
X"08e4050c",
X"81c00b83",
X"c08c08ff",
X"a4050827",
X"913883c0",
X"8c08e405",
X"08840783",
X"c08c08e4",
X"050c83c0",
X"8c08ffbc",
X"05089005",
X"3383c08c",
X"08e40508",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"c4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"bc05088c",
X"05082e85",
X"e03883c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffbc",
X"05088c05",
X"0c83c08c",
X"08ffbc05",
X"08890533",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa80508",
X"802e859a",
X"3883c08c",
X"08e40583",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"a405088f",
X"0683c08c",
X"08e4050c",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"d0050c83",
X"c08c08ff",
X"a8050882",
X"2e098106",
X"81c23880",
X"0b83c08c",
X"08ffa405",
X"08862a70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"a805082e",
X"8c3881c0",
X"0b83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffb005",
X"08872a70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e943883",
X"c08c08ff",
X"a8050881",
X"903283c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffb0",
X"0508842a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9438",
X"83c08c08",
X"ffa80508",
X"80d03283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"b0050883",
X"c08c08ff",
X"a8050832",
X"83c08c08",
X"ffb0050c",
X"800b83c0",
X"8c08f005",
X"0c800b83",
X"c08c08f4",
X"0523800b",
X"81eeb433",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffb80508",
X"2e82d338",
X"83c08c08",
X"f00581ee",
X"b40b83c0",
X"8c08ffac",
X"050c83c0",
X"8c08c805",
X"0c83c08c",
X"08ffac05",
X"083383c0",
X"8c08ffac",
X"05088105",
X"3381722b",
X"81722b07",
X"7083c08c",
X"08ffb005",
X"08065283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"a805082e",
X"09810681",
X"be3883c0",
X"8c08ffb8",
X"05088526",
X"80f63883",
X"c08c08ff",
X"ac050882",
X"05337081",
X"ff0683c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"80ca3883",
X"c08c08ff",
X"b8050883",
X"c08c08ff",
X"b8050881",
X"057081ff",
X"0683c08c",
X"08c80508",
X"73055383",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b4050883",
X"c08c08ff",
X"a4050834",
X"83c08c08",
X"ffac0508",
X"83053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e9d3881",
X"0b83c08c",
X"08ffa405",
X"082b83c0",
X"8c08d005",
X"08080783",
X"c08c08d0",
X"05080c83",
X"c08c08ff",
X"ac050884",
X"05703383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a40508fd",
X"c83883c0",
X"8c08f005",
X"528051c1",
X"fb3f83c0",
X"8c08e405",
X"085283c0",
X"8c08c405",
X"0851c3b6",
X"3f83c08c",
X"08fb0533",
X"7081800a",
X"29810a05",
X"70982c55",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"f9053370",
X"81800a29",
X"810a0570",
X"982c5583",
X"c08c08ff",
X"a4050c83",
X"c08c08c4",
X"05085383",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a8050cc3",
X"8e3f83c0",
X"8c08ffbc",
X"05088805",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e84",
X"e13883c0",
X"8c08ffbc",
X"05089005",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08812684",
X"c1388070",
X"81eef40b",
X"81eef40b",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"b405082e",
X"81ae3883",
X"c08c08ff",
X"ac050884",
X"2983c08c",
X"08ffa805",
X"08057033",
X"83c08c08",
X"c0050805",
X"70337281",
X"05337072",
X"06515351",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802eaa38",
X"810b83c0",
X"8c08ffac",
X"05082b83",
X"c08c08ff",
X"b4050807",
X"7083ffff",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffac05",
X"08810570",
X"81ff0681",
X"eef47184",
X"29710570",
X"81053351",
X"5383c08c",
X"08ffa805",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08fed438",
X"83c08c08",
X"ffbc0508",
X"8a052283",
X"c08c08c0",
X"050c83c0",
X"8c08ffb4",
X"050883c0",
X"8c08c005",
X"082e82ae",
X"38800b83",
X"c08c08e8",
X"050c800b",
X"83c08c08",
X"ec052380",
X"7083c08c",
X"08e80583",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"b0050c81",
X"af3983c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffac",
X"05082c70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e80e738",
X"83c08c08",
X"ffb00508",
X"83c08c08",
X"ffb00508",
X"81057081",
X"ff0683c0",
X"8c08ffb8",
X"05087305",
X"83c08c08",
X"ffbc0508",
X"90053383",
X"c08c08ff",
X"ac050884",
X"29055353",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa80508",
X"81eef605",
X"3383c08c",
X"08ffa405",
X"083483c0",
X"8c08ffac",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa4050c",
X"8f0b83c0",
X"8c08ffac",
X"05082783",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b0050885",
X"268c3883",
X"c08c08ff",
X"a40508fe",
X"a93883c0",
X"8c08e805",
X"528051ff",
X"bcaa3f83",
X"c08c08ff",
X"b4050883",
X"c08c08ff",
X"bc05088a",
X"052383c0",
X"8c08ffbc",
X"050880d2",
X"053383c0",
X"8c08ffbc",
X"050880d4",
X"05080583",
X"c08c08ff",
X"bc050880",
X"d4050c83",
X"c08c08d8",
X"05080d83",
X"c08c08d4",
X"05088180",
X"0a298180",
X"0a057098",
X"2c83c08c",
X"08cc0508",
X"81053383",
X"c08c08ff",
X"a8050c51",
X"83c08c08",
X"d4050c83",
X"c08c08ff",
X"a8050883",
X"c08c08d4",
X"050824e1",
X"ae38800b",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"dc05080d",
X"83c08c08",
X"ffa80508",
X"83c0800c",
X"9c3d0d83",
X"c08c0c04",
X"f33d0d02",
X"bf053302",
X"840580c3",
X"053383cb",
X"90335a5b",
X"5979802e",
X"8d387878",
X"06577680",
X"2e8e3881",
X"8a397878",
X"06577680",
X"2e818038",
X"83cb9033",
X"707a0758",
X"58798838",
X"78097079",
X"06515776",
X"83cb9034",
X"92983f83",
X"c080085e",
X"805c8f5d",
X"7d1c8711",
X"33585876",
X"802e80c2",
X"38770881",
X"ecb82e09",
X"8106b738",
X"805b815a",
X"7d1c701c",
X"9a113359",
X"59597682",
X"2e098106",
X"953883cb",
X"90568155",
X"80547653",
X"97183352",
X"7851ffbd",
X"813fff1a",
X"80d81c5c",
X"5a798025",
X"cf38ff1d",
X"81c41d5d",
X"5d7c8025",
X"ffa6388f",
X"3d0d04e9",
X"3d0d696c",
X"02880580",
X"ea05225c",
X"5a5b8070",
X"71415e58",
X"ff78797a",
X"7b7c7d46",
X"4c4a4540",
X"5d436299",
X"3d346202",
X"840580dd",
X"05347779",
X"2280ffff",
X"06544572",
X"79237978",
X"2e888738",
X"7a708105",
X"5c337084",
X"2a718c06",
X"70822a5a",
X"56568306",
X"ff1b7083",
X"ffff065c",
X"54568054",
X"75742e91",
X"387a7081",
X"055c33ff",
X"1b7083ff",
X"ff065c54",
X"54817627",
X"9b387381",
X"ff067b70",
X"81055d33",
X"55748280",
X"2905ff1b",
X"7083ffff",
X"065c5454",
X"827627aa",
X"387383ff",
X"ff067b70",
X"81055d33",
X"70902b72",
X"077d7081",
X"055f3370",
X"982b7207",
X"fe1f7083",
X"ffff0640",
X"52525252",
X"54547e80",
X"2e80c438",
X"7686f738",
X"748a2e09",
X"81069438",
X"811f7081",
X"ff06811e",
X"7081ff06",
X"5f524053",
X"86dc3974",
X"8c2e0981",
X"0686d338",
X"ff1f7081",
X"ff06ff1e",
X"7081ff06",
X"5f524053",
X"7b632586",
X"bd38ff43",
X"86b83976",
X"812e83bb",
X"38768124",
X"89387680",
X"2e8d3886",
X"a5397682",
X"2e84a638",
X"869c39f8",
X"15537284",
X"26849538",
X"72842981",
X"efb40553",
X"72080464",
X"802e80cd",
X"38782283",
X"80800653",
X"72838080",
X"2e098106",
X"bc388056",
X"756427a4",
X"38751e70",
X"83ffff06",
X"77101b90",
X"1172832a",
X"58515751",
X"53737534",
X"72870681",
X"712b5153",
X"72811634",
X"81167081",
X"ff065753",
X"977627cc",
X"387f8407",
X"40800b99",
X"3d435661",
X"16703370",
X"982b7098",
X"2c515151",
X"53807324",
X"80fb3860",
X"73291e70",
X"83ffff06",
X"7a228380",
X"80065258",
X"53728380",
X"802e0981",
X"0680de38",
X"60883270",
X"30707207",
X"80256390",
X"32703070",
X"72078025",
X"73075354",
X"58515553",
X"73802ebd",
X"38768706",
X"5372b638",
X"75842976",
X"10057911",
X"84117983",
X"2a575751",
X"53737534",
X"60811634",
X"65861423",
X"66881423",
X"7587387f",
X"8107408d",
X"3975812e",
X"09810685",
X"387f8207",
X"40811670",
X"81ff0657",
X"53817627",
X"fee53863",
X"61291e70",
X"83ffff06",
X"5f538070",
X"4642ff02",
X"840580dd",
X"0534ff0b",
X"993d3483",
X"f539811c",
X"7081ff06",
X"5d538042",
X"73812e09",
X"81068e38",
X"7781800a",
X"2981800a",
X"055880d3",
X"3973802e",
X"89387382",
X"2e098106",
X"8d387c81",
X"800a2981",
X"800a055d",
X"a439815f",
X"83b839ff",
X"1c7081ff",
X"065d537b",
X"63258338",
X"ff437c80",
X"2e92387c",
X"81800a29",
X"81ff0a05",
X"5d7c982c",
X"5d839339",
X"77802e92",
X"38778180",
X"0a2981ff",
X"0a055877",
X"982c5882",
X"fd397753",
X"839e3974",
X"892680f4",
X"38748429",
X"81efc805",
X"53720804",
X"73872e82",
X"e1387385",
X"2e82db38",
X"73882e82",
X"d538738c",
X"2e82cf38",
X"73892e09",
X"81068638",
X"814582c2",
X"3973812e",
X"09810682",
X"b9386280",
X"2582b338",
X"7b982b70",
X"982c5143",
X"82a83973",
X"83ffff06",
X"46829f39",
X"7383ffff",
X"06478296",
X"397381ff",
X"0641828e",
X"3973811a",
X"34828739",
X"7381ff06",
X"4481ff39",
X"7e5382a0",
X"3974812e",
X"81e33874",
X"81248938",
X"74802e8d",
X"3881e739",
X"74822e81",
X"d83881de",
X"3974567b",
X"83388156",
X"74537386",
X"2e098106",
X"97387581",
X"06537280",
X"2e8e3878",
X"2282ffff",
X"06fe8080",
X"0753b639",
X"7b833881",
X"5373822e",
X"09810697",
X"38728106",
X"5372802e",
X"8e387822",
X"81ffff06",
X"81808007",
X"5393397b",
X"9638fc14",
X"53728126",
X"8e387822",
X"ff808007",
X"53727923",
X"80e53980",
X"5573812e",
X"09810683",
X"38735577",
X"5377802e",
X"89387481",
X"06537280",
X"ca3872d0",
X"15545572",
X"81268338",
X"81557780",
X"2eb93874",
X"81065372",
X"802eb038",
X"78228380",
X"80065372",
X"8380802e",
X"0981069f",
X"3873b02e",
X"09810687",
X"3861993d",
X"34913973",
X"b12e0981",
X"06893861",
X"02840580",
X"dd053461",
X"8105538c",
X"39617431",
X"81055384",
X"39611453",
X"7283ffff",
X"064279f7",
X"fb387d83",
X"2a537282",
X"1a347822",
X"83808006",
X"53728380",
X"802e0981",
X"06883881",
X"537f872e",
X"83388053",
X"7283c080",
X"0c993d0d",
X"04fd3d0d",
X"75831133",
X"82123371",
X"982b7190",
X"2b078114",
X"3370882b",
X"72077533",
X"710783c0",
X"800c5253",
X"54565452",
X"853d0d04",
X"f63d0d02",
X"b7053302",
X"8405bb05",
X"33028805",
X"bf05335b",
X"5b5b8058",
X"80577888",
X"2b7a0756",
X"80557a54",
X"8153a352",
X"7c5192cc",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8c3d0d04",
X"f63d0d02",
X"b7053302",
X"8405bb05",
X"33028805",
X"bf05335b",
X"5b5b8058",
X"80577888",
X"2b7a0756",
X"80557a54",
X"8353a352",
X"7c519290",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8c3d0d04",
X"f73d0d02",
X"b3053302",
X"8405b605",
X"22605a58",
X"56805580",
X"54805381",
X"a3527b51",
X"91e23f83",
X"c0800881",
X"ff0683c0",
X"800c8b3d",
X"0d04ee3d",
X"0d649011",
X"5c5c807b",
X"34800b84",
X"1c0c800b",
X"881c3481",
X"0b891c34",
X"880b8a1c",
X"34800b8b",
X"1c34881b",
X"08c10681",
X"07881c0c",
X"8f3d7054",
X"5d88527b",
X"519c923f",
X"83c08008",
X"81ff0670",
X"5b597881",
X"a938903d",
X"335e81db",
X"5a7d892e",
X"09810681",
X"99387c53",
X"92527b51",
X"9beb3f83",
X"c0800881",
X"ff06705b",
X"59788182",
X"387c5888",
X"577856a9",
X"55785486",
X"5381a052",
X"7b5190d0",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"80e03802",
X"ba05337b",
X"347c5478",
X"537d527b",
X"519bd33f",
X"83c08008",
X"81ff0670",
X"5b597880",
X"c13802bd",
X"0533527b",
X"519beb3f",
X"83c08008",
X"81ff0670",
X"5b5978aa",
X"38817b33",
X"5a5a7979",
X"26993880",
X"54795388",
X"527b51fd",
X"bb3f811a",
X"7081ff06",
X"7c33525b",
X"59e43981",
X"0b881c34",
X"805a7983",
X"c0800c94",
X"3d0d0480",
X"0b83c080",
X"0c04f93d",
X"0d790284",
X"05ab0533",
X"8e3d7054",
X"585858ff",
X"afec3f8a",
X"3d8a0551",
X"ffafe33f",
X"7551fc8d",
X"3f83c080",
X"08848681",
X"2ebe3883",
X"c0800884",
X"86812699",
X"3883c080",
X"08848280",
X"2e80e638",
X"83c08008",
X"8482812e",
X"9f3881b4",
X"3983c080",
X"0880c082",
X"832e80f4",
X"3883c080",
X"0880c086",
X"832e80e8",
X"38819939",
X"83c09c33",
X"55805674",
X"762e0981",
X"06818b38",
X"74547653",
X"91527751",
X"fbd63f74",
X"54765390",
X"527751fb",
X"cb3f7454",
X"76538452",
X"7751fbfc",
X"3f810b83",
X"c09c3481",
X"b15680de",
X"39805476",
X"53915277",
X"51fba93f",
X"80547653",
X"90527751",
X"fb9e3f80",
X"0b83c09c",
X"34765287",
X"18335197",
X"963fb539",
X"80547653",
X"94527751",
X"fb823f80",
X"54765390",
X"527751fa",
X"f73f7551",
X"ffae973f",
X"83c08008",
X"892a8106",
X"53765287",
X"18335190",
X"cd3f800b",
X"83c09c34",
X"80567583",
X"c0800c89",
X"3d0d04f2",
X"3d0d6090",
X"115a5880",
X"0b881a33",
X"71595656",
X"74762e82",
X"a53882ac",
X"3f841908",
X"83c08008",
X"26829538",
X"78335a81",
X"0b8e3d23",
X"903df811",
X"55f40553",
X"99185277",
X"518ae53f",
X"83c08008",
X"81ff0670",
X"57557477",
X"2e098106",
X"81d93886",
X"39745681",
X"d2398156",
X"82578e3d",
X"33770655",
X"74802ebb",
X"38800b8d",
X"3d34903d",
X"f0055484",
X"53755277",
X"51facd3f",
X"83c08008",
X"81ff0655",
X"749d387b",
X"53755277",
X"51fce73f",
X"83c08008",
X"81ff0655",
X"7481b12e",
X"818b3874",
X"ffb33876",
X"1081fc06",
X"81177081",
X"ff065856",
X"57877627",
X"ffa83881",
X"56757a26",
X"80eb3880",
X"0b8d3d34",
X"8c3d7055",
X"57845375",
X"527751f9",
X"f73f83c0",
X"800881ff",
X"06557480",
X"c1387651",
X"ffac933f",
X"83c08008",
X"82870655",
X"7482812e",
X"098106aa",
X"3802ae05",
X"33810755",
X"74028405",
X"ae05347b",
X"53755277",
X"51fbeb3f",
X"83c08008",
X"81ff0655",
X"7481b12e",
X"903874fe",
X"b8388116",
X"7081ff06",
X"5755ff91",
X"39805675",
X"81ff0656",
X"973f83c0",
X"80088fd0",
X"05841a0c",
X"75577683",
X"c0800c90",
X"3d0d0404",
X"9080a008",
X"83c0800c",
X"04ff3d0d",
X"7387e829",
X"51fefdc2",
X"3f833d0d",
X"040483cb",
X"940b83c0",
X"800c04fd",
X"3d0d7577",
X"5454800b",
X"83caf434",
X"728a3890",
X"90800b84",
X"150c9039",
X"72812e09",
X"81068838",
X"9098800b",
X"84150c84",
X"140883cb",
X"8c0c800b",
X"88150c80",
X"0b8c150c",
X"83cb8c08",
X"53820b87",
X"80143481",
X"51ff9e3f",
X"83cb8c08",
X"53800b88",
X"143483cb",
X"8c085381",
X"0b878014",
X"3483cb8c",
X"0853800b",
X"8c143483",
X"cb8c0853",
X"800ba414",
X"34917434",
X"800b83c0",
X"a034800b",
X"83c0a434",
X"800b83c0",
X"a8348054",
X"7381c429",
X"83cb9805",
X"53800b83",
X"14348114",
X"7081ff06",
X"55538f74",
X"27e63885",
X"3d0d04fe",
X"3d0d7476",
X"82113370",
X"bf068171",
X"2bff0556",
X"51515253",
X"90712783",
X"38ff5276",
X"51717123",
X"83cb8c08",
X"51871333",
X"90123480",
X"0b83c0a4",
X"34800b83",
X"c0a83488",
X"13338a14",
X"33525271",
X"802eaa38",
X"7081ff06",
X"51845270",
X"83387052",
X"7183c0a4",
X"348a1333",
X"70307080",
X"25842b70",
X"88075151",
X"52537083",
X"c0a83490",
X"397081ff",
X"06517083",
X"38985271",
X"83c0a834",
X"800b83c0",
X"800c843d",
X"0d04f13d",
X"0d616568",
X"028c0580",
X"cb053302",
X"900580ce",
X"05220294",
X"0580d605",
X"22424041",
X"5a4040fd",
X"8b3f83c0",
X"8008a788",
X"055b8070",
X"715b5b52",
X"83943983",
X"cb8c0851",
X"7d941234",
X"83c0a433",
X"81075580",
X"7054567f",
X"862680ea",
X"387f8429",
X"81effc05",
X"83cb8c08",
X"53517008",
X"04800b84",
X"1334a139",
X"77337030",
X"70802583",
X"71315151",
X"52537084",
X"13348d39",
X"810b8413",
X"34b83983",
X"0b841334",
X"81705456",
X"ad39810b",
X"841334a2",
X"39773370",
X"30708025",
X"83713151",
X"51525370",
X"84133480",
X"78335252",
X"70833881",
X"52717834",
X"81537488",
X"075583c0",
X"a83383cb",
X"8c085257",
X"810b81d0",
X"123483cb",
X"8c085181",
X"0b819012",
X"347e802e",
X"ae387280",
X"2ea9387e",
X"ff1e5254",
X"7083ffff",
X"06537283",
X"ffff2e97",
X"38737081",
X"05553383",
X"cb8c0853",
X"517081c0",
X"1334ff13",
X"51de3983",
X"cb8c08a8",
X"11335351",
X"76881234",
X"83cb8c08",
X"51747134",
X"81ff5291",
X"3983cb8c",
X"08a01133",
X"70810651",
X"5253708f",
X"38fafd3f",
X"7a83c080",
X"0826e638",
X"81883981",
X"0ba01434",
X"83cb8c08",
X"a8113380",
X"ff067078",
X"07525351",
X"70802e80",
X"ed387186",
X"2a708106",
X"51517080",
X"2e913880",
X"78335253",
X"70833881",
X"53727834",
X"80e03971",
X"842a7081",
X"06515170",
X"802e9b38",
X"81197083",
X"ffff067d",
X"30709f2a",
X"51525a51",
X"787c2e09",
X"8106af38",
X"a4397183",
X"2a708106",
X"51517080",
X"2e933881",
X"1a7081ff",
X"065b5179",
X"832e0981",
X"0690388a",
X"3971a306",
X"5170802e",
X"85387151",
X"9239f9e4",
X"3f7a83c0",
X"800826fc",
X"e2387181",
X"bf065170",
X"83c0800c",
X"913d0d04",
X"f63d0d02",
X"b3053302",
X"8405b705",
X"33028805",
X"ba052259",
X"5959800b",
X"8c3d348c",
X"3dfc0556",
X"80558054",
X"76537752",
X"7851fbf2",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8c3d0d04",
X"f33d0d7f",
X"6264028c",
X"0580c205",
X"22722281",
X"1533425f",
X"415e5959",
X"8078237d",
X"53783352",
X"8151ffa0",
X"3f83c080",
X"0881ff06",
X"5675802e",
X"86387554",
X"81ad3983",
X"cb8c08a8",
X"1133821b",
X"3370862a",
X"70810673",
X"982b5351",
X"575c5657",
X"79802583",
X"38815673",
X"762e8738",
X"81f05481",
X"8239818c",
X"17337081",
X"ff067922",
X"7d713190",
X"2b70902c",
X"7009709f",
X"2c720670",
X"52525351",
X"53575754",
X"75742483",
X"38755574",
X"84808029",
X"fc808005",
X"70902c51",
X"5574ff2e",
X"943883cb",
X"8c088180",
X"11335154",
X"737c7081",
X"055e34db",
X"39772276",
X"05547378",
X"23790970",
X"9f2a7081",
X"06821c33",
X"81bf0671",
X"862b0751",
X"51515473",
X"821a347c",
X"76268a38",
X"7722547a",
X"7426febb",
X"38805473",
X"83c0800c",
X"8f3d0d04",
X"f93d0d7a",
X"57800b89",
X"3d23893d",
X"fc055376",
X"527951f8",
X"da3f83c0",
X"800881ff",
X"06705755",
X"7496387c",
X"547b5388",
X"3d225276",
X"51fde53f",
X"83c08008",
X"81ff0656",
X"7583c080",
X"0c893d0d",
X"04f03d0d",
X"62660288",
X"0580ce05",
X"22415d5e",
X"80028405",
X"80d20522",
X"7f810533",
X"ff115a5d",
X"5a5d81da",
X"5876bf26",
X"80e93878",
X"802e80e1",
X"387a5878",
X"7b278338",
X"7858821e",
X"3370872a",
X"585a7692",
X"3d34923d",
X"fc055677",
X"557b547e",
X"537d3352",
X"8251f8de",
X"3f83c080",
X"0881ff06",
X"5d800b92",
X"3d33585a",
X"76802e83",
X"38815a82",
X"1e3380ff",
X"067a872b",
X"07577682",
X"1f347c91",
X"38787831",
X"7083ffff",
X"06791e5e",
X"5a57ff9b",
X"397c5877",
X"83c0800c",
X"923d0d04",
X"f83d0d7b",
X"028405b2",
X"05225858",
X"800b8a3d",
X"238a3dfc",
X"05537752",
X"7a51f6f7",
X"3f83c080",
X"0881ff06",
X"70575574",
X"96387d54",
X"7653893d",
X"22527751",
X"feaf3f83",
X"c0800881",
X"ff065675",
X"83c0800c",
X"8a3d0d04",
X"ec3d0d66",
X"6e028805",
X"80df0533",
X"028c0580",
X"e3053302",
X"900580e7",
X"05330294",
X"0580eb05",
X"33029805",
X"80ee0522",
X"4143415f",
X"5c405702",
X"80f20522",
X"963d2396",
X"3df00553",
X"84177053",
X"775259f6",
X"863f83c0",
X"800881ff",
X"06587781",
X"e538777a",
X"81800658",
X"40807725",
X"83388140",
X"79943d34",
X"7b028405",
X"80c90534",
X"7c028405",
X"80ca0534",
X"7d028405",
X"80cb0534",
X"7a953d34",
X"7a882a57",
X"76028405",
X"80cd0534",
X"953d2257",
X"76028405",
X"80ce0534",
X"76882a57",
X"76028405",
X"80cf0534",
X"77923d34",
X"963dec11",
X"57578855",
X"f4175492",
X"3d225377",
X"527751f6",
X"953f83c0",
X"800881ff",
X"06587780",
X"ed387e80",
X"2e80cb38",
X"923d2279",
X"0858587f",
X"802e9c38",
X"76818080",
X"07790c7e",
X"54963dfc",
X"05537783",
X"ffff0652",
X"7851f9fc",
X"3f993976",
X"82808007",
X"790c7e54",
X"953d2253",
X"7783ffff",
X"06527851",
X"fc8f3f83",
X"c0800881",
X"ff065877",
X"9d38923d",
X"22538052",
X"7f307080",
X"25847131",
X"535157f9",
X"873f83c0",
X"800881ff",
X"06587783",
X"c0800c96",
X"3d0d04f6",
X"3d0d7c02",
X"8405b705",
X"335b5b80",
X"58805780",
X"56805579",
X"54855380",
X"527a51fd",
X"a33f83c0",
X"800881ff",
X"06597885",
X"3879871c",
X"347883c0",
X"800c8c3d",
X"0d04f93d",
X"0d02a705",
X"33028405",
X"ab053302",
X"8805af05",
X"33585957",
X"800b83cb",
X"9b335454",
X"72742e9f",
X"38811470",
X"81ff0655",
X"53738f26",
X"81b63873",
X"81c42983",
X"cb980583",
X"11335153",
X"72e33873",
X"81c42983",
X"cb940555",
X"800b8716",
X"34768816",
X"34758a16",
X"34778916",
X"3480750c",
X"83cb8c08",
X"8c160c80",
X"0b841634",
X"880b8516",
X"34800b86",
X"16348415",
X"08ffa1ff",
X"06a08007",
X"84160c81",
X"147081ff",
X"06535374",
X"51febc3f",
X"83c08008",
X"81ff0670",
X"55537280",
X"cd388a39",
X"7308750c",
X"725480c2",
X"397281f7",
X"9c555681",
X"f79c0880",
X"2eb23875",
X"84291470",
X"08765370",
X"08515454",
X"722d83c0",
X"800881ff",
X"06537280",
X"2ece3881",
X"167081ff",
X"0681f79c",
X"71842911",
X"53565753",
X"7208d038",
X"80547383",
X"c0800c89",
X"3d0d04f9",
X"3d0d7957",
X"800b8418",
X"0883cb8c",
X"0c58f088",
X"3f881708",
X"83c08008",
X"2783ed38",
X"effa3f83",
X"c0800881",
X"0588180c",
X"83cb8c08",
X"b8113370",
X"81ff0651",
X"51547381",
X"2ea43873",
X"81248838",
X"73782e8a",
X"38b83973",
X"822e9538",
X"b1397633",
X"81f00654",
X"73902ea6",
X"38917734",
X"a1397358",
X"763381f0",
X"06547390",
X"2e098106",
X"9138efa8",
X"3f83c080",
X"0881c805",
X"8c180ca0",
X"77348056",
X"7581c429",
X"83cb9b11",
X"33555573",
X"802eaa38",
X"83cb9415",
X"70085654",
X"74802e9d",
X"38881508",
X"802e9638",
X"8c140883",
X"cb8c082e",
X"09810689",
X"38735188",
X"15085473",
X"2d811670",
X"81ff0657",
X"548f7627",
X"ffba3876",
X"335473b0",
X"2e819938",
X"73b0248f",
X"3873912e",
X"ab3873a0",
X"2e80f538",
X"82a63973",
X"80d02e81",
X"e4387380",
X"d0248b38",
X"7380c02e",
X"81993882",
X"8f397381",
X"802e81fb",
X"38828539",
X"80567581",
X"c42983cb",
X"98118311",
X"33565955",
X"73802ea8",
X"3883cb94",
X"15700856",
X"5474802e",
X"9b388c14",
X"0883cb8c",
X"082e0981",
X"068e3873",
X"51841508",
X"54732d80",
X"0b831934",
X"81167081",
X"ff065754",
X"8f7627ff",
X"b9389277",
X"3481b539",
X"edc23f8c",
X"170883c0",
X"80082781",
X"a738b077",
X"3481a139",
X"83cb8c08",
X"54800b8c",
X"153483cb",
X"8c085484",
X"0b881534",
X"80c07734",
X"ed963f83",
X"c08008b2",
X"058c180c",
X"80fa39ed",
X"873f8c17",
X"0883c080",
X"082780ec",
X"3883cb8c",
X"0854810b",
X"8c153483",
X"cb8c0854",
X"800b8815",
X"3483cb8c",
X"0854880b",
X"a01534ec",
X"db3f83c0",
X"80089405",
X"8c180c80",
X"d07734bc",
X"3983cb8c",
X"08a01133",
X"70832a70",
X"81065151",
X"55557380",
X"2ea63888",
X"0ba01634",
X"ecae3f8c",
X"170883c0",
X"80082794",
X"38ff8077",
X"348e3977",
X"53805280",
X"51fa8b3f",
X"ff907734",
X"83cb8c08",
X"a0113370",
X"832a7081",
X"06515155",
X"5573802e",
X"8638880b",
X"a0163489",
X"3d0d04f4",
X"3d0d02bb",
X"05330284",
X"05bf0533",
X"5d5d800b",
X"83cb980b",
X"83cb940b",
X"8c117271",
X"8814755c",
X"5a5b5f5c",
X"595b5883",
X"15335372",
X"802e8188",
X"38733353",
X"7c732e09",
X"810680fc",
X"38811433",
X"537b732e",
X"09810680",
X"ef387508",
X"83cb8c08",
X"2e098106",
X"80e23880",
X"567581c4",
X"2983cb9c",
X"11703383",
X"1e335b57",
X"55537478",
X"2e098106",
X"973883cb",
X"a0130879",
X"082e0981",
X"068a3881",
X"14335274",
X"51fef83f",
X"81167081",
X"ff065753",
X"8f7627c5",
X"38807708",
X"54547274",
X"2e913876",
X"51841308",
X"53722d83",
X"c0800881",
X"ff065480",
X"0b831b34",
X"7353a939",
X"811881c4",
X"1681c416",
X"81c41981",
X"c41f81c4",
X"1e81c41d",
X"6081c405",
X"415d5e5f",
X"59565658",
X"8f7825fe",
X"ca388053",
X"7283c080",
X"0c8e3d0d",
X"04f83d0d",
X"02ae0522",
X"7d595780",
X"56815580",
X"54865381",
X"80527a51",
X"f4ee3f83",
X"c0800881",
X"ff0683c0",
X"800c8a3d",
X"0d04f73d",
X"0d02b205",
X"22028405",
X"b7053360",
X"5a5b5780",
X"56825579",
X"54865381",
X"80527b51",
X"f4be3f83",
X"c0800881",
X"ff0683c0",
X"800c8b3d",
X"0d04f83d",
X"0d02af05",
X"33598058",
X"80578056",
X"80557854",
X"89538052",
X"7a51f494",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8a3d0d04",
X"ffb83d0d",
X"80cb3d08",
X"705381f3",
X"d85256fe",
X"aadc3f83",
X"c0800880",
X"f3387551",
X"fea4c73f",
X"83ffff0b",
X"83c08008",
X"2580e138",
X"7551fea4",
X"c63f83c0",
X"80085583",
X"c0800880",
X"cf388280",
X"5383c080",
X"08528a3d",
X"705257fe",
X"e69d3f74",
X"527551fe",
X"a3d73f80",
X"5980ca3d",
X"fdfc0554",
X"82805376",
X"527551fe",
X"a1de3f81",
X"15557488",
X"802e0981",
X"06e13880",
X"527551fe",
X"a3af3f80",
X"0b83e3d8",
X"0c7583e3",
X"d40c8739",
X"800b83e3",
X"d40c80ca",
X"3d0d04ff",
X"3d0d7370",
X"08535102",
X"93053372",
X"34700881",
X"05710c83",
X"3d0d04ff",
X"b83d0d80",
X"cb3d7070",
X"84055208",
X"585683e3",
X"d408802e",
X"80fa388a",
X"3d705a76",
X"55775481",
X"e9cb5380",
X"cb3dfdfc",
X"055255fe",
X"cfed3f80",
X"5280ca3d",
X"fdfc0551",
X"ffad3f83",
X"e3d80852",
X"83e3d408",
X"51fea2b5",
X"3f805874",
X"51fecdb3",
X"3f80ca3d",
X"fdf80554",
X"83c08008",
X"53745283",
X"e3d40851",
X"fea0b13f",
X"83e3d808",
X"1883e3d8",
X"0c80ca3d",
X"fdf80554",
X"815381f3",
X"e45283e3",
X"d40851fe",
X"a0923f83",
X"e3d80818",
X"83e3d80c",
X"80ca3d0d",
X"04000000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002d46",
X"00002d87",
X"00002da9",
X"00002dcb",
X"00002df1",
X"00002df1",
X"00002df1",
X"00002df1",
X"00002e62",
X"00002eb3",
X"00002ebd",
X"00004492",
X"00004eb2",
X"00004f7b",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3f00",
X"0c0c4000",
X"0a0a4100",
X"0b0b4100",
X"07074100",
X"0a0b4300",
X"080b4200",
X"06060004",
X"04044500",
X"05054400",
X"0e0f2900",
X"08080004",
X"09090004",
X"0a0f4300",
X"090f4200",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"0000615f",
X"00006466",
X"00006272",
X"00006466",
X"000062af",
X"00006300",
X"0000633f",
X"00006348",
X"00006466",
X"00006466",
X"00006466",
X"00006466",
X"00006351",
X"00006359",
X"00006360",
X"00006566",
X"0000665f",
X"00006773",
X"00006a69",
X"00006a84",
X"00006a70",
X"00006a84",
X"00006a8b",
X"00006a96",
X"00006a9d",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"25782e48",
X"75622e20",
X"25642070",
X"6f727473",
X"00000000",
X"25782e48",
X"49440000",
X"204d6f75",
X"73650000",
X"204b6579",
X"626f6172",
X"64000000",
X"204a6f79",
X"73746963",
X"6b3a2564",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"43505520",
X"54757262",
X"6f3a2564",
X"78000000",
X"44726976",
X"65205475",
X"72626f3a",
X"25730000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"526f7461",
X"74652055",
X"5342206a",
X"6f797374",
X"69636b73",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"66726565",
X"7a65722e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"4d454d00",
X"5374616e",
X"64617264",
X"00000000",
X"46617374",
X"28362900",
X"46617374",
X"28352900",
X"46617374",
X"28342900",
X"46617374",
X"28332900",
X"46617374",
X"28322900",
X"46617374",
X"28312900",
X"46617374",
X"28302900",
X"2f757362",
X"2e6c6f67",
X"00000000",
X"0a000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00007898",
X"0000789c",
X"000078a4",
X"000078b0",
X"000078bc",
X"000078c8",
X"000078d4",
X"000078d8",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00000028",
X"00000006",
X"00000005",
X"00000004",
X"00000003",
X"00000002",
X"00000001",
X"00000000",
X"00007994",
X"000079a0",
X"000079a8",
X"000079b0",
X"000079b8",
X"000079c0",
X"000079c8",
X"000079d0",
X"000077f0",
X"00007638",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"69383030",
X"00000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
