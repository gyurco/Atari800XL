
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81d3",
X"c8738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81da",
X"e00c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757580f3",
X"bb2d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7580f2fa",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80dbf104",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"775193c4",
X"3f83c080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3381dae8",
X"0b81dae8",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"52775192",
X"f33f83c0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583c0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"55b3a83f",
X"83c08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"811451b2",
X"c03f83c0",
X"80083070",
X"83c08008",
X"07802583",
X"c0800c53",
X"863d0d04",
X"fc3d0d76",
X"70525599",
X"e03f83c0",
X"80085481",
X"5383c080",
X"0880c738",
X"745199a3",
X"3f83c080",
X"080b0b81",
X"d8dc5383",
X"c0800852",
X"53ff8f3f",
X"83c08008",
X"a5380b0b",
X"81d8e052",
X"7251fefe",
X"3f83c080",
X"0894380b",
X"0b81d8e4",
X"527251fe",
X"ed3f83c0",
X"8008802e",
X"83388154",
X"73537283",
X"c0800c86",
X"3d0d04fd",
X"3d0d7570",
X"525498f9",
X"3f815383",
X"c0800898",
X"38735198",
X"c23f83c0",
X"b0085283",
X"c0800851",
X"feb43f83",
X"c0800853",
X"7283c080",
X"0c853d0d",
X"04df3d0d",
X"a43d0870",
X"525e8ee7",
X"3f83c080",
X"0833953d",
X"56547396",
X"3881ddf8",
X"527451b1",
X"9a3f9a39",
X"7d527851",
X"91e83f84",
X"e3397d51",
X"8ecd3f83",
X"c0800852",
X"74518dfd",
X"3f804380",
X"42804180",
X"4083c0b8",
X"0852943d",
X"70525d94",
X"d03f83c0",
X"80085980",
X"0b83c080",
X"08555b83",
X"c080087b",
X"2e943881",
X"1b74525b",
X"97d23f83",
X"c0800854",
X"83c08008",
X"ee38805a",
X"ff5f7909",
X"709f2c7b",
X"065b547a",
X"7a248438",
X"ff1b5af6",
X"1a700970",
X"9f2c7206",
X"7bff125a",
X"5a525555",
X"80752595",
X"38765197",
X"973f83c0",
X"800876ff",
X"18585557",
X"738024ed",
X"38747f2e",
X"873880c2",
X"fa3f745f",
X"78ff1b70",
X"585d5880",
X"7a259538",
X"775196ec",
X"3f83c080",
X"0876ff18",
X"58555873",
X"8024ed38",
X"800b83c7",
X"d00c800b",
X"83c8840c",
X"0b0b81d8",
X"e8518bbe",
X"3f81800b",
X"83c8840c",
X"0b0b81d8",
X"f0518bae",
X"3fa80b83",
X"c7d00c76",
X"802e80e8",
X"3883c7d0",
X"08777932",
X"70307072",
X"07802570",
X"872b83c8",
X"840c5156",
X"78535656",
X"969f3f83",
X"c0800880",
X"2e8a380b",
X"0b81d8f8",
X"518af33f",
X"765195df",
X"3f83c080",
X"08520b0b",
X"81da8451",
X"8ae03f76",
X"5195e53f",
X"83c08008",
X"83c7d008",
X"55577574",
X"258638a8",
X"1656f739",
X"7583c7d0",
X"0c86f076",
X"24ff9438",
X"87980b83",
X"c7d00c77",
X"802eb738",
X"7751959b",
X"3f83c080",
X"08785255",
X"95bb3f0b",
X"0b81d980",
X"5483c080",
X"088f3887",
X"39807634",
X"81d8390b",
X"0b81d8fc",
X"54745373",
X"520b0b81",
X"d8d05189",
X"f93f8054",
X"0b0b81da",
X"dc5189ee",
X"3f811454",
X"73a82e09",
X"8106ed38",
X"868da051",
X"beef3f80",
X"52903d70",
X"525780e1",
X"b93f8352",
X"765180e1",
X"b13f6281",
X"91386180",
X"2e80fd38",
X"7b5473ff",
X"2e963878",
X"802e818c",
X"38785194",
X"b73f83c0",
X"8008ff15",
X"5559e739",
X"78802e80",
X"f7387851",
X"94b33f83",
X"c0800880",
X"2efbfd38",
X"785193fb",
X"3f83c080",
X"08520b0b",
X"81d8d851",
X"abda3f83",
X"c08008a3",
X"387c51ad",
X"923f83c0",
X"80085574",
X"ff165654",
X"807425ae",
X"38741d70",
X"33555673",
X"af2efec5",
X"38e93978",
X"5193ba3f",
X"83c08008",
X"527c51ac",
X"ca3f8f39",
X"7f882960",
X"10057a05",
X"61055afb",
X"fd396280",
X"2efbbe38",
X"80527651",
X"80e08f3f",
X"a33d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"842a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"a80b9088",
X"b834b80b",
X"9088b834",
X"7083c080",
X"0c823d0d",
X"04803d0d",
X"9088b833",
X"7081ff06",
X"70852a81",
X"32708106",
X"51515151",
X"70802e8d",
X"38980b90",
X"88b834b8",
X"0b9088b8",
X"347083c0",
X"800c823d",
X"0d04930b",
X"9088bc34",
X"ff0b9088",
X"a83404ff",
X"3d0d028f",
X"05335280",
X"0b9088bc",
X"348a51bc",
X"b43fdf3f",
X"80f80b90",
X"88a03480",
X"0b908888",
X"34fa1252",
X"71908880",
X"34800b90",
X"88983471",
X"90889034",
X"9088b852",
X"807234b8",
X"7234833d",
X"0d04803d",
X"0d028b05",
X"33517090",
X"88b434fe",
X"bf3f83c0",
X"8008802e",
X"f638823d",
X"0d04803d",
X"0d853980",
X"c6873ffe",
X"d83f83c0",
X"8008802e",
X"f2389088",
X"b4337081",
X"ff0683c0",
X"800c5182",
X"3d0d0480",
X"3d0da30b",
X"9088bc34",
X"ff0b9088",
X"a8349088",
X"b851a871",
X"34b87134",
X"823d0d04",
X"803d0d90",
X"88bc3370",
X"81c00670",
X"30708025",
X"83c0800c",
X"51515182",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067083",
X"2a813270",
X"81065151",
X"51517080",
X"2ee838b0",
X"0b9088b8",
X"34b80b90",
X"88b83482",
X"3d0d0480",
X"3d0d9080",
X"ac088106",
X"83c0800c",
X"823d0d04",
X"fd3d0d75",
X"77545480",
X"73259438",
X"73708105",
X"55335281",
X"d9845185",
X"a13fff13",
X"53e93985",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"80de8f3f",
X"83c08008",
X"7a27ed38",
X"74802e80",
X"e0387452",
X"755180dd",
X"f93f83c0",
X"80087553",
X"76525480",
X"ddfc3f83",
X"c080087a",
X"53755256",
X"80dddf3f",
X"83c08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"c08008c2",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9c",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fbfd3f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd13f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbad3f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83c0900c",
X"7183c094",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383c090",
X"085283c0",
X"940851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"99e65351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fd3d",
X"0d757052",
X"54a3c43f",
X"83c08008",
X"14537274",
X"2e9238ff",
X"13703353",
X"5371af2e",
X"098106ee",
X"38811353",
X"7283c080",
X"0c853d0d",
X"04fd3d0d",
X"75777053",
X"5454c73f",
X"83c08008",
X"732ea138",
X"83c08008",
X"733152ff",
X"125271ff",
X"2e8f3872",
X"70810554",
X"33747081",
X"055634eb",
X"39ff1454",
X"80743485",
X"3d0d0480",
X"3d0d7251",
X"ff903f82",
X"3d0d0471",
X"83c0800c",
X"04803d0d",
X"72518071",
X"34810bbc",
X"120c800b",
X"80c0120c",
X"823d0d04",
X"800b83c2",
X"e408248a",
X"38a4ae3f",
X"ff0b83c2",
X"e40c800b",
X"83c0800c",
X"04ff3d0d",
X"735283c0",
X"c008722e",
X"8d38d93f",
X"71519699",
X"3f7183c0",
X"c00c833d",
X"0d04f43d",
X"0d7e6062",
X"5c5a5581",
X"54bc1508",
X"81913874",
X"51cf3f79",
X"58807a25",
X"80f73883",
X"c3940870",
X"892a5783",
X"ff067884",
X"80723156",
X"56577378",
X"25833873",
X"557583c2",
X"e4082e84",
X"38ff893f",
X"83c2e408",
X"8025a638",
X"75892b51",
X"98dc3f83",
X"c394088f",
X"3dfc1155",
X"5c548152",
X"f81b5196",
X"c63f7614",
X"83c3940c",
X"7583c2e4",
X"0c745376",
X"527851a2",
X"df3f83c0",
X"800883c3",
X"94081683",
X"c3940c78",
X"7631761b",
X"5b595677",
X"8024ff8b",
X"38617a71",
X"0c547554",
X"75802e83",
X"38815473",
X"83c0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"9b3f7651",
X"feaf3f86",
X"3dfc0553",
X"78527751",
X"95e93f79",
X"75710c54",
X"83c08008",
X"5483c080",
X"08802e83",
X"38815473",
X"83c0800c",
X"863d0d04",
X"fe3d0d75",
X"83c2e408",
X"53538072",
X"24893871",
X"732e8438",
X"fdd63f74",
X"51fdea3f",
X"725197ae",
X"3f83c080",
X"085283c0",
X"8008802e",
X"83388152",
X"7183c080",
X"0c843d0d",
X"04803d0d",
X"7280c011",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d72bc11",
X"0883c080",
X"0c51823d",
X"0d0480c4",
X"0b83c080",
X"0c04fd3d",
X"0d757771",
X"54705355",
X"539f9c3f",
X"82c81308",
X"bc150c82",
X"c0130880",
X"c0150cfc",
X"eb3f7351",
X"93ab3f73",
X"83c0c00c",
X"83c08008",
X"5383c080",
X"08802e83",
X"38815372",
X"83c0800c",
X"853d0d04",
X"fd3d0d75",
X"775553fc",
X"bf3f7280",
X"2ea538bc",
X"13085273",
X"519ea63f",
X"83c08008",
X"8f387752",
X"7251ff9a",
X"3f83c080",
X"08538a39",
X"82cc1308",
X"53d83981",
X"537283c0",
X"800c853d",
X"0d04fe3d",
X"0dff0b83",
X"c2e40c74",
X"83c0c40c",
X"7583c2e0",
X"0c9f933f",
X"83c08008",
X"81ff0652",
X"81537199",
X"3883c2fc",
X"518e943f",
X"83c08008",
X"5283c080",
X"08802e83",
X"38725271",
X"537283c0",
X"800c843d",
X"0d04fa3d",
X"0d787a82",
X"c4120882",
X"c4120870",
X"72245956",
X"56575773",
X"732e0981",
X"06913880",
X"c0165280",
X"c017519c",
X"973f83c0",
X"80085574",
X"83c0800c",
X"883d0d04",
X"f63d0d7c",
X"5b807b71",
X"5c54577a",
X"772e8c38",
X"811a82cc",
X"1408545a",
X"72f63880",
X"5980d939",
X"7a548157",
X"80707b7b",
X"315a5755",
X"ff185374",
X"732580c1",
X"3882cc14",
X"08527351",
X"ff8c3f80",
X"0b83c080",
X"0825a138",
X"82cc1408",
X"82cc1108",
X"82cc160c",
X"7482cc12",
X"0c537580",
X"2e863872",
X"82cc170c",
X"72548057",
X"7382cc15",
X"08811757",
X"5556ffb8",
X"39811959",
X"800bff1b",
X"54547873",
X"25833881",
X"54768132",
X"70750651",
X"5372ff90",
X"388c3d0d",
X"04f73d0d",
X"7b7d5a5a",
X"82d05283",
X"c2e00851",
X"80d1973f",
X"83c08008",
X"57f9e13f",
X"795283c2",
X"e85195b5",
X"3f83c080",
X"08548053",
X"83c08008",
X"732e0981",
X"06828338",
X"83c0c408",
X"0b0b81d8",
X"d8537052",
X"569bd43f",
X"0b0b81d8",
X"d85280c0",
X"16519bc7",
X"3f75bc17",
X"0c7382c0",
X"170c810b",
X"82c4170c",
X"810b82c8",
X"170c7382",
X"cc170cff",
X"1782d017",
X"55578191",
X"3983c0d0",
X"3370822a",
X"70810651",
X"54557281",
X"80387481",
X"2a810658",
X"7780f638",
X"74842a81",
X"0682c415",
X"0c83c0d0",
X"33810682",
X"c8150c79",
X"5273519a",
X"ee3f7351",
X"9b853f83",
X"c0800814",
X"53af7370",
X"81055534",
X"72bc150c",
X"83c0d152",
X"72519acf",
X"3f83c0c8",
X"0882c015",
X"0c83c0de",
X"5280c014",
X"519abc3f",
X"78802e8d",
X"38735178",
X"2d83c080",
X"08802e99",
X"387782cc",
X"150c7580",
X"2e863873",
X"82cc170c",
X"7382d015",
X"ff195955",
X"5676802e",
X"9b3883c0",
X"c85283c2",
X"e85194ab",
X"3f83c080",
X"088a3883",
X"c0d13353",
X"72fed238",
X"78802e89",
X"3883c0c4",
X"0851fcb8",
X"3f83c0c4",
X"08537283",
X"c0800c8b",
X"3d0d04ff",
X"3d0d8052",
X"7351fdb5",
X"3f833d0d",
X"04f03d0d",
X"62705254",
X"f6903f83",
X"c0800874",
X"53873d70",
X"535555f6",
X"b03ff790",
X"3f7351d3",
X"3f635374",
X"5283c080",
X"0851fab8",
X"3f923d0d",
X"047183c0",
X"800c0480",
X"c01283c0",
X"800c0480",
X"3d0d7282",
X"c0110883",
X"c0800c51",
X"823d0d04",
X"803d0d72",
X"82cc1108",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"7282c411",
X"0883c080",
X"0c51823d",
X"0d04f93d",
X"0d7983c0",
X"98085757",
X"81772781",
X"96387688",
X"17082781",
X"8e387533",
X"5574822e",
X"89387483",
X"2eb33880",
X"fe397454",
X"761083fe",
X"06537688",
X"2a8c1708",
X"0552893d",
X"fc055199",
X"c13f83c0",
X"800880df",
X"38029d05",
X"33893d33",
X"71882b07",
X"565680d1",
X"39845476",
X"822b83fc",
X"06537687",
X"2a8c1708",
X"0552893d",
X"fc055199",
X"913f83c0",
X"8008b038",
X"029f0533",
X"0284059e",
X"05337198",
X"2b71902b",
X"07028c05",
X"9d053370",
X"882b7207",
X"8d3d3371",
X"80fffffe",
X"80060751",
X"52535758",
X"56833981",
X"557483c0",
X"800c893d",
X"0d04fb3d",
X"0d83c098",
X"08fe1988",
X"1208fe05",
X"55565480",
X"56747327",
X"8d388214",
X"33757129",
X"94160805",
X"57537583",
X"c0800c87",
X"3d0d04fc",
X"3d0d7652",
X"800b83c0",
X"98087033",
X"51525370",
X"832e0981",
X"06913895",
X"12339413",
X"3371982b",
X"71902b07",
X"5555519b",
X"12339a13",
X"3371882b",
X"07740783",
X"c0800c55",
X"863d0d04",
X"fc3d0d76",
X"83c09808",
X"55558075",
X"23881508",
X"5372812e",
X"88388814",
X"08732685",
X"388152b2",
X"39729038",
X"73335271",
X"832e0981",
X"06853890",
X"14085372",
X"8c160c72",
X"802e8d38",
X"7251fed6",
X"3f83c080",
X"08528539",
X"90140852",
X"7190160c",
X"80527183",
X"c0800c86",
X"3d0d04fa",
X"3d0d7883",
X"c0980871",
X"22810570",
X"83ffff06",
X"57545755",
X"73802e88",
X"38901508",
X"53728638",
X"835280e7",
X"39738f06",
X"527180da",
X"38811390",
X"160c8c15",
X"08537290",
X"38830b84",
X"17225752",
X"73762780",
X"c638bf39",
X"821633ff",
X"0574842a",
X"065271b2",
X"387251fc",
X"b13f8152",
X"7183c080",
X"0827a838",
X"835283c0",
X"80088817",
X"08279c38",
X"83c08008",
X"8c160c83",
X"c0800851",
X"fdbc3f83",
X"c0800890",
X"160c7375",
X"23805271",
X"83c0800c",
X"883d0d04",
X"f23d0d60",
X"6264585e",
X"5b753355",
X"74a02e09",
X"81068838",
X"81167044",
X"56ef3962",
X"70335656",
X"74af2e09",
X"81068438",
X"81164380",
X"0b881c0c",
X"62703351",
X"55749f26",
X"91387a51",
X"fdd23f83",
X"c0800856",
X"807d3483",
X"8139933d",
X"841c0870",
X"58595f8a",
X"55a07670",
X"81055834",
X"ff155574",
X"ff2e0981",
X"06ef3880",
X"705a5c88",
X"7f085f5a",
X"7b811d70",
X"81ff0660",
X"13703370",
X"af327030",
X"a0732771",
X"80250751",
X"51525b53",
X"5e575574",
X"80e73876",
X"ae2e0981",
X"06833881",
X"55787a27",
X"75075574",
X"802e9f38",
X"79883270",
X"3078ae32",
X"70307073",
X"079f2a53",
X"51575156",
X"75bb3888",
X"598b5aff",
X"ab397698",
X"2b557480",
X"25873881",
X"d2d81733",
X"57ff9f17",
X"55749926",
X"8938e017",
X"7081ff06",
X"58557881",
X"1a7081ff",
X"06721b53",
X"5b575576",
X"7534fef8",
X"397b1e7f",
X"0c805576",
X"a0268338",
X"8155748b",
X"19347a51",
X"fc823f83",
X"c0800880",
X"f538a054",
X"7a227085",
X"2b83e006",
X"5455901b",
X"08527c51",
X"93cc3f83",
X"c0800857",
X"83c08008",
X"8181387c",
X"33557480",
X"2e80f438",
X"8b1d3370",
X"832a7081",
X"06515656",
X"74b4388b",
X"7d841d08",
X"83c08008",
X"595b5b58",
X"ff185877",
X"ff2e9a38",
X"79708105",
X"5b337970",
X"81055b33",
X"71713152",
X"56567580",
X"2ee23886",
X"3975802e",
X"96387a51",
X"fbe53fff",
X"863983c0",
X"80085683",
X"c08008b6",
X"38833976",
X"56841b08",
X"8b113351",
X"5574a738",
X"8b1d3370",
X"842a7081",
X"06515656",
X"74893883",
X"56943981",
X"5690397c",
X"51fa943f",
X"83c08008",
X"881c0cfd",
X"81397583",
X"c0800c90",
X"3d0d04f8",
X"3d0d7a7c",
X"59578254",
X"83fe5377",
X"52765192",
X"913f8356",
X"83c08008",
X"80ec3881",
X"17337733",
X"71882b07",
X"56568256",
X"7482d4d5",
X"2e098106",
X"80d43875",
X"54b65377",
X"52765191",
X"e53f83c0",
X"80089838",
X"81173377",
X"3371882b",
X"0783c080",
X"08525656",
X"748182c6",
X"2eac3882",
X"5480d253",
X"77527651",
X"91bc3f83",
X"c0800898",
X"38811733",
X"77337188",
X"2b0783c0",
X"80085256",
X"56748182",
X"c62e8338",
X"81567583",
X"c0800c8a",
X"3d0d04eb",
X"3d0d675a",
X"800b83c0",
X"980c90de",
X"3f83c080",
X"08810655",
X"82567483",
X"ef387475",
X"538f3d70",
X"535759fe",
X"ca3f83c0",
X"800881ff",
X"06577681",
X"2e098106",
X"80d43890",
X"5483be53",
X"74527551",
X"90d03f83",
X"c0800880",
X"c9388f3d",
X"33557480",
X"2e80c938",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"0770587b",
X"575e525e",
X"575957fd",
X"ee3f83c0",
X"800881ff",
X"06577683",
X"2e098106",
X"86388156",
X"82f23976",
X"802e8638",
X"865682e8",
X"39a4548d",
X"53785275",
X"518fe73f",
X"815683c0",
X"800882d4",
X"3802be05",
X"33028405",
X"bd053371",
X"882b0759",
X"5d77ab38",
X"0280ce05",
X"33028405",
X"80cd0533",
X"71982b71",
X"902b0797",
X"3d337088",
X"2b720702",
X"940580cb",
X"05337107",
X"54525e57",
X"595602b7",
X"05337871",
X"29028805",
X"b6053302",
X"8c05b505",
X"3371882b",
X"07701d70",
X"7f8c050c",
X"5f595759",
X"5d8e3d33",
X"821b3402",
X"b9053390",
X"3d337188",
X"2b075a5c",
X"78841b23",
X"02bb0533",
X"028405ba",
X"05337188",
X"2b07565c",
X"74ab3802",
X"80ca0533",
X"02840580",
X"c9053371",
X"982b7190",
X"2b07963d",
X"3370882b",
X"72070294",
X"0580c705",
X"33710751",
X"5253575e",
X"5c747631",
X"78317984",
X"2a903d33",
X"54717131",
X"53565680",
X"c1fc3f83",
X"c0800882",
X"0570881c",
X"0c83c080",
X"08e08a05",
X"56567483",
X"dffe2683",
X"38825783",
X"fff67627",
X"85388357",
X"89398656",
X"76802e80",
X"db38767a",
X"3476832e",
X"098106b0",
X"380280d6",
X"05330284",
X"0580d505",
X"3371982b",
X"71902b07",
X"993d3370",
X"882b7207",
X"02940580",
X"d3053371",
X"077f9005",
X"0c525e57",
X"58568639",
X"771b901b",
X"0c841a22",
X"8c1b0819",
X"71842a05",
X"941c0c5d",
X"800b811b",
X"347983c0",
X"980c8056",
X"7583c080",
X"0c973d0d",
X"04e93d0d",
X"83c09808",
X"56855475",
X"802e8182",
X"38800b81",
X"1734993d",
X"e011466a",
X"548a3d70",
X"5458ec05",
X"51f6e53f",
X"83c08008",
X"5483c080",
X"0880df38",
X"893d3354",
X"73802e91",
X"3802ab05",
X"3370842a",
X"81065155",
X"74802e86",
X"38835480",
X"c1397651",
X"f4893f83",
X"c08008a0",
X"170c02bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"3371079c",
X"1c0c5278",
X"981b0c53",
X"56595781",
X"0b811734",
X"74547383",
X"c0800c99",
X"3d0d04f5",
X"3d0d7d7f",
X"617283c0",
X"98085a5d",
X"5d595c80",
X"7b0c8557",
X"75802e81",
X"e0388116",
X"33810655",
X"84577480",
X"2e81d238",
X"91397481",
X"17348639",
X"800b8117",
X"34815781",
X"c0399c16",
X"08981708",
X"31557478",
X"27833874",
X"5877802e",
X"81a93898",
X"16087083",
X"ff065657",
X"7480cf38",
X"821633ff",
X"0577892a",
X"067081ff",
X"065a5578",
X"a0387687",
X"38a01608",
X"558d39a4",
X"160851f0",
X"e93f83c0",
X"80085581",
X"7527ffa8",
X"3874a417",
X"0ca41608",
X"51f2833f",
X"83c08008",
X"5583c080",
X"08802eff",
X"893883c0",
X"800819a8",
X"170c9816",
X"0883ff06",
X"84807131",
X"51557775",
X"27833877",
X"557483ff",
X"ff065498",
X"160883ff",
X"0653a816",
X"08527957",
X"7b83387b",
X"5776518a",
X"8d3f83c0",
X"8008fed0",
X"38981608",
X"1598170c",
X"741a7876",
X"317c0817",
X"7d0c595a",
X"fed33980",
X"577683c0",
X"800c8d3d",
X"0d04fa3d",
X"0d7883c0",
X"98085556",
X"85557380",
X"2e81e138",
X"81143381",
X"06538455",
X"72802e81",
X"d3389c14",
X"08537276",
X"27833872",
X"56981408",
X"57800b98",
X"150c7580",
X"2e81b738",
X"82143370",
X"892b5653",
X"76802eb5",
X"387452ff",
X"1651bcfe",
X"3f83c080",
X"08ff1876",
X"54705358",
X"53bcef3f",
X"83c08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed83f83",
X"c0800853",
X"810b83c0",
X"8008278b",
X"38881408",
X"83c08008",
X"26883880",
X"0b811534",
X"b03983c0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc73f",
X"83c08008",
X"8c3883c0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683c0",
X"800805a8",
X"150c8055",
X"7483c080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83c09808",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1d13f",
X"83c08008",
X"5583c080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef7",
X"3f83c080",
X"0888170c",
X"7551efa8",
X"3f83c080",
X"08557483",
X"c0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683c0",
X"9808802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f73f83c0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"86983f83",
X"c0800841",
X"83c08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"ede13f83",
X"c0800841",
X"83c08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"83a53f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f23f83c0",
X"80088332",
X"70307072",
X"079f2c83",
X"c0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"81b13f75",
X"83c0800c",
X"9e3d0d04",
X"fd3d0d75",
X"77535473",
X"33517089",
X"38713351",
X"70802ea1",
X"38733372",
X"33525372",
X"71278538",
X"ff519439",
X"70732785",
X"3881518b",
X"39811481",
X"135354d3",
X"39805170",
X"83c0800c",
X"853d0d04",
X"fd3d0d75",
X"77545472",
X"337081ff",
X"06525270",
X"802ea338",
X"7181ff06",
X"8114ffbf",
X"12535452",
X"70992689",
X"38a01270",
X"81ff0653",
X"51717470",
X"81055634",
X"d2398074",
X"34853d0d",
X"04ffbd3d",
X"0d80c63d",
X"0852a53d",
X"705254ff",
X"b33f80c7",
X"3d085285",
X"3d705253",
X"ffa63f72",
X"527351fe",
X"df3f80c5",
X"3d0d04fe",
X"3d0d7476",
X"53537170",
X"81055333",
X"51707370",
X"81055534",
X"70f03884",
X"3d0d04fe",
X"3d0d7452",
X"80723352",
X"5370732e",
X"8d388112",
X"81147133",
X"53545270",
X"f5387283",
X"c0800c84",
X"3d0d04fc",
X"3d0d7655",
X"7483c3a8",
X"082eaf38",
X"80537451",
X"87c13f83",
X"c0800881",
X"ff06ff14",
X"7081ff06",
X"7230709f",
X"2a515255",
X"53547280",
X"2e843871",
X"dd3873fe",
X"387483c3",
X"a80c863d",
X"0d04ff3d",
X"0dff0b83",
X"c3a80c84",
X"a53f8151",
X"87853f83",
X"c0800881",
X"ff065271",
X"ee3881d3",
X"3f7183c0",
X"800c833d",
X"0d04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"823f7280",
X"2ea03883",
X"c3bc1433",
X"75708105",
X"57348114",
X"7083ffff",
X"06ff1570",
X"83ffff06",
X"56525552",
X"dd39800b",
X"83c0800c",
X"863d0d04",
X"fc3d0d76",
X"787a1156",
X"53558053",
X"71742e93",
X"38721551",
X"703383c3",
X"bc133481",
X"12811454",
X"52ea3980",
X"0b83c080",
X"0c863d0d",
X"04fd3d0d",
X"905483c3",
X"a8085186",
X"f43f83c0",
X"800881ff",
X"06ff1571",
X"30713070",
X"73079f2a",
X"729f2a06",
X"52555255",
X"5372db38",
X"853d0d04",
X"803d0d83",
X"c3b40810",
X"83c3ac08",
X"079080a8",
X"0c823d0d",
X"04800b83",
X"c3b40ce4",
X"3f04810b",
X"83c3b40c",
X"db3f04ed",
X"3f047183",
X"c3b00c04",
X"803d0d80",
X"51f43f81",
X"0b83c3b4",
X"0c810b83",
X"c3ac0cff",
X"bb3f823d",
X"0d04803d",
X"0d723070",
X"74078025",
X"83c3ac0c",
X"51ffa53f",
X"823d0d04",
X"803d0d02",
X"8b053390",
X"80a40c90",
X"80a80870",
X"81065151",
X"70f53890",
X"80a40870",
X"81ff0683",
X"c0800c51",
X"823d0d04",
X"803d0d81",
X"ff51d13f",
X"83c08008",
X"81ff0683",
X"c0800c82",
X"3d0d0480",
X"3d0d7390",
X"2b730790",
X"80b40c82",
X"3d0d0404",
X"fb3d0d78",
X"0284059f",
X"05337098",
X"2b555755",
X"7280259b",
X"387580ff",
X"06568052",
X"80f751e0",
X"3f83c080",
X"0881ff06",
X"54738126",
X"80ff3880",
X"51fee73f",
X"ffa23f81",
X"51fedf3f",
X"ff9a3f75",
X"51feed3f",
X"74982a51",
X"fee63f74",
X"902a7081",
X"ff065253",
X"feda3f74",
X"882a7081",
X"ff065253",
X"fece3f74",
X"81ff0651",
X"fec63f81",
X"557580c0",
X"2e098106",
X"86388195",
X"558d3975",
X"80c82e09",
X"81068438",
X"81875574",
X"51fea53f",
X"8a55fec8",
X"3f83c080",
X"0881ff06",
X"70982b54",
X"54728025",
X"8c38ff15",
X"7081ff06",
X"565374e2",
X"387383c0",
X"800c873d",
X"0d04fa3d",
X"0dfdc53f",
X"8051fdda",
X"3f8a54fe",
X"933fff14",
X"7081ff06",
X"555373f3",
X"38737453",
X"5580c051",
X"fea63f83",
X"c0800881",
X"ff065473",
X"812e0981",
X"06829f38",
X"83aa5280",
X"c851fe8c",
X"3f83c080",
X"0881ff06",
X"5372812e",
X"09810681",
X"a8387454",
X"873d7411",
X"5456fdc8",
X"3f83c080",
X"08733481",
X"147081ff",
X"06555383",
X"7427e538",
X"029a0533",
X"5372812e",
X"09810681",
X"d938029b",
X"05335380",
X"ce905472",
X"81aa2e8d",
X"3881c739",
X"80e4518a",
X"cc3fff14",
X"5473802e",
X"81b83882",
X"0a5281e9",
X"51fda53f",
X"83c08008",
X"81ff0653",
X"72de3872",
X"5280fa51",
X"fd923f83",
X"c0800881",
X"ff065372",
X"81903872",
X"54731653",
X"fcd63f83",
X"c0800873",
X"34811470",
X"81ff0655",
X"53837427",
X"e838873d",
X"3370862a",
X"70810651",
X"54548c55",
X"7280e338",
X"845580de",
X"39745281",
X"e951fccc",
X"3f83c080",
X"0881ff06",
X"53825581",
X"e9568173",
X"27863873",
X"5580c156",
X"80ce9054",
X"8a3980e4",
X"5189be3f",
X"ff145473",
X"802ea938",
X"80527551",
X"fc9a3f83",
X"c0800881",
X"ff065372",
X"e1388480",
X"5280d051",
X"fc863f83",
X"c0800881",
X"ff065372",
X"802e8338",
X"80557483",
X"c3b83480",
X"51fb873f",
X"fbc23f88",
X"3d0d04fb",
X"3d0d7754",
X"800b83c3",
X"b8337083",
X"2a708106",
X"51555755",
X"72752e09",
X"81068538",
X"73892b54",
X"735280d1",
X"51fbbd3f",
X"83c08008",
X"81ff0653",
X"72bd3882",
X"b8c054fb",
X"833f83c0",
X"800881ff",
X"06537281",
X"ff2e0981",
X"068938ff",
X"145473e7",
X"389f3972",
X"81fe2e09",
X"81069638",
X"83c7bc52",
X"83c3bc51",
X"faed3ffa",
X"d33ffad0",
X"3f833981",
X"558051fa",
X"893ffac4",
X"3f7481ff",
X"0683c080",
X"0c873d0d",
X"04fb3d0d",
X"7783c3bc",
X"56548151",
X"f9ec3f83",
X"c3b83370",
X"832a7081",
X"06515456",
X"72853873",
X"892b5473",
X"5280d851",
X"fab63f83",
X"c0800881",
X"ff065372",
X"80e43881",
X"ff51f9d4",
X"3f81fe51",
X"f9ce3f84",
X"80537470",
X"81055633",
X"51f9c13f",
X"ff137083",
X"ffff0651",
X"5372eb38",
X"7251f9b0",
X"3f7251f9",
X"ab3ff9d0",
X"3f83c080",
X"089f0653",
X"a7885472",
X"852e8c38",
X"993980e4",
X"5186f63f",
X"ff1454f9",
X"b33f83c0",
X"800881ff",
X"2e843873",
X"e9388051",
X"f8e43ff9",
X"9f3f800b",
X"83c0800c",
X"873d0d04",
X"7183c7c0",
X"0c888080",
X"0b83c7bc",
X"0c848080",
X"0b83c7c4",
X"0c04fd3d",
X"0d777017",
X"557705ff",
X"1a535371",
X"ff2e9438",
X"73708105",
X"55335170",
X"73708105",
X"5534ff12",
X"52e93985",
X"3d0d04fc",
X"3d0d87a6",
X"81557433",
X"83c7c834",
X"a05483a0",
X"805383c7",
X"c0085283",
X"c7bc0851",
X"ffb83fa0",
X"5483a480",
X"5383c7c0",
X"085283c7",
X"bc0851ff",
X"a53f9054",
X"83a88053",
X"83c7c008",
X"5283c7bc",
X"0851ff92",
X"3fa05380",
X"5283c7c4",
X"0883a080",
X"055185ce",
X"3fa05380",
X"5283c7c4",
X"0883a480",
X"055185be",
X"3f905380",
X"5283c7c4",
X"0883a880",
X"055185ae",
X"3fff7534",
X"83a08054",
X"805383c7",
X"c0085283",
X"c7c40851",
X"fecc3f80",
X"d0805483",
X"b0805383",
X"c7c00852",
X"83c7c408",
X"51feb73f",
X"86e13fa2",
X"54805383",
X"c7c4088c",
X"80055281",
X"dbdc51fe",
X"a13f860b",
X"87a88334",
X"800b87a8",
X"8234800b",
X"87a09a34",
X"af0b87a0",
X"9634bf0b",
X"87a09734",
X"800b87a0",
X"98349f0b",
X"87a09934",
X"800b87a0",
X"9b34e00b",
X"87a88934",
X"a20b87a8",
X"8034830b",
X"87a48f34",
X"820b87a8",
X"8134863d",
X"0d04fd3d",
X"0d83a080",
X"54805383",
X"c7c40852",
X"83c7c008",
X"51fdbf3f",
X"80d08054",
X"83b08053",
X"83c7c408",
X"5283c7c0",
X"0851fdaa",
X"3fa05483",
X"a0805383",
X"c7c40852",
X"83c7c008",
X"51fd973f",
X"a05483a4",
X"805383c7",
X"c4085283",
X"c7c00851",
X"fd843f90",
X"5483a880",
X"5383c7c4",
X"085283c7",
X"c00851fc",
X"f13f83c7",
X"c83387a6",
X"8134853d",
X"0d04803d",
X"0d908090",
X"08810683",
X"c0800c82",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe067607",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"812c8106",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fd06",
X"76100772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087082",
X"2cbf0683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fe8306",
X"76822b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"882c8706",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f1ff",
X"0676882b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"708b2cbf",
X"0683c080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870f8",
X"8fff0676",
X"8b2b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087091",
X"2cbf0683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fc87ff",
X"ff067691",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870992c",
X"810683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"ffbf0a06",
X"76992b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80800870",
X"882c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"70892c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708a2c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708b",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8c2cbf06",
X"83c0800c",
X"51823d0d",
X"04fe3d0d",
X"7481e629",
X"872a9080",
X"a00c843d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"81055434",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727084",
X"05540cff",
X"1151f039",
X"843d0d04",
X"fe3d0d84",
X"80805380",
X"5288800a",
X"51ffb33f",
X"81808053",
X"80528280",
X"0a51c63f",
X"843d0d04",
X"803d0d81",
X"51fbfc3f",
X"72802e90",
X"388051fd",
X"fe3fcd3f",
X"83c7cc33",
X"51fdf43f",
X"8151fc8d",
X"3f8051fc",
X"883f8051",
X"fbd93f82",
X"3d0d04fd",
X"3d0d7552",
X"805480ff",
X"72258838",
X"810bff80",
X"135354ff",
X"bf125170",
X"99268638",
X"e012529e",
X"39ff9f12",
X"51997127",
X"9538d012",
X"e0137054",
X"54518971",
X"2788388f",
X"73278338",
X"80527380",
X"2e853881",
X"80125271",
X"81ff0683",
X"c0800c85",
X"3d0d0480",
X"3d0d84d8",
X"c0518071",
X"70810553",
X"347084e0",
X"c02e0981",
X"06f03882",
X"3d0d04fe",
X"3d0d0297",
X"053351ff",
X"863f83c0",
X"800881ff",
X"0683c7d0",
X"08545280",
X"73249b38",
X"83c88008",
X"137283c8",
X"84080753",
X"53717334",
X"83c7d008",
X"810583c7",
X"d00c843d",
X"0d04fa3d",
X"0d82800a",
X"1b558057",
X"883dfc05",
X"54795374",
X"527851cb",
X"d33f883d",
X"0d04fe3d",
X"0d83c7e8",
X"08527451",
X"d2b73f83",
X"c080088c",
X"38765375",
X"5283c7e8",
X"0851c73f",
X"843d0d04",
X"fe3d0d83",
X"c7e80853",
X"75527451",
X"ccf63f83",
X"c080088d",
X"38775376",
X"5283c7e8",
X"0851ffa2",
X"3f843d0d",
X"04fe3d0d",
X"83c7e808",
X"51cbea3f",
X"83c08008",
X"8180802e",
X"09810688",
X"3883c180",
X"80539b39",
X"83c7e808",
X"51cbce3f",
X"83c08008",
X"80d0802e",
X"09810693",
X"3883c1b0",
X"805383c0",
X"80085283",
X"c7e80851",
X"fed83f84",
X"3d0d0480",
X"3d0df9e4",
X"3f83c080",
X"08842981",
X"dc800570",
X"0883c080",
X"0c51823d",
X"0d04ed3d",
X"0d804480",
X"43804280",
X"4180705a",
X"5bfdd03f",
X"800b83c7",
X"d00c800b",
X"83c8840c",
X"81d9d051",
X"c6b83f81",
X"800b83c8",
X"840c81d9",
X"d451c6aa",
X"3f80d00b",
X"83c7d00c",
X"7830707a",
X"07802570",
X"872b83c8",
X"840c5155",
X"f8d53f83",
X"c0800852",
X"81d9dc51",
X"c6843f80",
X"f80b83c7",
X"d00c7881",
X"32703070",
X"72078025",
X"70872b83",
X"c8840c51",
X"5656feef",
X"3f83c080",
X"085281d9",
X"e851c5da",
X"3f81a00b",
X"83c7d00c",
X"78823270",
X"30707207",
X"80257087",
X"2b83c884",
X"0c515683",
X"c7e80852",
X"56c6f43f",
X"83c08008",
X"5281d9f0",
X"51c5ab3f",
X"81f00b83",
X"c7d00c81",
X"0b83c7d4",
X"5b5883c7",
X"d0088219",
X"7a327030",
X"70720780",
X"2570872b",
X"83c8840c",
X"51578e3d",
X"7055ff1b",
X"54575757",
X"9a953f79",
X"7084055b",
X"0851c6ab",
X"3f745483",
X"c0800853",
X"775281d9",
X"f851c4de",
X"3fa81783",
X"c7d00c81",
X"18587785",
X"2e098106",
X"ffb03883",
X"900b83c7",
X"d00c7887",
X"32703070",
X"72078025",
X"70872b83",
X"c8840c51",
X"5656f7fb",
X"3f81da88",
X"5583c080",
X"08802e8e",
X"3883c7e4",
X"0851c5d7",
X"3f83c080",
X"08557452",
X"81da9051",
X"c48c3f83",
X"e00b83c7",
X"d00c7888",
X"32703070",
X"72078025",
X"70872b83",
X"c8840c51",
X"5781da9c",
X"5255c3ea",
X"3f868da0",
X"51f8f63f",
X"8052913d",
X"7052559b",
X"c13f8352",
X"74519bba",
X"3f635574",
X"82fc3861",
X"19597880",
X"25853874",
X"59903988",
X"79258538",
X"88598739",
X"78882682",
X"db387882",
X"2b5581d4",
X"d8150804",
X"f5e93f83",
X"c0800861",
X"57557581",
X"2e098106",
X"893883c0",
X"80081055",
X"903975ff",
X"2e098106",
X"883883c0",
X"8008812c",
X"55907525",
X"85389055",
X"88397480",
X"24833881",
X"557451f5",
X"c33f8290",
X"39f5d53f",
X"83c08008",
X"61055574",
X"80258538",
X"80558839",
X"87752583",
X"38875574",
X"51f5ce3f",
X"81ee3960",
X"87386280",
X"2e81e538",
X"83c0b408",
X"83c0b00c",
X"8bdf0b83",
X"c0b80c83",
X"c7e80851",
X"ffb4ee3f",
X"fadf3f81",
X"c7396056",
X"80762599",
X"388af80b",
X"83c0b80c",
X"83c7c815",
X"70085255",
X"ffb4ce3f",
X"74085291",
X"39758025",
X"913883c7",
X"c8150851",
X"c3bf3f80",
X"52fd1951",
X"b8396280",
X"2e818d38",
X"83c7c815",
X"700883c7",
X"d408720c",
X"83c7d40c",
X"fd1a7053",
X"51558c82",
X"3f83c080",
X"08568051",
X"8bf83f83",
X"c0800852",
X"74518890",
X"3f755280",
X"5188893f",
X"80d63960",
X"55807525",
X"b83883c0",
X"bc0883c0",
X"b00c8bdf",
X"0b83c0b8",
X"0c83c7e4",
X"0851ffb3",
X"d83f83c7",
X"e40851ff",
X"b0f23f83",
X"c0800881",
X"ff067052",
X"55f4d93f",
X"74802e9c",
X"388155a0",
X"39748025",
X"933883c7",
X"e40851c2",
X"b03f8051",
X"f4be3f84",
X"39628738",
X"7a802efa",
X"84388055",
X"7483c080",
X"0c953d0d",
X"04fe3d0d",
X"83c7f051",
X"80f3ce3f",
X"f4e23f83",
X"c0800880",
X"2e863880",
X"51818b39",
X"f4e73f83",
X"c0800880",
X"ff38f587",
X"3f83c080",
X"08802eb9",
X"388151f2",
X"963f8051",
X"f49d3fef",
X"8a3f800b",
X"83c7d00c",
X"f9a43f83",
X"c0800853",
X"ff0b83c7",
X"d00cf0f6",
X"3f7280cc",
X"3883c7cc",
X"3351f3f7",
X"3f7251f1",
X"e63f80c1",
X"39f4af3f",
X"83c08008",
X"802eb638",
X"8151f1d3",
X"3f8051f3",
X"da3feec7",
X"3f8af80b",
X"83c0b80c",
X"83c7d408",
X"51ffb281",
X"3fff0b83",
X"c7d00cf0",
X"b13f83c7",
X"d4085280",
X"5185fd3f",
X"8151f5a0",
X"3f843d0d",
X"04fb3d0d",
X"805283c7",
X"f05180e2",
X"dc3f800b",
X"83c7cc34",
X"90808052",
X"86848080",
X"51c4d73f",
X"83c08008",
X"81933889",
X"be3f81dd",
X"e051c997",
X"3f83c080",
X"08559c80",
X"0a5480c0",
X"805381da",
X"a45283c0",
X"800851f6",
X"eb3f83c7",
X"e8085381",
X"dab45274",
X"51c3e13f",
X"83c08008",
X"8438f6f9",
X"3f83c7ec",
X"085381da",
X"c0527451",
X"c3ca3f83",
X"c08008b5",
X"38873dfc",
X"05548480",
X"805386a8",
X"80805283",
X"c7ec0851",
X"c1d63f83",
X"c0800893",
X"38758480",
X"802e0981",
X"06893881",
X"0b83c7cc",
X"34873980",
X"0b83c7cc",
X"3483c7cc",
X"3351f1fb",
X"3f8151f3",
X"e73f92fa",
X"3f8151f3",
X"df3f8151",
X"fd933ffa",
X"3983c08c",
X"080283c0",
X"8c0cfb3d",
X"0d0281da",
X"cc0b83c0",
X"b40c81da",
X"d00b83c0",
X"ac0c81da",
X"d40b83c0",
X"bc0c83c0",
X"8c08fc05",
X"0c800b83",
X"c7d40b83",
X"c08c08f8",
X"050c83c0",
X"8c08f405",
X"0cc1e73f",
X"83c08008",
X"8605fc06",
X"83c08c08",
X"f0050c02",
X"83c08c08",
X"f0050831",
X"0d833d70",
X"83c08c08",
X"f8050870",
X"840583c0",
X"8c08f805",
X"0c0c51ff",
X"beaf3f83",
X"c08c08f4",
X"05088105",
X"83c08c08",
X"f4050c83",
X"c08c08f4",
X"0508872e",
X"098106ff",
X"ac388694",
X"808051ea",
X"fb3fff0b",
X"83c7d00c",
X"800b83c8",
X"840c84d8",
X"c00b83c8",
X"800c8151",
X"eea53f81",
X"51eeca3f",
X"8051eec5",
X"3f8151ee",
X"eb3f8151",
X"efc03f82",
X"51ef8e3f",
X"8051efe4",
X"3f8051f0",
X"8e3f80d0",
X"e7528051",
X"ffbbe83f",
X"fcd73f83",
X"c08c08fc",
X"05080d80",
X"0b83c080",
X"0c873d0d",
X"83c08c0c",
X"04803d0d",
X"81ff5180",
X"0b83c890",
X"1234ff11",
X"5170f438",
X"823d0d04",
X"ff3d0d73",
X"70335351",
X"81113371",
X"34718112",
X"34833d0d",
X"04fb3d0d",
X"77795656",
X"80707155",
X"55527175",
X"25ac3872",
X"16703370",
X"147081ff",
X"06555151",
X"51717427",
X"89388112",
X"7081ff06",
X"53517181",
X"147083ff",
X"ff065552",
X"54747324",
X"d6387183",
X"c0800c87",
X"3d0d04fb",
X"3d0d7756",
X"ffb5943f",
X"83c08008",
X"802ef538",
X"83caac08",
X"86057081",
X"ff065253",
X"ffb3943f",
X"810b9088",
X"d4349088",
X"d4337081",
X"ff065153",
X"728638f9",
X"ec3fef39",
X"80557416",
X"75822b54",
X"549088c0",
X"13337434",
X"81155574",
X"852e0981",
X"06e83881",
X"0b9088d4",
X"34753383",
X"c8903481",
X"163383c8",
X"91348216",
X"3383c892",
X"34831633",
X"83c89334",
X"845283c8",
X"9051febd",
X"3f83c080",
X"0881ff06",
X"84173357",
X"5372762e",
X"0981068d",
X"38ffb3c0",
X"3f83c080",
X"08802e9a",
X"3883caac",
X"08a82e09",
X"81068938",
X"860b83ca",
X"ac0c8739",
X"a80b83ca",
X"ac0c80e4",
X"51eebe3f",
X"873d0d04",
X"f43d0d7e",
X"60595580",
X"5d807582",
X"2b7183ca",
X"b0120c83",
X"cac4175b",
X"5b577679",
X"3477772e",
X"83b83876",
X"527751ff",
X"bcf63f8e",
X"3dfc0554",
X"905383ca",
X"98527751",
X"ffbcb13f",
X"7c567590",
X"2e098106",
X"83943883",
X"ca9851fd",
X"973f83ca",
X"9a51fd90",
X"3f83ca9c",
X"51fd893f",
X"7683caa8",
X"0c7751ff",
X"b9fd3f81",
X"d8e05283",
X"c0800851",
X"ffa9a33f",
X"83c08008",
X"812e0981",
X"0680d438",
X"7683cac0",
X"0c820b83",
X"ca9834ff",
X"960b83ca",
X"99347751",
X"ffbcc23f",
X"83c08008",
X"5583c080",
X"08772588",
X"3883c080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"ca9a3474",
X"83ca9b34",
X"7683ca9c",
X"34ff800b",
X"83ca9d34",
X"81903983",
X"ca983383",
X"ca993371",
X"882b0756",
X"5b7483ff",
X"ff2e0981",
X"0680e838",
X"fe800b83",
X"cac00c81",
X"0b83caa8",
X"0cff0b83",
X"ca9834ff",
X"0b83ca99",
X"347751ff",
X"bbcf3f83",
X"c0800883",
X"cac80c83",
X"c0800855",
X"83c08008",
X"80258838",
X"83c08008",
X"8f055574",
X"842c7083",
X"ffff0670",
X"882a5851",
X"557583ca",
X"9a347483",
X"ca9b3476",
X"83ca9c34",
X"ff800b83",
X"ca9d3481",
X"0b83caa7",
X"34a53974",
X"85962e09",
X"810680fe",
X"387583ca",
X"c00c7751",
X"ffbb833f",
X"83caa733",
X"83c08008",
X"07557483",
X"caa73483",
X"caa73381",
X"06557480",
X"2e833884",
X"5783ca9c",
X"3383ca9d",
X"3371882b",
X"07565c74",
X"81802e09",
X"8106a138",
X"83ca9a33",
X"83ca9b33",
X"71882b07",
X"565bad80",
X"75278738",
X"76820757",
X"9c397681",
X"07579639",
X"7482802e",
X"09810687",
X"38768307",
X"57873974",
X"81ff268a",
X"387783ca",
X"b01b0c76",
X"79348e3d",
X"0d04803d",
X"0d728429",
X"83cab005",
X"700883c0",
X"800c5182",
X"3d0d04fe",
X"3d0d800b",
X"83ca940c",
X"800b83ca",
X"900cff0b",
X"83c88c0c",
X"a80b83ca",
X"ac0cae51",
X"ffade03f",
X"800b83ca",
X"b0545280",
X"73708405",
X"550c8112",
X"5271842e",
X"098106ef",
X"38843d0d",
X"04fe3d0d",
X"74028405",
X"96052253",
X"5371802e",
X"97387270",
X"81055433",
X"51ffadea",
X"3fff1270",
X"83ffff06",
X"5152e639",
X"843d0d04",
X"fe3d0d02",
X"92052253",
X"82ac51e9",
X"d03f80c3",
X"51ffadc6",
X"3f819651",
X"e9c33f72",
X"5283c890",
X"51ffb23f",
X"725283c8",
X"9051f8f1",
X"3f83c080",
X"0881ff06",
X"51ffada2",
X"3f843d0d",
X"04ffb13d",
X"0d80d13d",
X"f80551f9",
X"9a3f83ca",
X"94088105",
X"83ca940c",
X"80cf3d33",
X"cf117081",
X"ff065156",
X"56748326",
X"88ed3875",
X"8f06ff05",
X"567583c8",
X"8c082e9b",
X"38758326",
X"96387583",
X"c88c0c75",
X"842983ca",
X"b0057008",
X"53557551",
X"fa963f80",
X"762488c9",
X"38758429",
X"83cab005",
X"55740880",
X"2e88ba38",
X"83c88c08",
X"842983ca",
X"b0057008",
X"02880582",
X"b9053352",
X"5b557480",
X"d22e84b1",
X"387480d2",
X"24903874",
X"bf2e9c38",
X"7480d02e",
X"81d73887",
X"f8397480",
X"d32e80d2",
X"387480d7",
X"2e81c638",
X"87e73902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"5656ffac",
X"9e3f80c1",
X"51ffabd6",
X"3ff6ea3f",
X"860b83c8",
X"90348152",
X"83c89051",
X"ffacf93f",
X"8151fde4",
X"3f748938",
X"860b83ca",
X"ac0c8739",
X"a80b83ca",
X"ac0cffab",
X"ea3f80c1",
X"51ffaba2",
X"3ff6b63f",
X"900b83ca",
X"a7338106",
X"56567480",
X"2e833898",
X"5683ca9c",
X"3383ca9d",
X"3371882b",
X"07565974",
X"81802e09",
X"81069c38",
X"83ca9a33",
X"83ca9b33",
X"71882b07",
X"5657ad80",
X"75278c38",
X"75818007",
X"56853975",
X"a0075675",
X"83c89034",
X"ff0b83c8",
X"9134e00b",
X"83c89234",
X"800b83c8",
X"93348452",
X"83c89051",
X"ffabed3f",
X"8451869e",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055659",
X"ffaadc3f",
X"7951ffb5",
X"c93f83c0",
X"8008802e",
X"8b3880ce",
X"51ffaa86",
X"3f85f239",
X"80c151ff",
X"a9fc3fff",
X"aaf13fff",
X"a9a43f83",
X"cac00858",
X"8375259b",
X"3883ca9c",
X"3383ca9d",
X"3371882b",
X"07fc1771",
X"297a0583",
X"80055a51",
X"578d3974",
X"81802918",
X"ff800558",
X"81805780",
X"5676762e",
X"9338ffa9",
X"d53f83c0",
X"800883c8",
X"90173481",
X"1656ea39",
X"ffa9c33f",
X"83c08008",
X"81ff0677",
X"5383c890",
X"5256f4d9",
X"3f83c080",
X"0881ff06",
X"5575752e",
X"09810681",
X"8a38ffa9",
X"c23f80c1",
X"51ffa8fa",
X"3fffa9ef",
X"3f775279",
X"51ffb3d8",
X"3f805e80",
X"d13dfdf4",
X"05547653",
X"83c89052",
X"7951ffb1",
X"e53f0282",
X"b9053355",
X"81587480",
X"d72e0981",
X"06bd3880",
X"d13dfdf0",
X"05547653",
X"8f3d7053",
X"7a5259ff",
X"b2ea3f80",
X"5676762e",
X"a2387519",
X"83c89017",
X"33713370",
X"72327030",
X"70802570",
X"307e0681",
X"1d5d5e51",
X"5151525b",
X"55db3982",
X"ac51e489",
X"3f77802e",
X"863880c3",
X"51843980",
X"ce51ffa7",
X"f53fffa8",
X"ea3fffa7",
X"9d3f83dd",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055955",
X"80705d59",
X"ffa8903f",
X"80c151ff",
X"a7c83f83",
X"caa80879",
X"2e82de38",
X"83cac808",
X"80fc0555",
X"80fd5274",
X"5187b33f",
X"83c08008",
X"5b778224",
X"b238ff18",
X"70872b83",
X"ffff8006",
X"81dca005",
X"83c89059",
X"57558180",
X"55757081",
X"05573377",
X"70810559",
X"34ff1570",
X"81ff0651",
X"5574ea38",
X"828d3977",
X"82e82e81",
X"ab387782",
X"e92e0981",
X"0681b238",
X"81dad851",
X"ffadcb3f",
X"78587787",
X"32703070",
X"72078025",
X"7a8a3270",
X"30707207",
X"80257307",
X"53545a51",
X"57557580",
X"2e973878",
X"78269238",
X"a00b83c8",
X"901a3481",
X"197081ff",
X"065a55eb",
X"39811870",
X"81ff0659",
X"558a7827",
X"ffbc388f",
X"5883c88b",
X"183383c8",
X"901934ff",
X"187081ff",
X"06595577",
X"8426ea38",
X"9058800b",
X"83c89019",
X"34811870",
X"81ff0670",
X"982b5259",
X"55748025",
X"e93880c6",
X"557a858f",
X"24843880",
X"c2557483",
X"c8903480",
X"f10b83c8",
X"9334810b",
X"83c89434",
X"7a83c891",
X"347a882c",
X"557483c8",
X"923480cb",
X"3982f078",
X"2580c438",
X"7780fd29",
X"fd97d305",
X"527951ff",
X"b0863f80",
X"d13dfdec",
X"055480fd",
X"5383c890",
X"527951ff",
X"afbe3f7b",
X"81195956",
X"7580fc24",
X"83387858",
X"77882c55",
X"7483c98d",
X"347783c9",
X"8e347583",
X"c98f3481",
X"805980cc",
X"3983cac0",
X"08578378",
X"259b3883",
X"ca9c3383",
X"ca9d3371",
X"882b07fc",
X"1a712979",
X"05838005",
X"5951598d",
X"39778180",
X"2917ff80",
X"05578180",
X"59765279",
X"51ffaf94",
X"3f80d13d",
X"fdec0554",
X"785383c8",
X"90527951",
X"ffaecd3f",
X"7851f6b8",
X"3fffa587",
X"3fffa3ba",
X"3f8b3983",
X"ca900881",
X"0583ca90",
X"0c80d13d",
X"0d04f6d9",
X"3ffc39fc",
X"3d0d7678",
X"71842983",
X"cab00570",
X"08515353",
X"53709e38",
X"80ce7234",
X"80cf0b81",
X"133480ce",
X"0b821334",
X"80c50b83",
X"13347084",
X"133480e7",
X"3983cac4",
X"13335480",
X"d2723473",
X"822a7081",
X"06515180",
X"cf537084",
X"3880d753",
X"72811334",
X"a00b8213",
X"34738306",
X"5170812e",
X"9e387081",
X"24883870",
X"802e8f38",
X"9f397082",
X"2e923870",
X"832e9238",
X"933980d8",
X"558e3980",
X"d3558939",
X"80cd5584",
X"3980c455",
X"74831334",
X"80c40b84",
X"1334800b",
X"85133486",
X"3d0d04fc",
X"3d0d7655",
X"80750c80",
X"0b84160c",
X"800b8816",
X"0c800b8c",
X"160c83c7",
X"f05180dc",
X"bc3f87a6",
X"80337081",
X"ff065152",
X"de9a3f71",
X"812a8132",
X"72813271",
X"81067181",
X"06318418",
X"0c545471",
X"832a8132",
X"72822a81",
X"32718106",
X"71810631",
X"770c5353",
X"87a09033",
X"70098106",
X"88170c52",
X"83c08008",
X"802e80c2",
X"3883c080",
X"08812a70",
X"810683c0",
X"80088106",
X"3184170c",
X"5283c080",
X"08832a83",
X"c0800882",
X"2a718106",
X"71810631",
X"770c5353",
X"83c08008",
X"842a8106",
X"88160c83",
X"c0800885",
X"2a81068c",
X"160c863d",
X"0d04fe3d",
X"0d747654",
X"527151fe",
X"c63f7281",
X"2ea23881",
X"73268d38",
X"72822ea8",
X"3872832e",
X"9c38e639",
X"7108e238",
X"841208dd",
X"38881208",
X"d838a539",
X"88120881",
X"2e9e3891",
X"39881208",
X"812e9538",
X"71089138",
X"8412088c",
X"388c1208",
X"812e0981",
X"06ffb238",
X"843d0d04",
X"fc3d0d76",
X"78535481",
X"53805587",
X"39711073",
X"10545273",
X"72265172",
X"802ea738",
X"70802e86",
X"38718025",
X"e8387280",
X"2e983871",
X"74268938",
X"73723175",
X"74075654",
X"72812a72",
X"812a5353",
X"e5397351",
X"78833874",
X"517083c0",
X"800c863d",
X"0d04fe3d",
X"0d805375",
X"527451ff",
X"a33f843d",
X"0d04fe3d",
X"0d815375",
X"527451ff",
X"933f843d",
X"0d04fb3d",
X"0d777955",
X"55805674",
X"76258638",
X"74305581",
X"56738025",
X"88387330",
X"76813257",
X"54805373",
X"527451fe",
X"e73f83c0",
X"80085475",
X"802e8738",
X"83c08008",
X"30547383",
X"c0800c87",
X"3d0d04fa",
X"3d0d787a",
X"57558057",
X"74772586",
X"38743055",
X"8157759f",
X"2c548153",
X"75743274",
X"31527451",
X"feaa3f83",
X"c0800854",
X"76802e87",
X"3883c080",
X"08305473",
X"83c0800c",
X"883d0d04",
X"fb3d0d78",
X"0284059f",
X"05335556",
X"800b81d6",
X"e8565381",
X"732b7406",
X"5271802e",
X"83388152",
X"74708205",
X"56227073",
X"902b0790",
X"809c0c51",
X"81135372",
X"882e0981",
X"06d93880",
X"5383cad0",
X"13335170",
X"81ff2eb2",
X"38701081",
X"d5880570",
X"22555180",
X"73177033",
X"701081d5",
X"88057022",
X"51515152",
X"5273712e",
X"91388112",
X"5271862e",
X"098106f1",
X"38739080",
X"9c0c8113",
X"5372862e",
X"098106ff",
X"b8388053",
X"72167033",
X"51517081",
X"ff2e9438",
X"701081d5",
X"88057022",
X"70848080",
X"0790809c",
X"0c515181",
X"13537286",
X"2e098106",
X"d7388053",
X"72165170",
X"3383cad0",
X"14348113",
X"5372862e",
X"098106ec",
X"38873d0d",
X"0404ff3d",
X"0d740284",
X"058f0533",
X"52527088",
X"38719080",
X"940c8e39",
X"70812e09",
X"81068638",
X"71908098",
X"0c833d0d",
X"04fb3d0d",
X"029f0533",
X"79982b70",
X"982c7c98",
X"2b70982c",
X"83caec15",
X"70337098",
X"2b70982c",
X"51585c5a",
X"51555154",
X"5470732e",
X"09810694",
X"3883cacc",
X"14337098",
X"2b70982c",
X"51525670",
X"722eb138",
X"72753471",
X"83cacc15",
X"3483cacd",
X"3383caed",
X"3371982b",
X"71902b07",
X"83cacc33",
X"70882b72",
X"0783caec",
X"33710790",
X"80b80c52",
X"59535452",
X"873d0d04",
X"fe3d0d74",
X"81113371",
X"3371882b",
X"0783c080",
X"0c535184",
X"3d0d0483",
X"cad83383",
X"c0800c04",
X"f53d0d02",
X"bb053302",
X"8405bf05",
X"33028805",
X"80c30533",
X"028c0580",
X"c6052266",
X"5c5a5e5c",
X"567a557b",
X"548953a1",
X"527d5180",
X"d0c03f83",
X"c0800881",
X"ff0683c0",
X"800c8d3d",
X"0d0483c0",
X"8c080283",
X"c08c0cf5",
X"3d0d83c0",
X"8c088805",
X"0883c08c",
X"088f0533",
X"83c08c08",
X"92052202",
X"8c057390",
X"0583c08c",
X"08e8050c",
X"83c08c08",
X"f8050c83",
X"c08c08f0",
X"050c83c0",
X"8c08ec05",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08f005",
X"0883c08c",
X"08e0050c",
X"83c08c08",
X"fc050c83",
X"c08c08f0",
X"05088927",
X"8a38890b",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"05088605",
X"87fffc06",
X"83c08c08",
X"e0050c02",
X"83c08c08",
X"e0050831",
X"0d853d70",
X"5583c08c",
X"08ec0508",
X"5483c08c",
X"08f00508",
X"5383c08c",
X"08f40508",
X"5283c08c",
X"08e4050c",
X"80d9f23f",
X"83c08008",
X"81ff0683",
X"c08c08e4",
X"050883c0",
X"8c08ec05",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"e0050880",
X"2e8c3883",
X"c08c08f8",
X"05080d89",
X"c83983c0",
X"8c08f005",
X"08802e89",
X"a63883c0",
X"8c08ec05",
X"08810533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508842e",
X"a938840b",
X"83c08c08",
X"e0050825",
X"88c73883",
X"c08c08e0",
X"0508852e",
X"859b3883",
X"c08c08e0",
X"0508a12e",
X"87ad3888",
X"ac39800b",
X"83c08c08",
X"ec050885",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08fc050c",
X"83c08c08",
X"e0050883",
X"2e098106",
X"88833883",
X"c08c08e8",
X"05088105",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e0050881",
X"2687e638",
X"810b83c0",
X"8c08e005",
X"0880d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08fc",
X"050c83c0",
X"8c08ec05",
X"08820533",
X"83c08c08",
X"e0050887",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088b",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"e005088c",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088d",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"e005088e",
X"052383c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088a",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"70940508",
X"fcffff06",
X"7194050c",
X"83c08c08",
X"e0050c83",
X"c08c08ec",
X"05088605",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"f4050c83",
X"c08c08e0",
X"050883c0",
X"8c08fc05",
X"082e0981",
X"06b63883",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c83",
X"c08c08fc",
X"050883c0",
X"8c08e005",
X"088b0534",
X"83c08c08",
X"ec050887",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"812e8f38",
X"83c08c08",
X"e0050882",
X"2eb73884",
X"8c3983c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c820b",
X"83c08c08",
X"e005088a",
X"053483d9",
X"3983c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08fc0508",
X"83c08c08",
X"e005088a",
X"053483a1",
X"3983c08c",
X"08fc0508",
X"802e8395",
X"3883c08c",
X"08ec0508",
X"83053383",
X"0683c08c",
X"08e0050c",
X"83c08c08",
X"e0050883",
X"2e098106",
X"82f33883",
X"c08c08ec",
X"05088205",
X"3370982b",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c83c0",
X"8c08e005",
X"08802582",
X"cc3883c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c83c0",
X"8c08ec05",
X"08860533",
X"83c08c08",
X"e0050880",
X"d6053483",
X"c08c08e0",
X"05088405",
X"83c08c08",
X"ec050882",
X"05338f06",
X"83c08c08",
X"e4050c83",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0883c08c",
X"08e00508",
X"3483c08c",
X"08ec0508",
X"84053383",
X"c08c08e0",
X"05088105",
X"34800b83",
X"c08c08e0",
X"05088205",
X"3483c08c",
X"08e00508",
X"08ff83ff",
X"06828007",
X"83c08c08",
X"e005080c",
X"83c08c08",
X"e8050881",
X"05338105",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"050883c0",
X"8c08e805",
X"08810534",
X"81833983",
X"c08c08fc",
X"0508802e",
X"80f73883",
X"c08c08ec",
X"05088605",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e00508a2",
X"2e098106",
X"80d73883",
X"c08c08ec",
X"05088805",
X"3383c08c",
X"08ec0508",
X"87053371",
X"82802905",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c5283c0",
X"8c08e405",
X"0c83c08c",
X"08f4050c",
X"83c08c08",
X"e4050883",
X"c08c08e0",
X"05088805",
X"2383c08c",
X"08ec0508",
X"3383c08c",
X"08f00508",
X"71317083",
X"ffff0683",
X"c08c08f0",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08ec0508",
X"0583c08c",
X"08ec050c",
X"f6d03983",
X"c08c08f8",
X"05080d83",
X"c08c08f0",
X"050883c0",
X"8c08e005",
X"0c83c08c",
X"08f80508",
X"0d83c08c",
X"08e00508",
X"83c0800c",
X"8d3d0d83",
X"c08c0c04",
X"83c08c08",
X"0283c08c",
X"0ce63d0d",
X"83c08c08",
X"88050802",
X"840583c0",
X"8c08e805",
X"0c83c08c",
X"08d4050c",
X"800b83ca",
X"f43483c0",
X"8c08d405",
X"08900583",
X"c08c08c0",
X"050c800b",
X"83c08c08",
X"c0050834",
X"800b83c0",
X"8c08c005",
X"08810534",
X"800b83c0",
X"8c08c405",
X"0c83c08c",
X"08c40508",
X"80d82983",
X"c08c08c0",
X"05080583",
X"c08c08ff",
X"b4050c80",
X"0b83c08c",
X"08ffb405",
X"0880d805",
X"0c83c08c",
X"08ffb405",
X"08840583",
X"c08c08ff",
X"b4050c83",
X"c08c08c4",
X"050883c0",
X"8c08ffb4",
X"05083488",
X"0b83c08c",
X"08ffb405",
X"08810534",
X"800b83c0",
X"8c08ffb4",
X"05088205",
X"3483c08c",
X"08ffb405",
X"0808ffa1",
X"ff06a080",
X"0783c08c",
X"08ffb405",
X"080c83c0",
X"8c08c405",
X"08810570",
X"81ff0683",
X"c08c08c4",
X"050c83c0",
X"8c08ffb4",
X"050c810b",
X"83c08c08",
X"c4050827",
X"fedb3883",
X"c08c08ec",
X"05705483",
X"c08c08c8",
X"050c9252",
X"83c08c08",
X"d4050851",
X"80cd993f",
X"83c08008",
X"81ff0670",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"8dea3883",
X"c08c08f4",
X"0551f18c",
X"3f83c080",
X"0883ffff",
X"0683c08c",
X"08f60552",
X"83c08c08",
X"e4050cf0",
X"f33f83c0",
X"800883ff",
X"ff0683c0",
X"8c08fd05",
X"3383c08c",
X"08ffb805",
X"0883c08c",
X"08c4050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"e0050c83",
X"c08c08c4",
X"050883c0",
X"8c08ffbc",
X"05082780",
X"fe3883c0",
X"8c08c805",
X"085483c0",
X"8c08c405",
X"08538952",
X"83c08c08",
X"d4050851",
X"80cc9e3f",
X"83c08008",
X"81ff0683",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b8050880",
X"f23883c0",
X"8c08ee05",
X"51eff13f",
X"83c08008",
X"83ffff06",
X"5383c08c",
X"08c40508",
X"5283c08c",
X"08d40508",
X"51f0b33f",
X"83c08c08",
X"c4050881",
X"057081ff",
X"0683c08c",
X"08c4050c",
X"83c08c08",
X"ffb4050c",
X"fef13983",
X"c08c08c0",
X"05088105",
X"3383c08c",
X"08ffb405",
X"0c81db0b",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb40508",
X"802e8be0",
X"38943983",
X"c08c08ff",
X"b8050883",
X"c08c08ff",
X"bc050c8b",
X"cb3983c0",
X"8c08f105",
X"335283c0",
X"8c08d405",
X"085180cb",
X"9c3f800b",
X"83c08c08",
X"c0050881",
X"053383c0",
X"8c08ffb4",
X"050c83c0",
X"8c08c405",
X"0c83c08c",
X"08c40508",
X"83c08c08",
X"ffb40508",
X"2789e638",
X"83c08c08",
X"c4050880",
X"d8297083",
X"c08c08c0",
X"05080570",
X"88057083",
X"053383c0",
X"8c08cc05",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"d8050c83",
X"c08c08cc",
X"050887a6",
X"3883c08c",
X"08c80508",
X"22028405",
X"71860587",
X"fffc0683",
X"c08c08ff",
X"b4050c83",
X"c08c08dc",
X"050c83c0",
X"8c08ffb8",
X"050c0283",
X"c08c08ff",
X"b4050831",
X"0d893d70",
X"5983c08c",
X"08ffb805",
X"085883c0",
X"8c08ffbc",
X"05088705",
X"335783c0",
X"8c08ffb4",
X"050ca255",
X"83c08c08",
X"cc050854",
X"86538181",
X"5283c08c",
X"08d40508",
X"51be933f",
X"83c08008",
X"81ff0683",
X"c08c08d0",
X"050c83c0",
X"8c08d005",
X"0881c138",
X"83c08c08",
X"ffbc0508",
X"96055383",
X"c08c08ff",
X"b8050852",
X"83c08c08",
X"ffb40508",
X"51a1c63f",
X"83c08008",
X"81ff0683",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b4050880",
X"2e818538",
X"83c08c08",
X"ffbc0508",
X"940583c0",
X"8c08ffbc",
X"05089605",
X"3370862a",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"cc050c83",
X"c08c08ff",
X"b4050883",
X"2e098106",
X"80c63883",
X"c08c08ff",
X"b4050883",
X"c08c08c8",
X"05088205",
X"3483cad8",
X"33708105",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb40508",
X"83cad834",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"cc050834",
X"83c08c08",
X"dc05080d",
X"83c08c08",
X"d0050881",
X"ff0683c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"0508fbff",
X"3883c08c",
X"08d80508",
X"83c08c08",
X"c0050805",
X"88057082",
X"05335183",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b4050883",
X"2e098106",
X"80e33883",
X"c08c08ff",
X"b8050883",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b4050881",
X"057081ff",
X"065183c0",
X"8c08ffb4",
X"050c810b",
X"83c08c08",
X"ffb40508",
X"27dd3880",
X"0b83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb405",
X"08810570",
X"81ff0651",
X"83c08c08",
X"ffb4050c",
X"970b83c0",
X"8c08ffb4",
X"050827dd",
X"3883c08c",
X"08e40508",
X"80f93270",
X"30708025",
X"515183c0",
X"8c08ffb4",
X"050c83c0",
X"8c08e005",
X"08912e09",
X"810680f9",
X"3883c08c",
X"08ffb405",
X"08802e80",
X"ec3883c0",
X"8c08c405",
X"0880e238",
X"850b83c0",
X"8c08c005",
X"08a60534",
X"a00b83c0",
X"8c08c005",
X"08a70534",
X"850b83c0",
X"8c08c005",
X"08a80534",
X"80c00b83",
X"c08c08c0",
X"0508a905",
X"34860b83",
X"c08c08c0",
X"0508aa05",
X"34900b83",
X"c08c08c0",
X"0508ab05",
X"34860b83",
X"c08c08c0",
X"0508ac05",
X"34a00b83",
X"c08c08c0",
X"0508ad05",
X"3483c08c",
X"08e40508",
X"89d83270",
X"30708025",
X"515183c0",
X"8c08ffb4",
X"050c83c0",
X"8c08e005",
X"0883edec",
X"2e098106",
X"80f63881",
X"7083c08c",
X"08ffb405",
X"080683c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb4",
X"0508802e",
X"80ce3883",
X"c08c08c4",
X"050880c4",
X"38840b83",
X"c08c08c0",
X"0508aa05",
X"3480c00b",
X"83c08c08",
X"c00508ab",
X"0534840b",
X"83c08c08",
X"c00508ac",
X"0534900b",
X"83c08c08",
X"c00508ad",
X"053483c0",
X"8c08ffb8",
X"050883c0",
X"8c08c005",
X"088c0534",
X"83c08c08",
X"e4050880",
X"f9327030",
X"70802551",
X"5183c08c",
X"08ffb405",
X"0c83c08c",
X"08e00508",
X"862e0981",
X"0680c338",
X"817083c0",
X"8c08ffb4",
X"05080683",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b4050880",
X"2e9c3883",
X"c08c08c4",
X"05089338",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"c005088d",
X"053483c0",
X"8c08c405",
X"0880d829",
X"83c08c08",
X"c0050805",
X"70840570",
X"83053383",
X"c08c08ff",
X"b4050c83",
X"c08c08c8",
X"050c83c0",
X"8c08ffbc",
X"050c8058",
X"805783c0",
X"8c08ffb4",
X"05085680",
X"5580548a",
X"53a15283",
X"c08c08d4",
X"050851b7",
X"8d3f83c0",
X"800881ff",
X"06703070",
X"9f2a5183",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b80508a0",
X"2e8c3883",
X"c08c08ff",
X"b40508f6",
X"c23883c0",
X"8c08ffbc",
X"05088b05",
X"3383c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb405",
X"08802eb3",
X"3883c08c",
X"08c80508",
X"83053383",
X"c08c08ff",
X"b4050c80",
X"58805783",
X"c08c08ff",
X"b4050856",
X"80558054",
X"8b53a152",
X"83c08c08",
X"d4050851",
X"b6883f83",
X"c08c08c4",
X"05088105",
X"7081ff06",
X"83c08c08",
X"c0050881",
X"05335283",
X"c08c08c4",
X"050c83c0",
X"8c08ffb4",
X"050cf689",
X"39800b83",
X"c08c08c4",
X"050c83c0",
X"8c08c405",
X"0880d829",
X"83c08c08",
X"d4050805",
X"709a0533",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb40508",
X"822e0981",
X"06a93883",
X"caf45681",
X"55805483",
X"c08c08ff",
X"b4050853",
X"83c08c08",
X"ffb80508",
X"97053352",
X"83c08c08",
X"d4050851",
X"e48a3f83",
X"c08c08c4",
X"05088105",
X"7081ff06",
X"83c08c08",
X"c4050c83",
X"c08c08ff",
X"b4050c81",
X"0b83c08c",
X"08c40508",
X"27fefb38",
X"810b83c0",
X"8c08c005",
X"0834800b",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"e805080d",
X"83c08c08",
X"ffbc0508",
X"83c0800c",
X"9c3d0d83",
X"c08c0c04",
X"f53d0d90",
X"1e57800b",
X"81183354",
X"59787327",
X"819d3878",
X"80d82917",
X"8a113354",
X"5472832e",
X"09810680",
X"f8389414",
X"335ba98c",
X"3f83c080",
X"085a8056",
X"7581c429",
X"1a871133",
X"54547280",
X"2e80c038",
X"730881d4",
X"fc2e0981",
X"06b53880",
X"74595574",
X"80d82918",
X"9a113354",
X"5472832e",
X"09810692",
X"38a41470",
X"3354547a",
X"73278738",
X"ff135372",
X"74348115",
X"7081ff06",
X"56538175",
X"27d13881",
X"167081ff",
X"0657538f",
X"7627ffa4",
X"3883cad8",
X"33ff0553",
X"7283cad8",
X"34811970",
X"81ff0681",
X"19335e5a",
X"537b7926",
X"fee53880",
X"0b83c080",
X"0c8d3d0d",
X"0483c08c",
X"080283c0",
X"8c0ce63d",
X"0d83c08c",
X"08880508",
X"02840571",
X"90057033",
X"7083c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"dc050c83",
X"c08c08e0",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"94b53880",
X"0b83c08c",
X"08c80508",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08d4",
X"050c83c0",
X"8c08d405",
X"0883c08c",
X"08ffa405",
X"082593fd",
X"3883c08c",
X"08d40508",
X"80d82983",
X"c08c08c8",
X"05080584",
X"05708605",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffa405",
X"08802e93",
X"8938a6b2",
X"3f83c08c",
X"08ffb805",
X"0880d405",
X"0883c080",
X"082692f2",
X"380283c0",
X"8c08ffb8",
X"05088105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08d8050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"fc052383",
X"c08c08ff",
X"a4050886",
X"0583fc06",
X"83c08c08",
X"ffa4050c",
X"0283c08c",
X"08ffa405",
X"08310d85",
X"3d705583",
X"c08c08fc",
X"055483c0",
X"8c08ffb8",
X"05085383",
X"c08c08e0",
X"05085283",
X"c08c08c0",
X"050cae8a",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"91bb3883",
X"c08c08ff",
X"b8050887",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"80d53883",
X"c08c08ff",
X"b8050886",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508822e",
X"098106b3",
X"3883c08c",
X"08fc0522",
X"83c08c08",
X"ffa4050c",
X"870b83c0",
X"8c08ffa4",
X"05082797",
X"3883c08c",
X"08c00508",
X"82055283",
X"c08c08c0",
X"05083351",
X"dba63f83",
X"c08c08ff",
X"b8050886",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508832e",
X"09810690",
X"a43883c0",
X"8c08ffb8",
X"05089205",
X"70820533",
X"83c08c08",
X"fc052283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08c4",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffa8",
X"0508268f",
X"e438800b",
X"83c08c08",
X"e4050c80",
X"0b83c08c",
X"08ffb005",
X"0c83c08c",
X"08ffb005",
X"081083c0",
X"8c0805f8",
X"0583c08c",
X"08ffb005",
X"08842983",
X"c08c08ff",
X"b0050810",
X"0583c08c",
X"08c40508",
X"05708405",
X"703383c0",
X"8c08c005",
X"08057033",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffbc0508",
X"2383c08c",
X"08ffa805",
X"08810533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"902e0981",
X"06be3883",
X"c08c08ff",
X"a8050833",
X"83c08c08",
X"c0050805",
X"81057033",
X"70828029",
X"83c08c08",
X"ffb40508",
X"05515183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"bc050823",
X"83c08c08",
X"ffac0508",
X"86052283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a80508a2",
X"3883c08c",
X"08ffac05",
X"08880522",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"81ff2e80",
X"e53883c0",
X"8c08ffbc",
X"05082270",
X"83c08c08",
X"ffa80508",
X"31708280",
X"29713183",
X"c08c08ff",
X"ac050888",
X"05227083",
X"c08c08ff",
X"a8050831",
X"70733553",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffbc05",
X"082383c0",
X"8c08ffb0",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa4050c",
X"810b83c0",
X"8c08ffb0",
X"050827fc",
X"e03883c0",
X"8c08f805",
X"2283c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08bf2691",
X"3883c08c",
X"08e40508",
X"820783c0",
X"8c08e405",
X"0c81c00b",
X"83c08c08",
X"ffa40508",
X"27913883",
X"c08c08e4",
X"05088107",
X"83c08c08",
X"e4050c83",
X"c08c08fa",
X"052283c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508bf26",
X"913883c0",
X"8c08e405",
X"08880783",
X"c08c08e4",
X"050c81c0",
X"0b83c08c",
X"08ffa405",
X"08279138",
X"83c08c08",
X"e4050884",
X"0783c08c",
X"08e4050c",
X"800b83c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffb0",
X"05081083",
X"c08c08c4",
X"05080570",
X"90057033",
X"83c08c08",
X"c0050805",
X"70337281",
X"05337072",
X"06515351",
X"83c08c08",
X"ffa8050c",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e9b",
X"38900b83",
X"c08c08ff",
X"b005082b",
X"83c08c08",
X"e4050807",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"b0050881",
X"057081ff",
X"0683c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa405",
X"0c970b83",
X"c08c08ff",
X"b0050827",
X"fef43883",
X"c08c08ff",
X"b8050890",
X"053383c0",
X"8c08e405",
X"0883c08c",
X"08ffb405",
X"0c83c08c",
X"08c4050c",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffb80508",
X"8c05082e",
X"83ff3883",
X"c08c08ff",
X"b4050883",
X"c08c08ff",
X"b805088c",
X"050c83c0",
X"8c08ffb8",
X"05088905",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e83",
X"b93883c0",
X"8c08e405",
X"83c08c08",
X"ffb40508",
X"8f0683c0",
X"8c08e405",
X"0c83c08c",
X"08cc050c",
X"800b83c0",
X"8c08f005",
X"0c800b83",
X"c08c08f4",
X"0523800b",
X"81d6f833",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffbc0508",
X"2e82d338",
X"83c08c08",
X"f00581d6",
X"f80b83c0",
X"8c08ffac",
X"050c83c0",
X"8c08d005",
X"0c83c08c",
X"08ffac05",
X"083383c0",
X"8c08ffac",
X"05088105",
X"3381722b",
X"81722b07",
X"7083c08c",
X"08ffb405",
X"08065283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"a805082e",
X"09810681",
X"be3883c0",
X"8c08ffbc",
X"05088526",
X"80f63883",
X"c08c08ff",
X"ac050882",
X"05337081",
X"ff0683c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"80ca3883",
X"c08c08ff",
X"bc050883",
X"c08c08ff",
X"bc050881",
X"057081ff",
X"0683c08c",
X"08d00508",
X"73055383",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b0050883",
X"c08c08ff",
X"a4050834",
X"83c08c08",
X"ffac0508",
X"83053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e9d3881",
X"0b83c08c",
X"08ffa405",
X"082b83c0",
X"8c08cc05",
X"08080783",
X"c08c08cc",
X"05080c83",
X"c08c08ff",
X"ac050884",
X"05703383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a40508fd",
X"c83883c0",
X"8c08f005",
X"528051d0",
X"c33f83c0",
X"8c08e405",
X"085283c0",
X"8c08c405",
X"0851d1fe",
X"3f83c08c",
X"08fb0533",
X"7081800a",
X"29810a05",
X"70982c55",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"f9053370",
X"81800a29",
X"810a0570",
X"982c5583",
X"c08c08ff",
X"a4050c83",
X"c08c08c4",
X"05085383",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a8050cd1",
X"d43f83c0",
X"8c08ffb8",
X"05088805",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e84",
X"e03883c0",
X"8c08ffb8",
X"05089005",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08812684",
X"c0388070",
X"81d7ac0b",
X"81d7ac0b",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"b405082e",
X"81ae3883",
X"c08c08ff",
X"ac050884",
X"2983c08c",
X"08ffa805",
X"08057033",
X"83c08c08",
X"c0050805",
X"70337281",
X"05337072",
X"06515351",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802eaa38",
X"810b83c0",
X"8c08ffac",
X"05082b83",
X"c08c08ff",
X"b4050807",
X"7083ffff",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffac05",
X"08810570",
X"81ff0681",
X"d7ac7184",
X"29710570",
X"81053351",
X"5383c08c",
X"08ffa805",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08fed438",
X"83c08c08",
X"ffb80508",
X"8a052283",
X"c08c08c0",
X"050c83c0",
X"8c08ffb4",
X"050883c0",
X"8c08c005",
X"082e82ad",
X"38800b83",
X"c08c08e8",
X"050c800b",
X"83c08c08",
X"ec052380",
X"7083c08c",
X"08e80583",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"b0050c81",
X"af3983c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffac",
X"05082c70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e80e738",
X"83c08c08",
X"ffb00508",
X"83c08c08",
X"ffb00508",
X"81057081",
X"ff0683c0",
X"8c08ffbc",
X"05087305",
X"83c08c08",
X"ffb80508",
X"90053383",
X"c08c08ff",
X"ac050884",
X"29055353",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa80508",
X"81d7ae05",
X"3383c08c",
X"08ffa405",
X"083483c0",
X"8c08ffac",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa4050c",
X"8f0b83c0",
X"8c08ffac",
X"05082783",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b0050885",
X"268c3883",
X"c08c08ff",
X"a40508fe",
X"a93883c0",
X"8c08e805",
X"528051ca",
X"f33f83c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffb8",
X"05088a05",
X"2383c08c",
X"08ffb805",
X"0880d205",
X"3383c08c",
X"08ffb805",
X"0880d405",
X"080583c0",
X"8c08ffb8",
X"050880d4",
X"050c83c0",
X"8c08d805",
X"080d83c0",
X"8c08d405",
X"0881800a",
X"2981800a",
X"0570982c",
X"83c08c08",
X"c8050881",
X"053383c0",
X"8c08ffa8",
X"050c5183",
X"c08c08d4",
X"050c83c0",
X"8c08ffa8",
X"050883c0",
X"8c08d405",
X"0824ec85",
X"38800b83",
X"c08c08ff",
X"a8050c83",
X"c08c08dc",
X"05080d83",
X"c08c08ff",
X"a8050883",
X"c0800c9c",
X"3d0d83c0",
X"8c0c04f3",
X"3d0d02bf",
X"05330284",
X"0580c305",
X"3383caf4",
X"335a5b59",
X"79802e8d",
X"38787806",
X"5776802e",
X"8e388189",
X"39787806",
X"5776802e",
X"80ff3883",
X"caf43370",
X"7a075858",
X"79883878",
X"09707906",
X"51577683",
X"caf43492",
X"973f83c0",
X"80085e80",
X"5c8f5d7d",
X"1c871133",
X"58587680",
X"2e80c138",
X"770881d4",
X"fc2e0981",
X"06b63880",
X"5b815a7d",
X"1c701c9a",
X"11335959",
X"5976822e",
X"09810694",
X"3883caf4",
X"56815580",
X"54765397",
X"18335278",
X"51cbc53f",
X"ff1a80d8",
X"1c5c5a79",
X"8025d038",
X"ff1d81c4",
X"1d5d5d7c",
X"8025ffa7",
X"388f3d0d",
X"04e93d0d",
X"696c0288",
X"0580ea05",
X"225c5a5b",
X"80707141",
X"5e58ff78",
X"797a7b7c",
X"7d464c4a",
X"45405d43",
X"62993d34",
X"62028405",
X"80dd0534",
X"77792280",
X"ffff0654",
X"45727923",
X"79782e88",
X"87387a70",
X"81055c33",
X"70842a71",
X"8c067082",
X"2a5a5656",
X"8306ff1b",
X"7083ffff",
X"065c5456",
X"80547574",
X"2e91387a",
X"7081055c",
X"33ff1b70",
X"83ffff06",
X"5c545481",
X"76279b38",
X"7381ff06",
X"7b708105",
X"5d335574",
X"82802905",
X"ff1b7083",
X"ffff065c",
X"54548276",
X"27aa3873",
X"83ffff06",
X"7b708105",
X"5d337090",
X"2b72077d",
X"7081055f",
X"3370982b",
X"7207fe1f",
X"7083ffff",
X"06405252",
X"52525454",
X"7e802e80",
X"c4387686",
X"f738748a",
X"2e098106",
X"9438811f",
X"7081ff06",
X"811e7081",
X"ff065f52",
X"405386dc",
X"39748c2e",
X"09810686",
X"d338ff1f",
X"7081ff06",
X"ff1e7081",
X"ff065f52",
X"40537b63",
X"2586bd38",
X"ff4386b8",
X"3976812e",
X"83bb3876",
X"81248938",
X"76802e8d",
X"3886a539",
X"76822e84",
X"a638869c",
X"39f81553",
X"72842684",
X"95387284",
X"2981d7ec",
X"05537208",
X"0464802e",
X"80cd3878",
X"22838080",
X"06537283",
X"80802e09",
X"8106bc38",
X"80567564",
X"27a43875",
X"1e7083ff",
X"ff067710",
X"1b901172",
X"832a5851",
X"57515373",
X"75347287",
X"0681712b",
X"51537281",
X"16348116",
X"7081ff06",
X"57539776",
X"27cc387f",
X"84074080",
X"0b993d43",
X"56611670",
X"3370982b",
X"70982c51",
X"51515380",
X"732480fb",
X"38607329",
X"1e7083ff",
X"ff067a22",
X"83808006",
X"52585372",
X"8380802e",
X"09810680",
X"de386088",
X"32703070",
X"72078025",
X"63903270",
X"30707207",
X"80257307",
X"53545851",
X"55537380",
X"2ebd3876",
X"87065372",
X"b6387584",
X"29761005",
X"79118411",
X"79832a57",
X"57515373",
X"75346081",
X"16346586",
X"14236688",
X"14237587",
X"387f8107",
X"408d3975",
X"812e0981",
X"0685387f",
X"82074081",
X"167081ff",
X"06575381",
X"7627fee5",
X"38636129",
X"1e7083ff",
X"ff065f53",
X"80704642",
X"ff028405",
X"80dd0534",
X"ff0b993d",
X"3483f539",
X"811c7081",
X"ff065d53",
X"80427381",
X"2e098106",
X"8e387781",
X"800a2981",
X"800a0558",
X"80d33973",
X"802e8938",
X"73822e09",
X"81068d38",
X"7c81800a",
X"2981800a",
X"055da439",
X"815f83b8",
X"39ff1c70",
X"81ff065d",
X"537b6325",
X"8338ff43",
X"7c802e92",
X"387c8180",
X"0a2981ff",
X"0a055d7c",
X"982c5d83",
X"93397780",
X"2e923877",
X"81800a29",
X"81ff0a05",
X"5877982c",
X"5882fd39",
X"7753839e",
X"39748926",
X"80f43874",
X"842981d8",
X"80055372",
X"08047387",
X"2e82e138",
X"73852e82",
X"db387388",
X"2e82d538",
X"738c2e82",
X"cf387389",
X"2e098106",
X"86388145",
X"82c23973",
X"812e0981",
X"0682b938",
X"62802582",
X"b3387b98",
X"2b70982c",
X"514382a8",
X"397383ff",
X"ff064682",
X"9f397383",
X"ffff0647",
X"82963973",
X"81ff0641",
X"828e3973",
X"811a3482",
X"87397381",
X"ff064481",
X"ff397e53",
X"82a03974",
X"812e81e3",
X"38748124",
X"89387480",
X"2e8d3881",
X"e7397482",
X"2e81d838",
X"81de3974",
X"567b8338",
X"81567453",
X"73862e09",
X"81069738",
X"75810653",
X"72802e8e",
X"38782282",
X"ffff06fe",
X"80800753",
X"b6397b83",
X"38815373",
X"822e0981",
X"06973872",
X"81065372",
X"802e8e38",
X"782281ff",
X"ff068180",
X"80075393",
X"397b9638",
X"fc145372",
X"81268e38",
X"7822ff80",
X"80075372",
X"792380e5",
X"39805573",
X"812e0981",
X"06833873",
X"55775377",
X"802e8938",
X"74810653",
X"7280ca38",
X"72d01554",
X"55728126",
X"83388155",
X"77802eb9",
X"38748106",
X"5372802e",
X"b0387822",
X"83808006",
X"53728380",
X"802e0981",
X"069f3873",
X"b02e0981",
X"06873861",
X"993d3491",
X"3973b12e",
X"09810689",
X"38610284",
X"0580dd05",
X"34618105",
X"538c3961",
X"74318105",
X"53843961",
X"14537283",
X"ffff0642",
X"79f7fb38",
X"7d832a53",
X"72821a34",
X"78228380",
X"80065372",
X"8380802e",
X"09810688",
X"3881537f",
X"872e8338",
X"80537283",
X"c0800c99",
X"3d0d04fd",
X"3d0d7583",
X"11338212",
X"3371982b",
X"71902b07",
X"81143370",
X"882b7207",
X"75337107",
X"83c0800c",
X"52535456",
X"5452853d",
X"0d04f63d",
X"0d02b705",
X"33028405",
X"bb053302",
X"8805bf05",
X"335b5b5b",
X"80588057",
X"78882b7a",
X"07568055",
X"7a548153",
X"a3527c51",
X"92cc3f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f63d",
X"0d02b705",
X"33028405",
X"bb053302",
X"8805bf05",
X"335b5b5b",
X"80588057",
X"78882b7a",
X"07568055",
X"7a548353",
X"a3527c51",
X"92903f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f73d",
X"0d02b305",
X"33028405",
X"b6052260",
X"5a585680",
X"55805480",
X"5381a352",
X"7b5191e2",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8b3d0d04",
X"ee3d0d64",
X"90115c5c",
X"807b3480",
X"0b841c0c",
X"800b881c",
X"34810b89",
X"1c34880b",
X"8a1c3480",
X"0b8b1c34",
X"881b08c1",
X"06810788",
X"1c0c8f3d",
X"70545d88",
X"527b519b",
X"eb3f83c0",
X"800881ff",
X"06705b59",
X"7881a938",
X"903d335e",
X"81db5a7d",
X"892e0981",
X"06819938",
X"7c539252",
X"7b519bc4",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"8182387c",
X"58885778",
X"56a95578",
X"54865381",
X"a0527b51",
X"90d03f83",
X"c0800881",
X"ff06705b",
X"597880e0",
X"3802ba05",
X"337b347c",
X"5478537d",
X"527b519b",
X"ac3f83c0",
X"800881ff",
X"06705b59",
X"7880c138",
X"02bd0533",
X"527b519b",
X"c43f83c0",
X"800881ff",
X"06705b59",
X"78aa3881",
X"7b335a5a",
X"79792699",
X"38805479",
X"5388527b",
X"51fdbb3f",
X"811a7081",
X"ff067c33",
X"525b59e4",
X"39810b88",
X"1c34805a",
X"7983c080",
X"0c943d0d",
X"04800b83",
X"c0800c04",
X"f93d0d79",
X"028405ab",
X"05338e3d",
X"70545858",
X"58ffbeb0",
X"3f8a3d8a",
X"0551ffbe",
X"a73f7551",
X"fc8d3f83",
X"c0800884",
X"86812ebe",
X"3883c080",
X"08848681",
X"26993883",
X"c0800884",
X"82802e80",
X"e63883c0",
X"80088482",
X"812e9f38",
X"81b43983",
X"c0800880",
X"c082832e",
X"80f43883",
X"c0800880",
X"c086832e",
X"80e83881",
X"993983c0",
X"9c335580",
X"5674762e",
X"09810681",
X"8b387454",
X"76539152",
X"7751fbd6",
X"3f745476",
X"53905277",
X"51fbcb3f",
X"74547653",
X"84527751",
X"fbfc3f81",
X"0b83c09c",
X"3481b156",
X"80de3980",
X"54765391",
X"527751fb",
X"a93f8054",
X"76539052",
X"7751fb9e",
X"3f800b83",
X"c09c3476",
X"52871833",
X"5197963f",
X"b5398054",
X"76539452",
X"7751fb82",
X"3f805476",
X"53905277",
X"51faf73f",
X"7551ffbc",
X"db3f83c0",
X"8008892a",
X"81065376",
X"52871833",
X"5190cd3f",
X"800b83c0",
X"9c348056",
X"7583c080",
X"0c893d0d",
X"04f23d0d",
X"6090115a",
X"58800b88",
X"1a337159",
X"56567476",
X"2e82a538",
X"82ac3f84",
X"190883c0",
X"80082682",
X"95387833",
X"5a810b8e",
X"3d23903d",
X"f81155f4",
X"05539918",
X"5277518a",
X"e53f83c0",
X"800881ff",
X"06705755",
X"74772e09",
X"810681d9",
X"38863974",
X"5681d239",
X"81568257",
X"8e3d3377",
X"06557480",
X"2ebb3880",
X"0b8d3d34",
X"903df005",
X"54845375",
X"527751fa",
X"cd3f83c0",
X"800881ff",
X"0655749d",
X"387b5375",
X"527751fc",
X"e73f83c0",
X"800881ff",
X"06557481",
X"b12e818b",
X"3874ffb3",
X"38761081",
X"fc068117",
X"7081ff06",
X"58565787",
X"7627ffa8",
X"38815675",
X"7a2680eb",
X"38800b8d",
X"3d348c3d",
X"70555784",
X"53755277",
X"51f9f73f",
X"83c08008",
X"81ff0655",
X"7480c138",
X"7651ffba",
X"d73f83c0",
X"80088287",
X"06557482",
X"812e0981",
X"06aa3802",
X"ae053381",
X"07557402",
X"8405ae05",
X"347b5375",
X"527751fb",
X"eb3f83c0",
X"800881ff",
X"06557481",
X"b12e9038",
X"74feb838",
X"81167081",
X"ff065755",
X"ff913980",
X"567581ff",
X"0656973f",
X"83c08008",
X"8fd00584",
X"1a0c7557",
X"7683c080",
X"0c903d0d",
X"04049080",
X"a00883c0",
X"800c04ff",
X"3d0d7387",
X"e82951ff",
X"91d33f83",
X"3d0d0404",
X"83caf80b",
X"83c0800c",
X"04fd3d0d",
X"75775454",
X"800b83ca",
X"d834728a",
X"38909080",
X"0b84150c",
X"90397281",
X"2e098106",
X"88389098",
X"800b8415",
X"0c841408",
X"83caf00c",
X"800b8815",
X"0c800b8c",
X"150c83ca",
X"f0085382",
X"0b878014",
X"348151ff",
X"9e3f83ca",
X"f0085380",
X"0b881434",
X"83caf008",
X"53810b87",
X"80143483",
X"caf00853",
X"800b8c14",
X"3483caf0",
X"0853800b",
X"a4143491",
X"7434800b",
X"83c0a034",
X"800b83c0",
X"a434800b",
X"83c0a834",
X"80547381",
X"c42983ca",
X"fc055380",
X"0b831434",
X"81147081",
X"ff065553",
X"8f7427e6",
X"38853d0d",
X"04fe3d0d",
X"74768211",
X"3370bf06",
X"81712bff",
X"05565151",
X"52539071",
X"278338ff",
X"52765171",
X"712383ca",
X"f0085187",
X"13339012",
X"34800b83",
X"c0a43480",
X"0b83c0a8",
X"34881333",
X"8a143352",
X"5271802e",
X"aa387081",
X"ff065184",
X"52708338",
X"70527183",
X"c0a4348a",
X"13337030",
X"70802584",
X"2b708807",
X"51515253",
X"7083c0a8",
X"34903970",
X"81ff0651",
X"70833898",
X"527183c0",
X"a834800b",
X"83c0800c",
X"843d0d04",
X"f13d0d61",
X"6568028c",
X"0580cb05",
X"33029005",
X"80ce0522",
X"02940580",
X"d6052242",
X"40415a40",
X"40fd8b3f",
X"83c08008",
X"a788055b",
X"8070715b",
X"5b528394",
X"3983caf0",
X"08517d94",
X"123483c0",
X"a4338107",
X"55807054",
X"567f8626",
X"80ea387f",
X"842981d8",
X"b40583ca",
X"f0085351",
X"70080480",
X"0b841334",
X"a1397733",
X"70307080",
X"25837131",
X"51515253",
X"70841334",
X"8d39810b",
X"841334b8",
X"39830b84",
X"13348170",
X"5456ad39",
X"810b8413",
X"34a23977",
X"33703070",
X"80258371",
X"31515152",
X"53708413",
X"34807833",
X"52527083",
X"38815271",
X"78348153",
X"74880755",
X"83c0a833",
X"83caf008",
X"5257810b",
X"81d01234",
X"83caf008",
X"51810b81",
X"9012347e",
X"802eae38",
X"72802ea9",
X"387eff1e",
X"52547083",
X"ffff0653",
X"7283ffff",
X"2e973873",
X"70810555",
X"3383caf0",
X"08535170",
X"81c01334",
X"ff1351de",
X"3983caf0",
X"08a81133",
X"53517688",
X"123483ca",
X"f0085174",
X"713481ff",
X"52913983",
X"caf008a0",
X"11337081",
X"06515253",
X"708f38fa",
X"fd3f7a83",
X"c0800826",
X"e6388188",
X"39810ba0",
X"143483ca",
X"f008a811",
X"3380ff06",
X"70780752",
X"53517080",
X"2e80ed38",
X"71862a70",
X"81065151",
X"70802e91",
X"38807833",
X"52537083",
X"38815372",
X"783480e0",
X"3971842a",
X"70810651",
X"5170802e",
X"9b388119",
X"7083ffff",
X"067d3070",
X"9f2a5152",
X"5a51787c",
X"2e098106",
X"af38a439",
X"71832a70",
X"81065151",
X"70802e93",
X"38811a70",
X"81ff065b",
X"5179832e",
X"09810690",
X"388a3971",
X"a3065170",
X"802e8538",
X"71519239",
X"f9e43f7a",
X"83c08008",
X"26fce238",
X"7181bf06",
X"517083c0",
X"800c913d",
X"0d04f63d",
X"0d02b305",
X"33028405",
X"b7053302",
X"8805ba05",
X"22595959",
X"800b8c3d",
X"348c3dfc",
X"05568055",
X"80547653",
X"77527851",
X"fbf23f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f33d",
X"0d7f6264",
X"028c0580",
X"c2052272",
X"22811533",
X"425f415e",
X"59598078",
X"237d5378",
X"33528151",
X"ffa03f83",
X"c0800881",
X"ff065675",
X"802e8638",
X"755481ad",
X"3983caf0",
X"08a81133",
X"821b3370",
X"862a7081",
X"0673982b",
X"5351575c",
X"56577980",
X"25833881",
X"5673762e",
X"873881f0",
X"54818239",
X"818c1733",
X"7081ff06",
X"79227d71",
X"31902b70",
X"902c7009",
X"709f2c72",
X"06705252",
X"53515357",
X"57547574",
X"24833875",
X"55748480",
X"8029fc80",
X"80057090",
X"2c515574",
X"ff2e9438",
X"83caf008",
X"81801133",
X"5154737c",
X"7081055e",
X"34db3977",
X"22760554",
X"73782379",
X"09709f2a",
X"70810682",
X"1c3381bf",
X"0671862b",
X"07515151",
X"5473821a",
X"347c7626",
X"8a387722",
X"547a7426",
X"febb3880",
X"547383c0",
X"800c8f3d",
X"0d04f93d",
X"0d7a5780",
X"0b893d23",
X"893dfc05",
X"53765279",
X"51f8da3f",
X"83c08008",
X"81ff0670",
X"57557496",
X"387c547b",
X"53883d22",
X"527651fd",
X"e53f83c0",
X"800881ff",
X"06567583",
X"c0800c89",
X"3d0d04f0",
X"3d0d6266",
X"02880580",
X"ce052241",
X"5d5e8002",
X"840580d2",
X"05227f81",
X"0533ff11",
X"5a5d5a5d",
X"81da5876",
X"bf2680e9",
X"3878802e",
X"80e1387a",
X"58787b27",
X"83387858",
X"821e3370",
X"872a585a",
X"76923d34",
X"923dfc05",
X"5677557b",
X"547e537d",
X"33528251",
X"f8de3f83",
X"c0800881",
X"ff065d80",
X"0b923d33",
X"585a7680",
X"2e833881",
X"5a821e33",
X"80ff067a",
X"872b0757",
X"76821f34",
X"7c913878",
X"78317083",
X"ffff0679",
X"1e5e5a57",
X"ff9b397c",
X"587783c0",
X"800c923d",
X"0d04f83d",
X"0d7b0284",
X"05b20522",
X"5858800b",
X"8a3d238a",
X"3dfc0553",
X"77527a51",
X"f6f73f83",
X"c0800881",
X"ff067057",
X"55749638",
X"7d547653",
X"893d2252",
X"7751feaf",
X"3f83c080",
X"0881ff06",
X"567583c0",
X"800c8a3d",
X"0d04ec3d",
X"0d666e02",
X"880580df",
X"0533028c",
X"0580e305",
X"33029005",
X"80e70533",
X"02940580",
X"eb053302",
X"980580ee",
X"05224143",
X"415f5c40",
X"570280f2",
X"0522963d",
X"23963df0",
X"05538417",
X"70537752",
X"59f6863f",
X"83c08008",
X"81ff0658",
X"7781e538",
X"777a8180",
X"06584080",
X"77258338",
X"81407994",
X"3d347b02",
X"840580c9",
X"05347c02",
X"840580ca",
X"05347d02",
X"840580cb",
X"05347a95",
X"3d347a88",
X"2a577602",
X"840580cd",
X"0534953d",
X"22577602",
X"840580ce",
X"05347688",
X"2a577602",
X"840580cf",
X"05347792",
X"3d34963d",
X"ec115757",
X"8855f417",
X"54923d22",
X"53775277",
X"51f6953f",
X"83c08008",
X"81ff0658",
X"7780ed38",
X"7e802e80",
X"cb38923d",
X"22790858",
X"587f802e",
X"9c387681",
X"80800779",
X"0c7e5496",
X"3dfc0553",
X"7783ffff",
X"06527851",
X"f9fc3f99",
X"39768280",
X"8007790c",
X"7e54953d",
X"22537783",
X"ffff0652",
X"7851fc8f",
X"3f83c080",
X"0881ff06",
X"58779d38",
X"923d2253",
X"80527f30",
X"70802584",
X"71315351",
X"57f9873f",
X"83c08008",
X"81ff0658",
X"7783c080",
X"0c963d0d",
X"04f63d0d",
X"7c028405",
X"b705335b",
X"5b805880",
X"57805680",
X"55795485",
X"5380527a",
X"51fda33f",
X"83c08008",
X"81ff0659",
X"78853879",
X"871c3478",
X"83c0800c",
X"8c3d0d04",
X"f93d0d02",
X"a7053302",
X"8405ab05",
X"33028805",
X"af053358",
X"5957800b",
X"83caff33",
X"54547274",
X"2e9f3881",
X"147081ff",
X"06555373",
X"8f2681b6",
X"387381c4",
X"2983cafc",
X"05831133",
X"515372e3",
X"387381c4",
X"2983caf8",
X"0555800b",
X"87163476",
X"88163475",
X"8a163477",
X"89163480",
X"750c83ca",
X"f0088c16",
X"0c800b84",
X"1634880b",
X"85163480",
X"0b861634",
X"841508ff",
X"a1ff06a0",
X"80078416",
X"0c811470",
X"81ff0653",
X"537451fe",
X"bc3f83c0",
X"800881ff",
X"06705553",
X"7280cd38",
X"8a397308",
X"750c7254",
X"80c23972",
X"81ddd455",
X"5681ddd4",
X"08802eb2",
X"38758429",
X"14700876",
X"53700851",
X"5454722d",
X"83c08008",
X"81ff0653",
X"72802ece",
X"38811670",
X"81ff0681",
X"ddd47184",
X"29115356",
X"57537208",
X"d0388054",
X"7383c080",
X"0c893d0d",
X"04f93d0d",
X"7957800b",
X"84180883",
X"caf00c58",
X"f0883f88",
X"170883c0",
X"80082783",
X"ed38effa",
X"3f83c080",
X"08810588",
X"180c83ca",
X"f008b811",
X"337081ff",
X"06515154",
X"73812ea4",
X"38738124",
X"88387378",
X"2e8a38b8",
X"3973822e",
X"9538b139",
X"763381f0",
X"06547390",
X"2ea63891",
X"7734a139",
X"73587633",
X"81f00654",
X"73902e09",
X"81069138",
X"efa83f83",
X"c0800881",
X"c8058c18",
X"0ca07734",
X"80567581",
X"c42983ca",
X"ff113355",
X"5573802e",
X"aa3883ca",
X"f8157008",
X"56547480",
X"2e9d3888",
X"1508802e",
X"96388c14",
X"0883caf0",
X"082e0981",
X"06893873",
X"51881508",
X"54732d81",
X"167081ff",
X"0657548f",
X"7627ffba",
X"38763354",
X"73b02e81",
X"993873b0",
X"248f3873",
X"912eab38",
X"73a02e80",
X"f53882a6",
X"397380d0",
X"2e81e438",
X"7380d024",
X"8b387380",
X"c02e8199",
X"38828f39",
X"7381802e",
X"81fb3882",
X"85398056",
X"7581c429",
X"83cafc11",
X"83113356",
X"59557380",
X"2ea83883",
X"caf81570",
X"08565474",
X"802e9b38",
X"8c140883",
X"caf0082e",
X"0981068e",
X"38735184",
X"15085473",
X"2d800b83",
X"19348116",
X"7081ff06",
X"57548f76",
X"27ffb938",
X"92773481",
X"b539edc2",
X"3f8c1708",
X"83c08008",
X"2781a738",
X"b0773481",
X"a13983ca",
X"f0085480",
X"0b8c1534",
X"83caf008",
X"54840b88",
X"153480c0",
X"7734ed96",
X"3f83c080",
X"08b2058c",
X"180c80fa",
X"39ed873f",
X"8c170883",
X"c0800827",
X"80ec3883",
X"caf00854",
X"810b8c15",
X"3483caf0",
X"0854800b",
X"88153483",
X"caf00854",
X"880ba015",
X"34ecdb3f",
X"83c08008",
X"94058c18",
X"0c80d077",
X"34bc3983",
X"caf008a0",
X"11337083",
X"2a708106",
X"51515555",
X"73802ea6",
X"38880ba0",
X"1634ecae",
X"3f8c1708",
X"83c08008",
X"279438ff",
X"8077348e",
X"39775380",
X"528051fa",
X"8b3fff90",
X"773483ca",
X"f008a011",
X"3370832a",
X"70810651",
X"51555573",
X"802e8638",
X"880ba016",
X"34893d0d",
X"04f63d0d",
X"02b30533",
X"028405b7",
X"05335b5b",
X"800b83ca",
X"fc708412",
X"72745d59",
X"575b5856",
X"83153353",
X"72802e80",
X"f3387333",
X"537a732e",
X"09810680",
X"e7388114",
X"33537973",
X"2e098106",
X"80da3880",
X"557481c4",
X"2983cb80",
X"05703383",
X"1b335855",
X"5373762e",
X"0981068a",
X"38811333",
X"527351ff",
X"9c3f8115",
X"7081ff06",
X"56538f75",
X"27d33880",
X"0b83caf8",
X"19700856",
X"54557375",
X"2e913872",
X"51841408",
X"53722d83",
X"c0800881",
X"ff065580",
X"0b831834",
X"7453a039",
X"811681c4",
X"1981c417",
X"81c41781",
X"c41d81c4",
X"1c5c5d57",
X"5759568f",
X"7625fee8",
X"38805372",
X"83c0800c",
X"8c3d0d04",
X"f83d0d02",
X"ae05227d",
X"59578056",
X"81558054",
X"86538180",
X"527a51f5",
X"953f83c0",
X"800881ff",
X"0683c080",
X"0c8a3d0d",
X"04f73d0d",
X"02b20522",
X"028405b7",
X"0533605a",
X"5b578056",
X"82557954",
X"86538180",
X"527b51f4",
X"e53f83c0",
X"800881ff",
X"0683c080",
X"0c8b3d0d",
X"04f83d0d",
X"02af0533",
X"59805880",
X"57805680",
X"55785489",
X"5380527a",
X"51f4bb3f",
X"83c08008",
X"81ff0683",
X"c0800c8a",
X"3d0d0400",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002b20",
X"00002b61",
X"00002b83",
X"00002baa",
X"00002baa",
X"00002baa",
X"00002baa",
X"00002c1b",
X"00002c6d",
X"00004190",
X"000049d4",
X"00004a8d",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3f00",
X"0c0c4000",
X"0a0a4100",
X"0b0b4100",
X"07074100",
X"0a0b4300",
X"080b4200",
X"04044500",
X"05054400",
X"06060004",
X"08080004",
X"09090004",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"00005719",
X"00005a20",
X"0000582c",
X"00005a20",
X"00005869",
X"000058ba",
X"000058f9",
X"00005902",
X"00005a20",
X"00005a20",
X"00005a20",
X"00005a20",
X"0000590b",
X"00005913",
X"0000591a",
X"00005b20",
X"00005c19",
X"00005d2d",
X"00006023",
X"0000603e",
X"0000602a",
X"0000603e",
X"00006045",
X"00006050",
X"00006057",
X"25732025",
X"73000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"66726565",
X"7a65722e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"6e616d65",
X"20000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00006c8c",
X"00006c90",
X"00006c98",
X"00006ca4",
X"00006cb0",
X"00006cbc",
X"00006cc8",
X"00006ccc",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00006c28",
X"00006a7c",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"69383030",
X"00000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
