-- megafunction wizard: %ALTIOBUF%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altiobuf_out 

-- ============================================================
-- File Name: altiobufo.vhd
-- Megafunction Name(s):
-- 			altiobuf_out
--
-- Simulation Library Files(s):
-- 			cyclonev
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 14.0.0 Build 200 06/17/2014 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus II License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


--altiobuf_out CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" ENABLE_BUS_HOLD="FALSE" LEFT_SHIFT_SERIES_TERMINATION_CONTROL="FALSE" NUMBER_OF_CHANNELS=1 OPEN_DRAIN_OUTPUT="FALSE" PSEUDO_DIFFERENTIAL_MODE="TRUE" USE_DIFFERENTIAL_MODE="TRUE" USE_OE="TRUE" USE_TERMINATION_CONTROL="FALSE" datain dataout dataout_b oe oe_b
--VERSION_BEGIN 14.0 cbx_altiobuf_out 2014:06:05:09:45:41:SJ cbx_mgl 2014:06:05:10:17:12:SJ cbx_stratixiii 2014:06:05:09:45:41:SJ cbx_stratixv 2014:06:05:09:45:41:SJ  VERSION_END

 LIBRARY cyclonev;
 USE cyclonev.all;

--synthesis_resources = cyclonev_io_obuf 2 cyclonev_pseudo_diff_out 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altiobufo_iobuf_out_h5u IS 
	 PORT 
	 ( 
		 datain	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 dataout	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 dataout_b	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 oe	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '1');
		 oe_b	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '1')
	 ); 
 END altiobufo_iobuf_out_h5u;

 ARCHITECTURE RTL OF altiobufo_iobuf_out_h5u IS

	 SIGNAL  wire_obuf_ba_o	:	STD_LOGIC;
	 SIGNAL  wire_obuf_ba_oe	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pseudo_diffa_w_lg_oebout3w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_obufa_o	:	STD_LOGIC;
	 SIGNAL  wire_obufa_oe	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pseudo_diffa_w_lg_oeout2w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pseudo_diffa_o	:	STD_LOGIC;
	 SIGNAL  wire_pseudo_diffa_obar	:	STD_LOGIC;
	 SIGNAL  wire_pseudo_diffa_oebout	:	STD_LOGIC;
	 SIGNAL  wire_pseudo_diffa_oein	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_oe_w1w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pseudo_diffa_oeout	:	STD_LOGIC;
	 SIGNAL  oe_w :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  cyclonev_io_obuf
	 GENERIC 
	 (
		bus_hold	:	STRING := "false";
		open_drain_output	:	STRING := "false";
		shift_series_termination_control	:	STRING := "false";
		lpm_type	:	STRING := "cyclonev_io_obuf"
	 );
	 PORT
	 ( 
		dynamicterminationcontrol	:	IN STD_LOGIC := '0';
		i	:	IN STD_LOGIC := '0';
		o	:	OUT STD_LOGIC;
		obar	:	OUT STD_LOGIC;
		oe	:	IN STD_LOGIC := '1';
		parallelterminationcontrol	:	IN STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
		seriesterminationcontrol	:	IN STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  cyclonev_pseudo_diff_out
	 PORT
	 ( 
		dtc	:	OUT STD_LOGIC;
		dtcbar	:	OUT STD_LOGIC;
		dtcin	:	IN STD_LOGIC := '0';
		i	:	IN STD_LOGIC := '0';
		o	:	OUT STD_LOGIC;
		obar	:	OUT STD_LOGIC;
		oebout	:	OUT STD_LOGIC;
		oein	:	IN STD_LOGIC := '0';
		oeout	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	dataout(0) <= wire_obufa_o;
	dataout_b(0) <= wire_obuf_ba_o;
	oe_w <= oe;
	wire_obuf_ba_oe <= wire_pseudo_diffa_w_lg_oebout3w;
	wire_pseudo_diffa_w_lg_oebout3w(0) <= NOT wire_pseudo_diffa_oebout;
	obuf_ba :  cyclonev_io_obuf
	  GENERIC MAP (
		bus_hold => "false",
		open_drain_output => "false"
	  )
	  PORT MAP ( 
		i => wire_pseudo_diffa_obar,
		o => wire_obuf_ba_o,
		oe => wire_obuf_ba_oe(0)
	  );
	wire_obufa_oe <= wire_pseudo_diffa_w_lg_oeout2w;
	wire_pseudo_diffa_w_lg_oeout2w(0) <= NOT wire_pseudo_diffa_oeout;
	obufa :  cyclonev_io_obuf
	  GENERIC MAP (
		bus_hold => "false",
		open_drain_output => "false"
	  )
	  PORT MAP ( 
		i => wire_pseudo_diffa_o,
		o => wire_obufa_o,
		oe => wire_obufa_oe(0)
	  );
	wire_pseudo_diffa_oein <= wire_w_lg_oe_w1w;
	wire_w_lg_oe_w1w(0) <= NOT oe_w(0);
	pseudo_diffa :  cyclonev_pseudo_diff_out
	  PORT MAP ( 
		i => datain(0),
		o => wire_pseudo_diffa_o,
		obar => wire_pseudo_diffa_obar,
		oebout => wire_pseudo_diffa_oebout,
		oein => wire_pseudo_diffa_oein(0),
		oeout => wire_pseudo_diffa_oeout
	  );

 END RTL; --altiobufo_iobuf_out_h5u
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY altiobufo IS
	PORT
	(
		datain		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		oe		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		oe_b		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		dataout		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		dataout_b		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0)
	);
END altiobufo;


ARCHITECTURE RTL OF altiobufo IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (0 DOWNTO 0);



	COMPONENT altiobufo_iobuf_out_h5u
	PORT (
			datain	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			oe	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			oe_b	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			dataout	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			dataout_b	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	dataout    <= sub_wire0(0 DOWNTO 0);
	dataout_b    <= sub_wire1(0 DOWNTO 0);

	altiobufo_iobuf_out_h5u_component : altiobufo_iobuf_out_h5u
	PORT MAP (
		datain => datain,
		oe => oe,
		oe_b => oe_b,
		dataout => sub_wire0,
		dataout_b => sub_wire1
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: enable_bus_hold STRING "FALSE"
-- Retrieval info: CONSTANT: left_shift_series_termination_control STRING "FALSE"
-- Retrieval info: CONSTANT: number_of_channels NUMERIC "1"
-- Retrieval info: CONSTANT: open_drain_output STRING "FALSE"
-- Retrieval info: CONSTANT: pseudo_differential_mode STRING "TRUE"
-- Retrieval info: CONSTANT: use_differential_mode STRING "TRUE"
-- Retrieval info: CONSTANT: use_oe STRING "TRUE"
-- Retrieval info: CONSTANT: use_termination_control STRING "FALSE"
-- Retrieval info: USED_PORT: datain 0 0 1 0 INPUT NODEFVAL "datain[0..0]"
-- Retrieval info: USED_PORT: dataout 0 0 1 0 OUTPUT NODEFVAL "dataout[0..0]"
-- Retrieval info: USED_PORT: dataout_b 0 0 1 0 OUTPUT NODEFVAL "dataout_b[0..0]"
-- Retrieval info: USED_PORT: oe 0 0 1 0 INPUT NODEFVAL "oe[0..0]"
-- Retrieval info: USED_PORT: oe_b 0 0 1 0 INPUT NODEFVAL "oe_b[0..0]"
-- Retrieval info: CONNECT: @datain 0 0 1 0 datain 0 0 1 0
-- Retrieval info: CONNECT: @oe 0 0 1 0 oe 0 0 1 0
-- Retrieval info: CONNECT: @oe_b 0 0 1 0 oe_b 0 0 1 0
-- Retrieval info: CONNECT: dataout 0 0 1 0 @dataout 0 0 1 0
-- Retrieval info: CONNECT: dataout_b 0 0 1 0 @dataout_b 0 0 1 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altiobufo.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altiobufo.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altiobufo.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altiobufo.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altiobufo_inst.vhd FALSE
-- Retrieval info: LIB_FILE: cyclonev
