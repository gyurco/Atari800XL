
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f8",
X"bc738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80fc",
X"9c0c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f2",
X"ea2d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580f0fe",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"96d20480",
X"3d0d80fd",
X"c0087008",
X"810683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d80fd",
X"c0087008",
X"70fe0676",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80fdc008",
X"70087081",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80fdc008",
X"700870fd",
X"06761007",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"fdc00870",
X"0870822c",
X"bf0683e0",
X"800c5151",
X"823d0d04",
X"ff3d0d80",
X"fdc00870",
X"0870fe83",
X"0676822b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80fdc008",
X"70087088",
X"2c870683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80fdc008",
X"700870f1",
X"ff067688",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d80fdc0",
X"08700870",
X"8b2cbf06",
X"83e0800c",
X"5151823d",
X"0d04ff3d",
X"0d80fdc0",
X"08700870",
X"f88fff06",
X"768b2b07",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"fdd00870",
X"0870882c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fdd00870",
X"0870892c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fdd00870",
X"08708a2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fdd00870",
X"08708b2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"fd3d0d75",
X"81e62987",
X"2a80fdb0",
X"0854730c",
X"853d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d848080",
X"53805288",
X"800a51ff",
X"b33f8180",
X"80538052",
X"82800a51",
X"c63f843d",
X"0d04803d",
X"0d8151fc",
X"fc3f7280",
X"2e8338d2",
X"3f8051fc",
X"f03f8051",
X"fcbd3f82",
X"3d0d04fd",
X"3d0d7552",
X"805480ff",
X"72258838",
X"810bff80",
X"135354ff",
X"bf125170",
X"99268638",
X"e012529e",
X"39ff9f12",
X"51997127",
X"9538d012",
X"e0137054",
X"54518971",
X"2788388f",
X"73278338",
X"80527380",
X"2e853881",
X"80125271",
X"81ff0683",
X"e0800c85",
X"3d0d0480",
X"3d0d86b8",
X"c0518071",
X"70810553",
X"347086c0",
X"c02e0981",
X"06f03882",
X"3d0d04fe",
X"3d0d0297",
X"053351ff",
X"863f83e0",
X"800881ff",
X"0683e09c",
X"08545280",
X"73249b38",
X"83e0b408",
X"137283e0",
X"b8080753",
X"53717334",
X"83e09c08",
X"810583e0",
X"9c0c843d",
X"0d04fa3d",
X"0d82800a",
X"1b558057",
X"883dfc05",
X"54795374",
X"527851b7",
X"b63f883d",
X"0d04fe3d",
X"0d83e0b0",
X"08527451",
X"bdf03f83",
X"e080088c",
X"38765375",
X"5283e0b0",
X"0851c73f",
X"843d0d04",
X"fe3d0d83",
X"e0b00853",
X"75527451",
X"b8b73f83",
X"e080088d",
X"38775376",
X"5283e0b0",
X"0851ffa2",
X"3f843d0d",
X"04803d0d",
X"fb9b3f83",
X"e0800887",
X"2680cd38",
X"83e08008",
X"842980f8",
X"cc055170",
X"08040b0b",
X"80f9b451",
X"b7390b0b",
X"80f9b851",
X"af390b0b",
X"80f9c051",
X"a7390b0b",
X"80f9cc51",
X"9f390b0b",
X"80f9d851",
X"97390b0b",
X"80f9e451",
X"8f390b0b",
X"80f9f051",
X"87390b0b",
X"80f9f451",
X"7083e080",
X"0c823d0d",
X"04ee3d0d",
X"80438042",
X"80418070",
X"5a5bfdd3",
X"3f800b83",
X"e09c0c80",
X"0b83e0b8",
X"0c0b0b80",
X"f9f851b1",
X"ef3f8180",
X"0b83e0b8",
X"0c0b0b80",
X"f9fc51b1",
X"df3f80d0",
X"0b83e09c",
X"0c783070",
X"7a078025",
X"70872b83",
X"e0b80c51",
X"55f9bd3f",
X"83e08008",
X"520b0b80",
X"fa8451b1",
X"b73f80f8",
X"0b83e09c",
X"0c788132",
X"70307072",
X"07802570",
X"872b83e0",
X"b80c5156",
X"56fea23f",
X"83e08008",
X"520b0b80",
X"fa9051b1",
X"8b3f81a0",
X"0b83e09c",
X"0c788232",
X"70307072",
X"07802570",
X"872b83e0",
X"b80c5156",
X"56f9c73f",
X"83e08008",
X"520b0b80",
X"fa9851b0",
X"df3f81f0",
X"0b83e09c",
X"0c810b83",
X"e0a05b58",
X"83e09c08",
X"82197a32",
X"70307072",
X"07802570",
X"872b83e0",
X"b80c5157",
X"8e3d7055",
X"ff1b5457",
X"5757a6bd",
X"3f797084",
X"055b0851",
X"b28b3f74",
X"5483e080",
X"08537752",
X"0b0b80fa",
X"a451b090",
X"3fa81783",
X"e09c0c81",
X"18587785",
X"2e098106",
X"ffae3883",
X"900b83e0",
X"9c0c7887",
X"32703070",
X"72078025",
X"70872b83",
X"e0b80c51",
X"560b0b80",
X"fab45256",
X"afda3f83",
X"e00b83e0",
X"9c0c7888",
X"32703070",
X"72078025",
X"70872b83",
X"e0b80c51",
X"560b0b80",
X"fac85256",
X"afb63f86",
X"8da051f9",
X"9b3f8052",
X"913d7052",
X"558cbc3f",
X"83527451",
X"8cb53f61",
X"19597880",
X"25853880",
X"59903988",
X"79258538",
X"88598739",
X"78882682",
X"a1387882",
X"2b5580f8",
X"ec150804",
X"f6ee3f83",
X"e0800861",
X"57557581",
X"2e098106",
X"893883e0",
X"80081055",
X"903975ff",
X"2e098106",
X"883883e0",
X"8008812c",
X"55907525",
X"85389055",
X"88397480",
X"24833881",
X"557451f6",
X"cb3f81d6",
X"39f6de3f",
X"83e08008",
X"61055574",
X"80258538",
X"80558839",
X"87752583",
X"38875574",
X"51f6da3f",
X"81b439f6",
X"ed3f83e0",
X"80086105",
X"55748024",
X"85388155",
X"88398675",
X"25833886",
X"557451f6",
X"e93f8192",
X"39605680",
X"76259838",
X"a18b0b83",
X"e0cc0c83",
X"e0941570",
X"0852558d",
X"e43f7408",
X"52913975",
X"80259138",
X"83e09415",
X"0851afc3",
X"3f8052fd",
X"1951a739",
X"62802e80",
X"d93883e0",
X"a00883e0",
X"94167008",
X"83e0a00c",
X"71710c56",
X"52fd1951",
X"95813f83",
X"e0a00852",
X"805194f7",
X"3fb43962",
X"802eaf38",
X"a1ec0b83",
X"e0cc0c83",
X"e0b00851",
X"8d8b3f83",
X"e0b00851",
X"aee33f9c",
X"800a5380",
X"c0805283",
X"e0800851",
X"f9ac3f81",
X"558c3962",
X"87387a80",
X"2efad738",
X"80557483",
X"e0800c94",
X"3d0d04fe",
X"3d0df5d8",
X"3f83e080",
X"08802e86",
X"38805180",
X"f639f5e0",
X"3f83e080",
X"0880ea38",
X"f6863f83",
X"e0800880",
X"2eaa3881",
X"51f3d83f",
X"84903f80",
X"0b83e09c",
X"0cfa863f",
X"83e08008",
X"53ff0b83",
X"e09c0c86",
X"e33f72bd",
X"387251f3",
X"b63fbb39",
X"f5ba3f83",
X"e0800880",
X"2eb03881",
X"51f3a43f",
X"83dc3fa1",
X"8b0b83e0",
X"cc0c83e0",
X"a008518b",
X"e83fff0b",
X"83e09c0c",
X"86ae3f83",
X"e0a00852",
X"805193ab",
X"3f8151f6",
X"a53f843d",
X"0d0483e0",
X"8c080283",
X"e08c0cfa",
X"3d0d800b",
X"83e0a00b",
X"83e08c08",
X"fc050c83",
X"e08c08f8",
X"050cb08b",
X"3f83e080",
X"088605fc",
X"0683e08c",
X"08f4050c",
X"0283e08c",
X"08f40508",
X"310d853d",
X"7083e08c",
X"08fc0508",
X"70840583",
X"e08c08fc",
X"050c0c51",
X"ace93f83",
X"e08c08f8",
X"05088105",
X"83e08c08",
X"f8050c83",
X"e08c08f8",
X"0508852e",
X"098106ff",
X"ad388688",
X"80805182",
X"9f3fff0b",
X"83e09c0c",
X"800b83e0",
X"b80c86b8",
X"c00b83e0",
X"b40c8151",
X"f28f3f81",
X"51f2b93f",
X"8251f396",
X"3f8251f2",
X"e03f8dff",
X"528051aa",
X"8c3f8480",
X"80528684",
X"808051af",
X"f23f83e0",
X"800881d2",
X"3895d43f",
X"0b0b80fa",
X"d051b4a8",
X"3f83e080",
X"0883e08c",
X"08f4050c",
X"83c18080",
X"54818080",
X"530b0b80",
X"fae85283",
X"e0800851",
X"f6ba3f83",
X"c2808054",
X"81808053",
X"0b0b80fa",
X"f45283e0",
X"8c08f405",
X"0851f6a0",
X"3f83c380",
X"80548180",
X"80530b0b",
X"80fb8052",
X"83e08c08",
X"f4050851",
X"f6863f83",
X"c4808054",
X"81808053",
X"0b0b80fb",
X"8c5283e0",
X"8c08f405",
X"0851f5ec",
X"3f83c5b0",
X"805480d0",
X"80530b0b",
X"80fb9852",
X"83e08c08",
X"f4050851",
X"f5d23f83",
X"c6b08054",
X"80d08053",
X"0b0b80fb",
X"a45283e0",
X"8c08f405",
X"0851f5b8",
X"3f9c800a",
X"5480c080",
X"530b0b80",
X"fbb05283",
X"e08c08f4",
X"050851f5",
X"9f3f8151",
X"f3943f9e",
X"bc3f8151",
X"f38c3ffb",
X"da3ffc39",
X"7183e0c0",
X"0c888080",
X"0b83e0bc",
X"0c848080",
X"0b83e0c4",
X"0c04f03d",
X"0d80fcb8",
X"08547333",
X"83e0c834",
X"83a08056",
X"83e0c008",
X"1683e0bc",
X"08175654",
X"74337434",
X"83e0c408",
X"16548074",
X"34811656",
X"7583a0a0",
X"2e098106",
X"db3883a4",
X"805683e0",
X"c0081683",
X"e0bc0817",
X"56547433",
X"743483e0",
X"c4081654",
X"80743481",
X"16567583",
X"a4a02e09",
X"8106db38",
X"83a88056",
X"83e0c008",
X"1683e0bc",
X"08175654",
X"74337434",
X"83e0c408",
X"16548074",
X"34811656",
X"7583a890",
X"2e098106",
X"db3880fc",
X"b80854ff",
X"74348056",
X"83e0c008",
X"1683e0c4",
X"08175555",
X"73337534",
X"81165675",
X"83a0802e",
X"098106e4",
X"3883b080",
X"5683e0c0",
X"081683e0",
X"c4081755",
X"55733375",
X"34811656",
X"75848080",
X"2e098106",
X"e438f28b",
X"3f893d58",
X"a25380f9",
X"90527751",
X"80dbb83f",
X"80578c80",
X"5683e0c4",
X"08167719",
X"55557333",
X"75348116",
X"81185856",
X"76a22e09",
X"8106e638",
X"80fcdc08",
X"54867434",
X"80fce008",
X"54807434",
X"80fcd808",
X"54807434",
X"80fcc808",
X"54af7434",
X"80fcd408",
X"54bf7434",
X"80fcd008",
X"54807434",
X"80fccc08",
X"549f7434",
X"80fcc408",
X"54807434",
X"80fcb008",
X"54e07434",
X"80fca808",
X"54767434",
X"80fca408",
X"54837434",
X"80fcac08",
X"54827434",
X"923d0d04",
X"fe3d0d80",
X"5383e0c4",
X"081383e0",
X"c0081452",
X"52703372",
X"34811353",
X"7283a080",
X"2e098106",
X"e43883b0",
X"805383e0",
X"c4081383",
X"e0c00814",
X"52527033",
X"72348113",
X"53728480",
X"802e0981",
X"06e43883",
X"a0805383",
X"e0c40813",
X"83e0c008",
X"14525270",
X"33723481",
X"13537283",
X"a0a02e09",
X"8106e438",
X"83a48053",
X"83e0c408",
X"1383e0c0",
X"08145252",
X"70337234",
X"81135372",
X"83a4a02e",
X"098106e4",
X"3883a880",
X"5383e0c4",
X"081383e0",
X"c0081452",
X"52703372",
X"34811353",
X"7283a890",
X"2e098106",
X"e43880fc",
X"b8085183",
X"e0c83371",
X"34843d0d",
X"04fe3d0d",
X"74538073",
X"0c800b84",
X"140c800b",
X"88140c80",
X"fcbc0870",
X"337081ff",
X"0670812a",
X"81327081",
X"06515254",
X"51517080",
X"2e883881",
X"0b84140c",
X"93397181",
X"32708106",
X"51517080",
X"2e8638ff",
X"0b84140c",
X"71832a81",
X"32708106",
X"51517080",
X"2e863881",
X"730c9339",
X"71822a81",
X"32708106",
X"51517080",
X"2e8438ff",
X"730c80fc",
X"b4087033",
X"70097081",
X"06515151",
X"5170802e",
X"8638810b",
X"88140c84",
X"3d0d04fe",
X"3d0d7476",
X"54527151",
X"feeb3f72",
X"812ea238",
X"8173268d",
X"3872822e",
X"ab387283",
X"2e9f38e6",
X"397108e2",
X"38841208",
X"dd388812",
X"08d838a0",
X"39881208",
X"812e0981",
X"06cc3894",
X"39881208",
X"812e8d38",
X"71088938",
X"84120880",
X"2effb738",
X"843d0d04",
X"ffb83d0d",
X"800b80cc",
X"3d08538b",
X"3d705359",
X"5480c6ed",
X"3f80cc3d",
X"085280ca",
X"3dfdfc05",
X"5180c6dd",
X"3f893d33",
X"028405a1",
X"05330288",
X"05a20533",
X"59575573",
X"18703351",
X"5372802e",
X"be3872ae",
X"2e863881",
X"1454ec39",
X"80ca3dfe",
X"81111570",
X"33515458",
X"74732e09",
X"8106a038",
X"fe821814",
X"70335153",
X"75732e09",
X"81069038",
X"fe831814",
X"53817333",
X"54547673",
X"2e833880",
X"547383e0",
X"800c80ca",
X"3d0d04fc",
X"3d0d7670",
X"5255ac9e",
X"3f83e080",
X"08548153",
X"83e08008",
X"80c13874",
X"51abe13f",
X"83e08008",
X"80fbd053",
X"83e08008",
X"5253fec8",
X"3f83e080",
X"08a13880",
X"fbd45272",
X"51feb93f",
X"83e08008",
X"923880fb",
X"d8527251",
X"feaa3f83",
X"e0800880",
X"2e833881",
X"54735372",
X"83e0800c",
X"863d0d04",
X"fd3d0d75",
X"705254ab",
X"bd3f8153",
X"83e08008",
X"97387351",
X"ab863f80",
X"fbdc5283",
X"e0800851",
X"fdf23f83",
X"e0800853",
X"7283e080",
X"0c853d0d",
X"04e03d0d",
X"a33d0870",
X"525ea1d5",
X"3f83e080",
X"0833943d",
X"56547399",
X"388f5380",
X"fbe05274",
X"5180d4df",
X"3f9a397d",
X"527851a4",
X"be3f84db",
X"397d51a1",
X"b83f83e0",
X"80085274",
X"51a0e83f",
X"83e0cc08",
X"52933d70",
X"525ba79b",
X"3f83e080",
X"0859800b",
X"83e08008",
X"555c83e0",
X"80087c2e",
X"9438811c",
X"74525caa",
X"9c3f83e0",
X"80085483",
X"e08008ee",
X"38805aff",
X"7a437a42",
X"7a415f79",
X"09709f2c",
X"7b065b54",
X"7b7a2484",
X"38ff1c5a",
X"f61a7009",
X"709f2c72",
X"067bff12",
X"5a5a5255",
X"55807525",
X"95387651",
X"a9db3f83",
X"e0800876",
X"ff185855",
X"57738024",
X"ed38747f",
X"2e8638ea",
X"863f745f",
X"78ff1b70",
X"585e5880",
X"7a259538",
X"7751a9b1",
X"3f83e080",
X"0876ff18",
X"58555873",
X"8024ed38",
X"800b83e0",
X"9c0c800b",
X"83e0b80c",
X"80fbf051",
X"9e823f81",
X"800b83e0",
X"b80c80fb",
X"f8519df4",
X"3fa80b83",
X"e09c0c76",
X"802e80e4",
X"3883e09c",
X"08777932",
X"70307072",
X"07802570",
X"872b83e0",
X"b80c5156",
X"78535656",
X"a8e83f83",
X"e0800880",
X"2e883880",
X"fc80519d",
X"bb3f7651",
X"a8aa3f83",
X"e0800852",
X"80fab051",
X"9daa3f76",
X"51a8b23f",
X"83e08008",
X"83e09c08",
X"55577574",
X"258638a8",
X"1656f739",
X"7583e09c",
X"0c86f076",
X"24ff9838",
X"87980b83",
X"e09c0c77",
X"802eb138",
X"7751a7e8",
X"3f83e080",
X"08785255",
X"a8883f80",
X"fc885483",
X"e080088d",
X"38873980",
X"7634fda0",
X"3980fae4",
X"54745373",
X"5280fbc0",
X"519cc93f",
X"805480fc",
X"90519cc0",
X"3f811454",
X"73a82e09",
X"8106ef38",
X"868da051",
X"e69a3f80",
X"52903d70",
X"5254f9bb",
X"3f835273",
X"51f9b43f",
X"61802e81",
X"9c387c54",
X"73ff2e96",
X"3878802e",
X"819d3878",
X"51a7923f",
X"83e08008",
X"ff155559",
X"e7397880",
X"2e818838",
X"7851a78e",
X"3f83e080",
X"08802efc",
X"96387851",
X"a6d63f83",
X"e0800883",
X"e0800853",
X"80fbc852",
X"54bffe3f",
X"83e08008",
X"a5387a51",
X"80c1b53f",
X"83e08008",
X"5574ff16",
X"56548074",
X"25fbfd38",
X"741b7033",
X"555673af",
X"2efecc38",
X"e8397a51",
X"80c1913f",
X"825380fb",
X"cc5283e0",
X"80081b51",
X"80d09c3f",
X"7a5180c0",
X"fb3f7352",
X"83e08008",
X"1b5180c0",
X"d33ffbc4",
X"397f8829",
X"6010057a",
X"0561055a",
X"fbf539a2",
X"3d0d0480",
X"3d0d81ff",
X"51800b83",
X"e0d81234",
X"ff115170",
X"f438823d",
X"0d04ff3d",
X"0d737033",
X"53518111",
X"33713471",
X"81123483",
X"3d0d04fb",
X"3d0d7779",
X"56568070",
X"71555552",
X"717525ac",
X"38721670",
X"33701470",
X"81ff0655",
X"51515171",
X"74278938",
X"81127081",
X"ff065351",
X"71811470",
X"83ffff06",
X"55525474",
X"7324d638",
X"7183e080",
X"0c873d0d",
X"04fd3d0d",
X"755494a6",
X"3f83e080",
X"08802ef6",
X"3883e2f4",
X"08860570",
X"81ff0652",
X"5391ff3f",
X"8439ed83",
X"3f94873f",
X"83e08008",
X"812ef338",
X"92e23f83",
X"e0800874",
X"3492d93f",
X"83e08008",
X"81153492",
X"cf3f83e0",
X"80088215",
X"3492c53f",
X"83e08008",
X"83153492",
X"bb3f83e0",
X"80088415",
X"348439ec",
X"c23f93c6",
X"3f83e080",
X"08802ef3",
X"38733383",
X"e0d83481",
X"143383e0",
X"d9348214",
X"3383e0da",
X"34831433",
X"83e0db34",
X"845283e0",
X"d851fea7",
X"3f83e080",
X"0881ff06",
X"84153355",
X"5372742e",
X"0981068c",
X"3892b73f",
X"83e08008",
X"802e9a38",
X"83e2f408",
X"a82e0981",
X"06893886",
X"0b83e2f4",
X"0c8739a8",
X"0b83e2f4",
X"0c80e451",
X"e2923f85",
X"3d0d04f4",
X"3d0d7e60",
X"5a55805d",
X"8075822b",
X"7183e2f8",
X"120c83e3",
X"8c175c5c",
X"56757a34",
X"78762e83",
X"ce387552",
X"78519c98",
X"3f8e3dfc",
X"05549053",
X"83e2e052",
X"78519bdb",
X"3f7c5877",
X"902e0981",
X"0683ac38",
X"83e2e051",
X"fd843f83",
X"e2e251fc",
X"fd3f83e2",
X"e451fcf6",
X"3f7583e2",
X"f00c7851",
X"99a73f80",
X"fbd45283",
X"e0800851",
X"f59e3f83",
X"e0800881",
X"2e098106",
X"80e33875",
X"83e3880c",
X"820b83e2",
X"e034ff96",
X"0b83e2e1",
X"3478519b",
X"d93f83e0",
X"80085583",
X"e0800876",
X"25883883",
X"e080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583e2e2",
X"347483e2",
X"e334800b",
X"83e2e434",
X"ff800b83",
X"e2e53478",
X"519bac3f",
X"83e2ef33",
X"83e08008",
X"0755819f",
X"3983e2e0",
X"3383e2e1",
X"3371882b",
X"07565c74",
X"83ffff2e",
X"09810680",
X"e838fe80",
X"0b83e388",
X"0c810b83",
X"e2f00cff",
X"0b83e2e0",
X"34ff0b83",
X"e2e13478",
X"519ad73f",
X"83e08008",
X"83e3900c",
X"83e08008",
X"5583e080",
X"08802588",
X"3883e080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"e2e23474",
X"83e2e334",
X"800b83e2",
X"e434ff80",
X"0b83e2e5",
X"34810b83",
X"e2ef34a4",
X"39748596",
X"2e098106",
X"81893877",
X"83e3880c",
X"78519a8b",
X"3f83e2ef",
X"3383e080",
X"08075574",
X"83e2ef34",
X"83e2ef33",
X"81065574",
X"802e8a38",
X"76840770",
X"81ff0658",
X"5583e2e4",
X"3383e2e5",
X"3371882b",
X"07565674",
X"81802e09",
X"8106a138",
X"83e2e233",
X"83e2e333",
X"71882b07",
X"565cad80",
X"75278738",
X"76820755",
X"94397681",
X"07558e39",
X"7482802e",
X"0981068c",
X"38768307",
X"557481ff",
X"06578739",
X"7481ff26",
X"8a387883",
X"e2f81c0c",
X"767a348e",
X"3d0d04fe",
X"3d0d800b",
X"83e2dc0c",
X"800b83e2",
X"d80cff0b",
X"83e0d40c",
X"a80b83e2",
X"f40cae51",
X"8cb43f80",
X"0b83e2f8",
X"54528073",
X"70840555",
X"0c811252",
X"71842e09",
X"8106ef38",
X"843d0d04",
X"fe3d0d74",
X"02840596",
X"05225353",
X"71802e96",
X"38727081",
X"05543351",
X"8cd33fff",
X"127083ff",
X"ff065152",
X"e739843d",
X"0d04fe3d",
X"0d029205",
X"225382ac",
X"51dda53f",
X"80c3518c",
X"b03f8196",
X"51dd993f",
X"725283e0",
X"d851ffb4",
X"3f725283",
X"e0d851f8",
X"de3f83e0",
X"800881ff",
X"06518c8d",
X"3f843d0d",
X"04ffb13d",
X"0d80d13d",
X"f80551f9",
X"883f83e2",
X"dc088105",
X"83e2dc0c",
X"80cf3d33",
X"cf117081",
X"ff065156",
X"56748326",
X"88dc3875",
X"8f06ff05",
X"567583e0",
X"d4082e9b",
X"38758326",
X"96387583",
X"e0d40c75",
X"842983e2",
X"f8057008",
X"53557551",
X"fa993f80",
X"762488b8",
X"38758429",
X"83e2f805",
X"55740880",
X"2e88a938",
X"83e0d408",
X"842983e2",
X"f8057008",
X"02880582",
X"b9053352",
X"5b557480",
X"d22e84a4",
X"387480d2",
X"24903874",
X"bf2e9c38",
X"7480d02e",
X"81d63887",
X"e8397480",
X"d32e80d4",
X"387480d7",
X"2e81c538",
X"87d73902",
X"82bb0533",
X"70882b81",
X"fe800602",
X"880582ba",
X"05337105",
X"5156568b",
X"8a3f80c1",
X"518abe3f",
X"f6d53f86",
X"0b83e0d8",
X"34815283",
X"e0d8518b",
X"f93f8151",
X"fde43f74",
X"8938860b",
X"83e2f40c",
X"8739a80b",
X"83e2f40c",
X"8ad93f80",
X"c1518a8d",
X"3ff6a43f",
X"900b83e2",
X"ef338106",
X"56567480",
X"2e833898",
X"5683e2e4",
X"3383e2e5",
X"3371882b",
X"07565974",
X"81802e09",
X"81069c38",
X"83e2e233",
X"83e2e333",
X"71882b07",
X"5657ad80",
X"75278c38",
X"75818007",
X"56853975",
X"a0075675",
X"83e0d834",
X"ff0b83e0",
X"d934e00b",
X"83e0da34",
X"800b83e0",
X"db348452",
X"83e0d851",
X"8af03f84",
X"51869039",
X"0282bb05",
X"3370882b",
X"81fe8006",
X"02880582",
X"ba053371",
X"05515659",
X"89c93f79",
X"5194dc3f",
X"83e08008",
X"802e8a38",
X"80ce5188",
X"f03f85e2",
X"3980c151",
X"88e73f89",
X"ef3f87f3",
X"3f83e388",
X"08588375",
X"259b3883",
X"e2e43383",
X"e2e53371",
X"882b07fc",
X"1771297a",
X"05838005",
X"5a51578d",
X"39748180",
X"2918ff80",
X"05588180",
X"57805676",
X"762e9238",
X"88c63f83",
X"e0800883",
X"e0d81734",
X"811656eb",
X"3988b53f",
X"83e08008",
X"81ff0677",
X"5383e0d8",
X"5256f4cb",
X"3f83e080",
X"0881ff06",
X"5575752e",
X"09810681",
X"843888b7",
X"3f80c151",
X"87eb3f88",
X"f33f7752",
X"79519384",
X"3f805e80",
X"d13dfdf4",
X"05547653",
X"83e0d852",
X"79519198",
X"3f0282b9",
X"05335581",
X"587480d7",
X"2e098106",
X"bc3880d1",
X"3dfdf005",
X"5476538f",
X"3d70537a",
X"5259929f",
X"3f805676",
X"762ea238",
X"751983e0",
X"d8173371",
X"33707232",
X"70307080",
X"2570307e",
X"06811d5d",
X"5e515151",
X"525b55db",
X"3982ac51",
X"d7ea3f77",
X"802e8638",
X"80c35184",
X"3980ce51",
X"86eb3f87",
X"f33f85f7",
X"3f83da39",
X"0282bb05",
X"3370882b",
X"81fe8006",
X"02880582",
X"ba053359",
X"78055956",
X"80705d59",
X"87893f80",
X"c15186bd",
X"3f83e2f0",
X"08792e82",
X"db3883e3",
X"900880fc",
X"055580fd",
X"527451bb",
X"ab3f83e0",
X"80085b77",
X"8224b238",
X"ff187087",
X"2b83ffff",
X"800680fd",
X"d40583e0",
X"d8595755",
X"81805575",
X"70810557",
X"33777081",
X"055934ff",
X"157081ff",
X"06515574",
X"ea38828a",
X"397782e8",
X"2e81aa38",
X"7782e92e",
X"09810681",
X"b13880fc",
X"8c518cd4",
X"3f785877",
X"87327030",
X"70720780",
X"257a8a32",
X"70307072",
X"07802573",
X"0753545a",
X"51575575",
X"802e9738",
X"78782692",
X"38a00b83",
X"e0d81a34",
X"81197081",
X"ff065a55",
X"eb398118",
X"7081ff06",
X"59558a78",
X"27ffbc38",
X"8f5883e0",
X"d3183383",
X"e0d81934",
X"ff187081",
X"ff065955",
X"778426ea",
X"38905880",
X"0b83e0d8",
X"19348118",
X"7081ff06",
X"70982b52",
X"59557480",
X"25e93880",
X"c6557a85",
X"8f248438",
X"80c25574",
X"83e0d834",
X"80f10b83",
X"e0db3481",
X"0b83e0dc",
X"347a83e0",
X"d9347a88",
X"2c557483",
X"e0da3480",
X"c93982f0",
X"782580c2",
X"387780fd",
X"29fd97d3",
X"05527951",
X"8fb63f80",
X"d13dfdec",
X"055480fd",
X"5383e0d8",
X"5279518e",
X"f63f7b81",
X"19595675",
X"80fc2483",
X"38785877",
X"882c5574",
X"83e1d534",
X"7783e1d6",
X"347583e1",
X"d7348180",
X"5980ca39",
X"83e38808",
X"57837825",
X"9b3883e2",
X"e43383e2",
X"e5337188",
X"2b07fc1a",
X"71297905",
X"83800559",
X"51598d39",
X"77818029",
X"17ff8005",
X"57818059",
X"76527951",
X"8ec63f80",
X"d13dfdec",
X"05547853",
X"83e0d852",
X"79518e87",
X"3f7851f6",
X"c93f8494",
X"3f82983f",
X"8b3983e2",
X"d8088105",
X"83e2d80c",
X"80d13d0d",
X"04f6ea3f",
X"dda13ff9",
X"39fc3d0d",
X"76787184",
X"2983e2f8",
X"05700851",
X"53535370",
X"9e3880ce",
X"723480cf",
X"0b811334",
X"80ce0b82",
X"133480c5",
X"0b831334",
X"70841334",
X"80e73983",
X"e38c1333",
X"5480d272",
X"3473822a",
X"70810651",
X"5180cf53",
X"70843880",
X"d7537281",
X"1334a00b",
X"82133473",
X"83065170",
X"812e9e38",
X"70812488",
X"3870802e",
X"8f389f39",
X"70822e92",
X"3870832e",
X"92389339",
X"80d8558e",
X"3980d355",
X"893980cd",
X"55843980",
X"c4557483",
X"133480c4",
X"0b841334",
X"800b8513",
X"34863d0d",
X"04fe3d0d",
X"80fcec08",
X"70337081",
X"ff067084",
X"2a813281",
X"06555152",
X"5371802e",
X"8c38a873",
X"3480fcec",
X"0851b871",
X"347183e0",
X"800c843d",
X"0d04fe3d",
X"0d80fcec",
X"08703370",
X"81ff0670",
X"852a8132",
X"81065551",
X"52537180",
X"2e8c3898",
X"733480fc",
X"ec0851b8",
X"71347183",
X"e0800c84",
X"3d0d0480",
X"3d0d80fc",
X"e8085193",
X"713480fc",
X"f40851ff",
X"7134823d",
X"0d04fe3d",
X"0d029305",
X"3380fce8",
X"08535380",
X"72348a51",
X"d1b23fd3",
X"3f80fcf8",
X"085280f8",
X"723480fd",
X"90085280",
X"7234fa13",
X"80fd9808",
X"53537272",
X"3480fd80",
X"08528072",
X"3480fd88",
X"08527272",
X"3480fcec",
X"08528072",
X"3480fcec",
X"0852b872",
X"34843d0d",
X"04ff3d0d",
X"028f0533",
X"80fcf008",
X"52527171",
X"34fe9e3f",
X"83e08008",
X"802ef638",
X"833d0d04",
X"803d0d84",
X"39da8c3f",
X"feb83f83",
X"e0800880",
X"2ef33880",
X"fcf00870",
X"337081ff",
X"0683e080",
X"0c515182",
X"3d0d0480",
X"3d0d80fc",
X"e80851a3",
X"713480fc",
X"f40851ff",
X"713480fc",
X"ec0851a8",
X"713480fc",
X"ec0851b8",
X"7134823d",
X"0d04803d",
X"0d80fce8",
X"08703370",
X"81c00670",
X"30708025",
X"83e0800c",
X"51515151",
X"823d0d04",
X"ff3d0d80",
X"fcec0870",
X"337081ff",
X"0670832a",
X"81327081",
X"06515151",
X"52527080",
X"2ee538b0",
X"723480fc",
X"ec0851b8",
X"7134833d",
X"0d04803d",
X"0d80fda4",
X"08700881",
X"0683e080",
X"0c51823d",
X"0d04fd3d",
X"0d757754",
X"54807325",
X"94387370",
X"81055533",
X"5280fc94",
X"51859d3f",
X"ff1353e9",
X"39853d0d",
X"04f63d0d",
X"7c7e6062",
X"5a5d5b56",
X"80598155",
X"8539747a",
X"29557452",
X"7551b2fc",
X"3f83e080",
X"087a27ee",
X"3874802e",
X"80dd3874",
X"527551b2",
X"e73f83e0",
X"80087553",
X"765254b3",
X"8e3f83e0",
X"80087a53",
X"755256b2",
X"cf3f83e0",
X"80087930",
X"707b079f",
X"2a707780",
X"24075151",
X"54557287",
X"3883e080",
X"08c53876",
X"8118b016",
X"55585889",
X"74258b38",
X"b714537a",
X"853880d7",
X"14537278",
X"34811959",
X"ff9f3980",
X"77348c3d",
X"0d04f73d",
X"0d7b7d7f",
X"62029005",
X"bb053357",
X"59565a5a",
X"b0587283",
X"38a05875",
X"70708105",
X"52337159",
X"54559039",
X"8074258e",
X"38ff1477",
X"70810559",
X"33545472",
X"ef3873ff",
X"15555380",
X"73258938",
X"77527951",
X"782def39",
X"75337557",
X"5372802e",
X"90387252",
X"7951782d",
X"75708105",
X"573353ed",
X"398b3d0d",
X"04ee3d0d",
X"64666969",
X"70708105",
X"52335b4a",
X"5c5e5e76",
X"802e82f9",
X"3876a52e",
X"09810682",
X"e0388070",
X"41677070",
X"81055233",
X"714a5957",
X"5f76b02e",
X"0981068c",
X"38757081",
X"05573376",
X"4857815f",
X"d0175675",
X"892680da",
X"3876675c",
X"59805c93",
X"39778a24",
X"80c3387b",
X"8a29187b",
X"7081055d",
X"335a5cd0",
X"197081ff",
X"06585889",
X"7727a438",
X"ff9f1970",
X"81ff06ff",
X"a91b5a51",
X"56857627",
X"9238ffbf",
X"197081ff",
X"06515675",
X"85268a38",
X"c9195877",
X"8025ffb9",
X"387a477b",
X"407881ff",
X"06577680",
X"e42e80e5",
X"387680e4",
X"24a73876",
X"80d82e81",
X"86387680",
X"d8249038",
X"76802e81",
X"cc3876a5",
X"2e81b638",
X"81b93976",
X"80e32e81",
X"8c3881af",
X"397680f5",
X"2e9b3876",
X"80f5248b",
X"387680f3",
X"2e818138",
X"81993976",
X"80f82e80",
X"ca38818f",
X"39913d70",
X"55578053",
X"8a527984",
X"1b710853",
X"5b56fc81",
X"3f7655ab",
X"3979841b",
X"7108943d",
X"705b5b52",
X"5b567580",
X"258c3875",
X"3056ad78",
X"340280c1",
X"05577654",
X"80538a52",
X"7551fbd5",
X"3f77557e",
X"54b83991",
X"3d705577",
X"80d83270",
X"30708025",
X"56515856",
X"90527984",
X"1b710853",
X"5b57fbb1",
X"3f7555db",
X"3979841b",
X"83123354",
X"5b569839",
X"79841b71",
X"08575b56",
X"80547f53",
X"7c527d51",
X"fc9c3f87",
X"3976527d",
X"517c2d66",
X"70335881",
X"0547fd83",
X"39943d0d",
X"047283e0",
X"900c7183",
X"e0940c04",
X"fb3d0d88",
X"3d707084",
X"05520857",
X"54755383",
X"e0900852",
X"83e09408",
X"51fcc63f",
X"873d0d04",
X"ff3d0d73",
X"70085351",
X"02930533",
X"72347008",
X"8105710c",
X"833d0d04",
X"fc3d0d87",
X"3d881155",
X"785480c2",
X"b45351fc",
X"983f8052",
X"873d51d0",
X"3f863d0d",
X"04803d0d",
X"72517080",
X"2e833881",
X"517083e0",
X"800c823d",
X"0d04ff3d",
X"0d028f05",
X"33703070",
X"9f2a83e0",
X"800c5252",
X"833d0d04",
X"fd3d0d75",
X"705254a4",
X"e73f83e0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83e0",
X"8008732e",
X"a13883e0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183e0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83e5b808",
X"248a38a5",
X"cf3fff0b",
X"83e5b80c",
X"800b83e0",
X"800c04ff",
X"3d0d7352",
X"83e39408",
X"722e8d38",
X"d93f7151",
X"96de3f71",
X"83e3940c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"558154bc",
X"15088192",
X"387451cf",
X"3f795880",
X"7a2580f7",
X"3883e5e8",
X"0870892a",
X"5783ff06",
X"78848072",
X"31565657",
X"73782583",
X"38735575",
X"83e5b808",
X"2e8438ff",
X"893f83e5",
X"b8088025",
X"a6387589",
X"2b5199ca",
X"3f83e5e8",
X"088f3dfc",
X"11555c54",
X"8152f81b",
X"5197af3f",
X"761483e5",
X"e80c7583",
X"e5b80c74",
X"53765278",
X"51a4803f",
X"83e08008",
X"83e5e808",
X"1683e5e8",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8b3861",
X"7a710c54",
X"7551fcf1",
X"3f83e080",
X"08547383",
X"e0800c8e",
X"3d0d04fc",
X"3d0dfe9a",
X"3f7651fe",
X"ae3f863d",
X"fc055302",
X"a2052252",
X"775196ce",
X"3f79863d",
X"22710c54",
X"83e08008",
X"51fcba3f",
X"863d0d04",
X"fd3d0d76",
X"83e5b808",
X"53538072",
X"24893871",
X"732e8438",
X"fddc3f75",
X"51fdf03f",
X"725198a2",
X"3f7351fc",
X"903f853d",
X"0d04803d",
X"0d7280c0",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d72bc",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"c40b83e0",
X"800c04fd",
X"3d0d7577",
X"71547053",
X"5553a0d4",
X"3f82c813",
X"08bc150c",
X"82c01308",
X"80c0150c",
X"fd803f73",
X"5194853f",
X"7383e394",
X"0c83e080",
X"0851fbb1",
X"3f853d0d",
X"04fd3d0d",
X"75775553",
X"fce03f72",
X"802ea538",
X"bc130852",
X"73519fea",
X"3f83e080",
X"088f3877",
X"527251ff",
X"a63f83e0",
X"8008538a",
X"3982cc13",
X"0853d839",
X"81537283",
X"e0800c85",
X"3d0d04ff",
X"3d0dff0b",
X"83e5b80c",
X"7383e398",
X"0c7483e5",
X"b40ca0d7",
X"3f83e080",
X"0881ff06",
X"5271802e",
X"88387151",
X"fadc3f90",
X"3983e5d0",
X"518f823f",
X"83e08008",
X"51fab63f",
X"833d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"519de23f",
X"83e08008",
X"557483e0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"e0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283e5b4",
X"0851a684",
X"3f83e080",
X"0857fa8a",
X"3f795283",
X"e5bc5196",
X"c73f83e0",
X"80085380",
X"5483e080",
X"08742e09",
X"81068283",
X"3883e398",
X"080b0b80",
X"fbc85370",
X"52559da0",
X"3f0b0b80",
X"fbc85280",
X"c015519d",
X"933f74bc",
X"160c7282",
X"c0160c81",
X"0b82c416",
X"0c810b82",
X"c8160cff",
X"17735757",
X"81973983",
X"e3a43370",
X"822a7081",
X"06515454",
X"72818638",
X"73812a81",
X"06587780",
X"fc387680",
X"2e819038",
X"82d015ff",
X"1875842a",
X"810682c4",
X"130c83e3",
X"a4338106",
X"82c8130c",
X"7b547153",
X"58569cb4",
X"3f75519c",
X"cb3f83e0",
X"80081653",
X"af737081",
X"05553472",
X"bc170c83",
X"e3a55272",
X"519c953f",
X"83e39c08",
X"82c0170c",
X"83e3b252",
X"83901551",
X"9c823f77",
X"82cc170c",
X"78802e8d",
X"38755178",
X"2d83e080",
X"08802e8d",
X"3874802e",
X"86387582",
X"cc160c75",
X"5583e39c",
X"5283e5bc",
X"5195e73f",
X"83e08008",
X"8a3883e3",
X"a5335372",
X"fed13880",
X"0b82cc17",
X"0c78802e",
X"893883e3",
X"980851fc",
X"b93f83e3",
X"98085473",
X"83e0800c",
X"8b3d0d04",
X"ff3d0d80",
X"527351fd",
X"b63f833d",
X"0d04f03d",
X"0d627052",
X"54f6b93f",
X"83e08008",
X"7453873d",
X"70535555",
X"f6d93ff7",
X"b93f7351",
X"d33f6353",
X"745283e0",
X"800851fa",
X"c03f923d",
X"0d047183",
X"e0800c04",
X"80c01283",
X"e0800c04",
X"803d0d72",
X"82c01108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"7282cc11",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282c4",
X"110883e0",
X"800c5182",
X"3d0d04f6",
X"3d0d7c83",
X"e0980859",
X"59817927",
X"82a93878",
X"88190827",
X"82a13877",
X"33567582",
X"2e819b38",
X"75822489",
X"3875812e",
X"8d38828b",
X"3975832e",
X"81b73882",
X"82397883",
X"ffff0670",
X"812a1170",
X"83ffff06",
X"7083ff06",
X"71892a90",
X"3d5f525a",
X"51515576",
X"83ff2e8e",
X"38825476",
X"538c1808",
X"15527951",
X"a9397554",
X"76538c18",
X"08155279",
X"519ad63f",
X"83e08008",
X"81bd3875",
X"5483e080",
X"08538c18",
X"08158105",
X"528c3dfd",
X"05519ab9",
X"3f83e080",
X"0881a038",
X"02a90533",
X"8c3d3371",
X"882b077a",
X"81067184",
X"2a535758",
X"56748638",
X"769fff06",
X"56755581",
X"80397554",
X"781083fe",
X"06537888",
X"2a8c1908",
X"05528c3d",
X"fc055199",
X"f83f83e0",
X"800880df",
X"3802a905",
X"338c3d33",
X"71882b07",
X"565780d1",
X"39845478",
X"822b83fc",
X"06537887",
X"2a8c1908",
X"05528c3d",
X"fc055199",
X"c83f83e0",
X"8008b038",
X"02ab0533",
X"028405aa",
X"05337198",
X"2b71902b",
X"07028c05",
X"a9053370",
X"882b7207",
X"903d3371",
X"80fffffe",
X"80060751",
X"52535758",
X"56833981",
X"557483e0",
X"800c8c3d",
X"0d04fb3d",
X"0d83e098",
X"08fe1988",
X"1208fe05",
X"55565480",
X"56747327",
X"8d388214",
X"33757129",
X"94160805",
X"57537583",
X"e0800c87",
X"3d0d04fc",
X"3d0d7683",
X"e0980855",
X"55807523",
X"88150853",
X"72812e88",
X"38881408",
X"73268538",
X"8152b239",
X"72903873",
X"33527183",
X"2e098106",
X"85389014",
X"0853728c",
X"160c7280",
X"2e8d3872",
X"51ff933f",
X"83e08008",
X"52853990",
X"14085271",
X"90160c80",
X"527183e0",
X"800c863d",
X"0d04fa3d",
X"0d7883e0",
X"98087122",
X"81057083",
X"ffff0657",
X"54575573",
X"802e8838",
X"90150853",
X"72863883",
X"5280e739",
X"738f0652",
X"7180da38",
X"81139016",
X"0c8c1508",
X"53729038",
X"830b8417",
X"22575273",
X"762780c6",
X"38bf3982",
X"1633ff05",
X"74842a06",
X"5271b238",
X"7251fbdb",
X"3f815271",
X"83e08008",
X"27a83883",
X"5283e080",
X"08881708",
X"279c3883",
X"e080088c",
X"160c83e0",
X"800851fd",
X"f93f83e0",
X"80089016",
X"0c737523",
X"80527183",
X"e0800c88",
X"3d0d04f2",
X"3d0d6062",
X"64585d5b",
X"75335574",
X"a02e0981",
X"06883881",
X"16704456",
X"ef396270",
X"33565674",
X"af2e0981",
X"06843881",
X"1643800b",
X"881c0c62",
X"70335155",
X"74a02691",
X"387a51fd",
X"d23f83e0",
X"80085680",
X"7c3483a8",
X"39933d84",
X"1c087058",
X"5a5f8a55",
X"a0767081",
X"055834ff",
X"155574ff",
X"2e098106",
X"ef388070",
X"595d887f",
X"085f5a7c",
X"811e7081",
X"ff066013",
X"703370af",
X"327030a0",
X"73277180",
X"25075151",
X"525b535f",
X"57557480",
X"d83876ae",
X"2e098106",
X"83388155",
X"777a2775",
X"07557480",
X"2e9f3879",
X"88327030",
X"78ae3270",
X"30707307",
X"9f2a5351",
X"57515675",
X"ac388858",
X"8b5affab",
X"39ff9f17",
X"55749926",
X"8938e017",
X"7081ff06",
X"58557781",
X"197081ff",
X"06721c53",
X"5a575576",
X"7534ff87",
X"397c1e7f",
X"0c805576",
X"a0268338",
X"8155748b",
X"1a347a51",
X"fc913f83",
X"e0800880",
X"f538a054",
X"7a227085",
X"2b83e006",
X"5455901b",
X"08527b51",
X"94cf3f83",
X"e0800857",
X"83e08008",
X"8182387b",
X"33557480",
X"2e80f538",
X"8b1c3370",
X"832a7081",
X"06515656",
X"74b4388b",
X"7c841d08",
X"83e08008",
X"595b5b58",
X"ff185877",
X"ff2e9a38",
X"79708105",
X"5b337970",
X"81055b33",
X"71713152",
X"56567580",
X"2ee23886",
X"3975802e",
X"bc387a51",
X"fbf43fff",
X"863983e0",
X"80085683",
X"e0800880",
X"2ea93883",
X"e0800883",
X"2e098106",
X"80de3884",
X"1b088b11",
X"33515574",
X"80d23884",
X"5680cd39",
X"8356ec39",
X"815680c4",
X"39765684",
X"1b088b11",
X"33515574",
X"b7388b1c",
X"3370842a",
X"70810651",
X"56577480",
X"2ed53895",
X"1c33941d",
X"3371982b",
X"71902b07",
X"9b1f337f",
X"9a053371",
X"882b0772",
X"077f8805",
X"0c5a5856",
X"58fcda39",
X"7583e080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"5192de3f",
X"835683e0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"5192b23f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"76519289",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583e080",
X"0c8a3d0d",
X"04ec3d0d",
X"6659800b",
X"83e0980c",
X"78567880",
X"2e83e838",
X"91a53f83",
X"e0800881",
X"06558256",
X"7483d838",
X"7475538e",
X"3d705358",
X"58fec23f",
X"83e08008",
X"81ff0656",
X"75812e09",
X"810680d4",
X"38905483",
X"be537452",
X"76519195",
X"3f83e080",
X"0880c938",
X"8e3d3355",
X"74802e80",
X"c93802bb",
X"05330284",
X"05ba0533",
X"71982b71",
X"902b0702",
X"8c05b905",
X"3370882b",
X"7207943d",
X"33710770",
X"587c5754",
X"525d5759",
X"56fde63f",
X"83e08008",
X"81ff0656",
X"75832e09",
X"81068638",
X"815682db",
X"3975802e",
X"86388756",
X"82d139a4",
X"548d5377",
X"52765190",
X"ac3f8156",
X"83e08008",
X"82bd3802",
X"ba053302",
X"8405b905",
X"3371882b",
X"07585c76",
X"ab380280",
X"ca053302",
X"840580c9",
X"05337198",
X"2b71902b",
X"07963d33",
X"70882b72",
X"07029405",
X"80c70533",
X"71075452",
X"5d575856",
X"02b30533",
X"77712902",
X"8805b205",
X"33028c05",
X"b1053371",
X"882b0770",
X"1c708c1f",
X"0c5e5957",
X"585c8d3d",
X"33821a34",
X"02b50533",
X"8f3d3371",
X"882b0759",
X"5b77841a",
X"2302b705",
X"33028405",
X"b6053371",
X"882b0756",
X"5b74ab38",
X"0280c605",
X"33028405",
X"80c50533",
X"71982b71",
X"902b0795",
X"3d337088",
X"2b720702",
X"940580c3",
X"05337107",
X"51525357",
X"5d5b7476",
X"31773178",
X"842a8f3d",
X"33547171",
X"31535656",
X"95e63f83",
X"e0800882",
X"0570881b",
X"0c709ff6",
X"26810557",
X"5583fff6",
X"75278338",
X"83567579",
X"3475832e",
X"098106af",
X"380280d2",
X"05330284",
X"0580d105",
X"3371982b",
X"71902b07",
X"983d3370",
X"882b7207",
X"02940580",
X"cf053371",
X"07901f0c",
X"525d5759",
X"56863976",
X"1a901a0c",
X"8419228c",
X"1a081871",
X"842a0594",
X"1b0c5c80",
X"0b811a34",
X"7883e098",
X"0c805675",
X"83e0800c",
X"963d0d04",
X"e93d0d83",
X"e0980856",
X"86547580",
X"2e81a638",
X"800b8117",
X"34993de0",
X"11466a54",
X"c01153ec",
X"0551f6cf",
X"3f83e080",
X"085483e0",
X"80088185",
X"38893d33",
X"5473802e",
X"933802ab",
X"05337084",
X"2a708106",
X"51555573",
X"802e8638",
X"835480e5",
X"3902b505",
X"338f3d33",
X"71982b71",
X"902b0702",
X"8c05bb05",
X"33029005",
X"ba053371",
X"882b0772",
X"07a01b0c",
X"029005bf",
X"05330294",
X"05be0533",
X"71982b71",
X"902b0702",
X"9c05bd05",
X"3370882b",
X"7207993d",
X"3371077f",
X"9c050c52",
X"83e08008",
X"981f0c56",
X"5a525253",
X"57595781",
X"0b811734",
X"83e08008",
X"547383e0",
X"800c993d",
X"0d04f53d",
X"0d7d6002",
X"8805ba05",
X"227283e0",
X"98085b5d",
X"5a5c5c80",
X"7b238656",
X"76802e81",
X"e0388117",
X"33810655",
X"85567480",
X"2e81d238",
X"9c170898",
X"18083155",
X"74782787",
X"387483ff",
X"ff065877",
X"802e81ae",
X"38981708",
X"7083ff06",
X"56567480",
X"ca388217",
X"33ff0576",
X"892a0670",
X"81ff065a",
X"5578a038",
X"758738a0",
X"1708558d",
X"39a41708",
X"51efe03f",
X"83e08008",
X"55817527",
X"80f83874",
X"a4180ca4",
X"170851f2",
X"8d3f83e0",
X"8008802e",
X"80e43883",
X"e0800819",
X"a8180c98",
X"170883ff",
X"06848071",
X"317083ff",
X"ff065851",
X"55777627",
X"83387756",
X"75549817",
X"0883ff06",
X"53a81708",
X"5279557b",
X"83387b55",
X"74518ad1",
X"3f83e080",
X"08a43898",
X"17081698",
X"180c751a",
X"78773170",
X"83ffff06",
X"7d227905",
X"525a565a",
X"747b23fe",
X"ce398056",
X"8839800b",
X"81183481",
X"567583e0",
X"800c8d3d",
X"0d04fa3d",
X"0d7883e0",
X"98085556",
X"86557380",
X"2e81dc38",
X"81143381",
X"06538555",
X"72802e81",
X"ce389c14",
X"08537276",
X"27833872",
X"56981408",
X"57800b98",
X"150c7580",
X"2e81a938",
X"82143370",
X"892b5653",
X"76802eb5",
X"387452ff",
X"165190d4",
X"3f83e080",
X"08ff1876",
X"54705358",
X"5390c53f",
X"83e08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b4387251",
X"edc13f83",
X"e0800853",
X"810b83e0",
X"80082780",
X"cb3883e0",
X"80088815",
X"082780c0",
X"3883e080",
X"08a4150c",
X"98140815",
X"98150c75",
X"753156c9",
X"39981408",
X"16709816",
X"0c735256",
X"efc83f83",
X"e0800880",
X"2e963882",
X"1433ff05",
X"76892a06",
X"83e08008",
X"05a8150c",
X"80558839",
X"800b8115",
X"34815574",
X"83e0800c",
X"883d0d04",
X"ee3d0d64",
X"56865583",
X"e0980880",
X"2e80f638",
X"943df411",
X"84180c66",
X"54d40552",
X"7551f197",
X"3f83e080",
X"085583e0",
X"800880cf",
X"38893d33",
X"5473802e",
X"bc3802ab",
X"05337084",
X"2a708106",
X"51555584",
X"5573802e",
X"bc3802b5",
X"05338f3d",
X"3371982b",
X"71902b07",
X"028c05bb",
X"05330290",
X"05ba0533",
X"71882b07",
X"7207881b",
X"0c535759",
X"577551ee",
X"d23f83e0",
X"80085574",
X"832e0981",
X"06833884",
X"557483e0",
X"800c943d",
X"0d04e43d",
X"0d6ea13d",
X"08405d86",
X"5683e098",
X"08802e84",
X"9b389e3d",
X"f405841e",
X"0c7e9838",
X"7c51ee97",
X"3f83e080",
X"08568484",
X"39814182",
X"80398341",
X"81fb3993",
X"3d7f9605",
X"4159807f",
X"8295055f",
X"56756081",
X"ff053483",
X"41901d08",
X"762e81dd",
X"38a0547c",
X"2270852b",
X"83e00654",
X"58901d08",
X"52785186",
X"ac3f83e0",
X"80084183",
X"e08008ff",
X"b8387833",
X"5c7b802e",
X"ffb4388b",
X"193370bf",
X"06718106",
X"52435574",
X"802e80e8",
X"387b81bf",
X"0655748f",
X"2480dd38",
X"9a193355",
X"7480d538",
X"9c193355",
X"74802e80",
X"cb38f31e",
X"70585e81",
X"56758b2e",
X"09810685",
X"388e568b",
X"39759a2e",
X"09810683",
X"389c5675",
X"19707081",
X"05523371",
X"33811a82",
X"1a5f5b52",
X"5b557486",
X"38797734",
X"853980df",
X"7734777b",
X"57577aa0",
X"2e098106",
X"c0388156",
X"7b81e532",
X"7030709f",
X"2a515155",
X"7bae2e93",
X"3874802e",
X"8e386183",
X"2a708106",
X"51557480",
X"2e97387c",
X"51ecf73f",
X"83e08008",
X"4183e080",
X"08873890",
X"1d08fea5",
X"38806034",
X"75802e88",
X"387d527f",
X"5183b13f",
X"60802e86",
X"38800b90",
X"1e0c6056",
X"60832e09",
X"81068838",
X"800b901e",
X"0c853960",
X"81d23889",
X"1f57901d",
X"08802e81",
X"a8388056",
X"75197033",
X"515574a0",
X"2ea03874",
X"852e0981",
X"06843881",
X"e5557477",
X"70810559",
X"34811670",
X"81ff0657",
X"55877627",
X"d7388819",
X"335574a0",
X"2ea938ae",
X"77708105",
X"59348856",
X"75197033",
X"515574a0",
X"2e953874",
X"77708105",
X"59348116",
X"7081ff06",
X"57558a76",
X"27e2388b",
X"19337f88",
X"05349f19",
X"339e1a33",
X"71982b71",
X"902b079d",
X"1c337088",
X"2b72079c",
X"1e337107",
X"640c5299",
X"1d33981e",
X"3371882b",
X"07535153",
X"57595674",
X"7f840523",
X"97193396",
X"1a337188",
X"2b075656",
X"747f8605",
X"23807734",
X"7c51eafe",
X"3f83e080",
X"085683e0",
X"8008832e",
X"09810688",
X"38800b90",
X"1e0c8056",
X"961f3355",
X"748a3889",
X"1f52961f",
X"5181b13f",
X"7583e080",
X"0c9e3d0d",
X"04fd3d0d",
X"75775354",
X"73335170",
X"89387133",
X"5170802e",
X"a1387333",
X"72335253",
X"72712785",
X"38ff5194",
X"39707327",
X"85388151",
X"8b398114",
X"81135354",
X"d3398051",
X"7083e080",
X"0c853d0d",
X"04fd3d0d",
X"75775454",
X"72337081",
X"ff065252",
X"70802ea3",
X"387181ff",
X"068114ff",
X"bf125354",
X"52709926",
X"8938a012",
X"7081ff06",
X"53517174",
X"70810556",
X"34d23980",
X"7434853d",
X"0d04ffbd",
X"3d0d80c6",
X"3d0852a5",
X"3d705254",
X"ffb33f80",
X"c73d0852",
X"853d7052",
X"53ffa63f",
X"72527351",
X"fedf3f80",
X"c53d0d04",
X"fe3d0d74",
X"76535371",
X"70810553",
X"33517073",
X"70810555",
X"3470f038",
X"843d0d04",
X"fe3d0d74",
X"52807233",
X"52537073",
X"2e8d3881",
X"12811471",
X"33535452",
X"70f53872",
X"83e0800c",
X"843d0d04",
X"fc3d0d76",
X"557483e5",
X"fc082eaf",
X"38805374",
X"5184cd3f",
X"83e08008",
X"81ff06ff",
X"147081ff",
X"06723070",
X"9f2a5152",
X"55535472",
X"802e8438",
X"71dd3873",
X"fe387483",
X"e5fc0c86",
X"3d0d0480",
X"3d0dff0b",
X"83e5fc0c",
X"82f63f85",
X"883f83e0",
X"800881ff",
X"065170f0",
X"3881d63f",
X"7083e080",
X"0c823d0d",
X"04fc3d0d",
X"76028405",
X"a2052202",
X"8805a605",
X"227a5455",
X"5555ff84",
X"3f72802e",
X"a03883e6",
X"8c143375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552dd",
X"39800b83",
X"e0800c86",
X"3d0d04fc",
X"3d0d7678",
X"7a115653",
X"55805371",
X"742e9338",
X"72155170",
X"3383e68c",
X"13348112",
X"81145452",
X"ea39800b",
X"83e0800c",
X"863d0d04",
X"fd3d0d90",
X"5483e5fc",
X"0851858a",
X"3f83e080",
X"0881ff06",
X"ff157130",
X"71307073",
X"079f2a72",
X"9f2a0652",
X"55525553",
X"72db3885",
X"3d0d04ff",
X"3d0d83e6",
X"88081083",
X"e6800807",
X"80fda808",
X"52710c83",
X"3d0d0480",
X"0b83e688",
X"0ce13f04",
X"810b83e6",
X"880cd83f",
X"04ed3f04",
X"7183e684",
X"0c04803d",
X"0d8051f4",
X"3f810b83",
X"e6880c81",
X"0b83e680",
X"0cffb83f",
X"823d0d04",
X"803d0d72",
X"30707407",
X"802583e6",
X"800c51ff",
X"a23f823d",
X"0d04fe3d",
X"0d029305",
X"3380fdac",
X"0854730c",
X"80fda808",
X"52710870",
X"81065151",
X"70f73872",
X"087081ff",
X"0683e080",
X"0c51843d",
X"0d04803d",
X"0d81ff51",
X"cd3f83e0",
X"800881ff",
X"0683e080",
X"0c823d0d",
X"04ff3d0d",
X"74902b74",
X"0780fd9c",
X"0852710c",
X"833d0d04",
X"803d0dfe",
X"f53f8051",
X"ff8a3f82",
X"3d0d04fe",
X"3d0d83e6",
X"8c0b8480",
X"115351d1",
X"3f843d0d",
X"04fd3d0d",
X"76028405",
X"97053353",
X"5381ff54",
X"ffa43fff",
X"a13fff9e",
X"3fff9b3f",
X"7180c007",
X"51fee73f",
X"72982a51",
X"fee03f72",
X"902a7081",
X"ff065252",
X"fed43f72",
X"882a7081",
X"ff065252",
X"fec83f72",
X"81ff0651",
X"fec03f81",
X"9551feba",
X"3ffee33f",
X"83e08008",
X"81ff06ff",
X"157081ff",
X"06703070",
X"9f2a5152",
X"56535372",
X"81ff2e09",
X"81068438",
X"71db3872",
X"83e0800c",
X"853d0d04",
X"fd3d0d81",
X"51fded3f",
X"75892b52",
X"9151fef1",
X"3f83e080",
X"0881ff06",
X"70555372",
X"a538fe96",
X"3f83e080",
X"0881ff06",
X"537281fe",
X"2e098106",
X"ed38febb",
X"3ffdff3f",
X"fdfc3f80",
X"51fdb53f",
X"80547383",
X"e0800c85",
X"3d0d04fe",
X"3d0d0293",
X"05335381",
X"51fd9d3f",
X"75527251",
X"fea33f83",
X"e0800881",
X"ff065380",
X"51fd893f",
X"7283e080",
X"0c843d0d",
X"04fd3d0d",
X"81ff53fd",
X"b93fff13",
X"7081ff06",
X"515372f3",
X"38725272",
X"51ffbc3f",
X"83e08008",
X"81ff0653",
X"81ff5472",
X"812e0981",
X"0680e238",
X"83ffff54",
X"8052b751",
X"ff9d3f83",
X"e0800881",
X"ff065372",
X"812e0981",
X"06a13880",
X"52a951ff",
X"863f83e0",
X"800881ff",
X"06537280",
X"2e8d38ff",
X"147083ff",
X"ff065553",
X"73ca3880",
X"528151fe",
X"e63f83e0",
X"800881ff",
X"065381ff",
X"54729238",
X"7252bb51",
X"fed13f84",
X"80529051",
X"fec93f72",
X"547383e0",
X"800c853d",
X"0d04fb3d",
X"0d83e68c",
X"568151fb",
X"db3f7789",
X"2b529851",
X"fcdf3f83",
X"e0800881",
X"ff067056",
X"547380d7",
X"38fc833f",
X"81fe51fb",
X"d13f8480",
X"53757081",
X"05573351",
X"fbc43fff",
X"137083ff",
X"ff065153",
X"72eb38fb",
X"e13ffbde",
X"3ffbdb3f",
X"83e08008",
X"81ff0670",
X"9f065455",
X"72852e09",
X"81069838",
X"fbc43f83",
X"e0800881",
X"ff065372",
X"802ef138",
X"8051faf0",
X"3f805574",
X"83e0800c",
X"873d0d04",
X"83e08c08",
X"0283e08c",
X"0cfd3d0d",
X"805383e0",
X"8c088c05",
X"085283e0",
X"8c088805",
X"085183d4",
X"3f83e080",
X"087083e0",
X"800c5485",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"fd3d0d81",
X"5383e08c",
X"088c0508",
X"5283e08c",
X"08880508",
X"5183a13f",
X"83e08008",
X"7083e080",
X"0c54853d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cf9",
X"3d0d800b",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"05088025",
X"b93883e0",
X"8c088805",
X"083083e0",
X"8c088805",
X"0c800b83",
X"e08c08f4",
X"050c83e0",
X"8c08fc05",
X"088a3881",
X"0b83e08c",
X"08f4050c",
X"83e08c08",
X"f4050883",
X"e08c08fc",
X"050c83e0",
X"8c088c05",
X"088025b9",
X"3883e08c",
X"088c0508",
X"3083e08c",
X"088c050c",
X"800b83e0",
X"8c08f005",
X"0c83e08c",
X"08fc0508",
X"8a38810b",
X"83e08c08",
X"f0050c83",
X"e08c08f0",
X"050883e0",
X"8c08fc05",
X"0c805383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"05085181",
X"df3f83e0",
X"80087083",
X"e08c08f8",
X"050c5483",
X"e08c08fc",
X"0508802e",
X"903883e0",
X"8c08f805",
X"083083e0",
X"8c08f805",
X"0c83e08c",
X"08f80508",
X"7083e080",
X"0c54893d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cfb",
X"3d0d800b",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"05088025",
X"993883e0",
X"8c088805",
X"083083e0",
X"8c088805",
X"0c810b83",
X"e08c08fc",
X"050c83e0",
X"8c088c05",
X"08802590",
X"3883e08c",
X"088c0508",
X"3083e08c",
X"088c050c",
X"815383e0",
X"8c088c05",
X"085283e0",
X"8c088805",
X"0851bd3f",
X"83e08008",
X"7083e08c",
X"08f8050c",
X"5483e08c",
X"08fc0508",
X"802e9038",
X"83e08c08",
X"f8050830",
X"83e08c08",
X"f8050c83",
X"e08c08f8",
X"05087083",
X"e0800c54",
X"873d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cfd3d0d",
X"810b83e0",
X"8c08fc05",
X"0c800b83",
X"e08c08f8",
X"050c83e0",
X"8c088c05",
X"0883e08c",
X"08880508",
X"27b93883",
X"e08c08fc",
X"0508802e",
X"ae38800b",
X"83e08c08",
X"8c050824",
X"a23883e0",
X"8c088c05",
X"081083e0",
X"8c088c05",
X"0c83e08c",
X"08fc0508",
X"1083e08c",
X"08fc050c",
X"ffb83983",
X"e08c08fc",
X"0508802e",
X"80e13883",
X"e08c088c",
X"050883e0",
X"8c088805",
X"0826ad38",
X"83e08c08",
X"88050883",
X"e08c088c",
X"05083183",
X"e08c0888",
X"050c83e0",
X"8c08f805",
X"0883e08c",
X"08fc0508",
X"0783e08c",
X"08f8050c",
X"83e08c08",
X"fc050881",
X"2a83e08c",
X"08fc050c",
X"83e08c08",
X"8c050881",
X"2a83e08c",
X"088c050c",
X"ff953983",
X"e08c0890",
X"0508802e",
X"933883e0",
X"8c088805",
X"087083e0",
X"8c08f405",
X"0c519139",
X"83e08c08",
X"f8050870",
X"83e08c08",
X"f4050c51",
X"83e08c08",
X"f4050883",
X"e0800c85",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"ff3d0d80",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"88050881",
X"06ff1170",
X"097083e0",
X"8c088c05",
X"080683e0",
X"8c08fc05",
X"081183e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"812a83e0",
X"8c088805",
X"0c83e08c",
X"088c0508",
X"1083e08c",
X"088c050c",
X"51515151",
X"83e08c08",
X"88050880",
X"2e8438ff",
X"ab3983e0",
X"8c08fc05",
X"087083e0",
X"800c5183",
X"3d0d83e0",
X"8c0c04fc",
X"3d0d7670",
X"797b5555",
X"55558f72",
X"278c3872",
X"75078306",
X"5170802e",
X"a938ff12",
X"5271ff2e",
X"98387270",
X"81055433",
X"74708105",
X"5634ff12",
X"5271ff2e",
X"098106ea",
X"387483e0",
X"800c863d",
X"0d047451",
X"72708405",
X"54087170",
X"8405530c",
X"72708405",
X"54087170",
X"8405530c",
X"72708405",
X"54087170",
X"8405530c",
X"72708405",
X"54087170",
X"8405530c",
X"f0125271",
X"8f26c938",
X"83722795",
X"38727084",
X"05540871",
X"70840553",
X"0cfc1252",
X"718326ed",
X"387054ff",
X"81390000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"000007ba",
X"000007c2",
X"000007ca",
X"000007d2",
X"000007da",
X"000007e2",
X"000007ea",
X"000007f2",
X"0000099c",
X"000009dd",
X"000009ff",
X"00000a21",
X"00000a21",
X"00000a21",
X"00000a21",
X"00000a7f",
X"00000aaf",
X"70704740",
X"9c704268",
X"9c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d20",
X"62616e6b",
X"3a256400",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"43617274",
X"72696467",
X"6520386b",
X"2073696d",
X"706c6500",
X"45786974",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"69383030",
X"00000000",
X"786c6f72",
X"69672e72",
X"6f6d0000",
X"786c6869",
X"61732e72",
X"6f6d0000",
X"756c7469",
X"6d6f6e2e",
X"726f6d00",
X"6f736268",
X"6961732e",
X"726f6d00",
X"6f73626f",
X"7269672e",
X"726f6d00",
X"6f73616f",
X"7269672e",
X"726f6d00",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"25732025",
X"73000000",
X"2e2e0000",
X"2f000000",
X"41545200",
X"58464400",
X"58455800",
X"524f4d00",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"6e616d65",
X"20000000",
X"25303278",
X"00000000",
X"00000000",
X"00000000",
X"0001d20f",
X"0001d400",
X"0001d401",
X"0001d409",
X"0001d010",
X"0001d301",
X"0001d300",
X"0001d20a",
X"0001d01b",
X"0001d016",
X"0001d019",
X"0001d018",
X"0001d017",
X"0001d01a",
X"0001d403",
X"0001d402",
X"0001d40e",
X"0004007c",
X"00040078",
X"00040074",
X"00040068",
X"00040060",
X"0004005c",
X"00040058",
X"00040054",
X"00040050",
X"0004004c",
X"00040048",
X"00040044",
X"00040040",
X"00040034",
X"00040030",
X"0004002c",
X"00040028",
X"00040024",
X"00040020",
X"0004001c",
X"00040018",
X"00040014",
X"00040010",
X"0004000c",
X"00040008",
X"00040004",
X"00040000",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
