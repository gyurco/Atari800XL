---------------------------------------------------------------------------
-- (c) 2013 mark watson
-- I am happy for anyone to use this for non-commercial use.
-- If my vhdl files are used commercially or otherwise sold,
-- please contact me for explicit permission at scrameta (gmail).
-- This applies for source and binary form and derived works.
---------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use IEEE.STD_LOGIC_MISC.all;

ENTITY pokey_mixer IS
PORT 
( 
	CHANNEL_0 : IN STD_LOGIC_VECTOR(3 downto 0);
	CHANNEL_1 : IN STD_LOGIC_VECTOR(3 downto 0);
	CHANNEL_2 : IN STD_LOGIC_VECTOR(3 downto 0);
	CHANNEL_3 : IN STD_LOGIC_VECTOR(3 downto 0);
	
	GTIA_SOUND : IN STD_LOGIC;

	COVOX_CHANNEL_0 : IN STD_LOGIC_VECTOR(7 downto 0);
	COVOX_CHANNEL_1 : IN STD_LOGIC_VECTOR(7 downto 0);
	
	VOLUME_OUT_NEXT : OUT STD_LOGIC_vector(15 downto 0)
);
END pokey_mixer;

ARCHITECTURE vhdl OF pokey_mixer IS
	signal volume_sum : std_logic_vector(9 downto 0);
	signal volume_next : std_logic_vector(15 downto 0);
BEGIN
	-- next state
	process (channel_0,channel_1,channel_2,channel_3,covox_CHANNEL_0,covox_channel_1,gtia_sound)
		variable channel0_en_long : unsigned(10 downto 0);
		variable channel1_en_long : unsigned(10 downto 0);
		variable channel2_en_long : unsigned(10 downto 0);
		variable channel3_en_long : unsigned(10 downto 0);
		variable gtia_sound_long : unsigned(10 downto 0);
		variable covox_0_long : unsigned(10 downto 0);
		variable covox_1_long : unsigned(10 downto 0);
		
		variable volume_int_sum : unsigned(10 downto 0);
	begin
		channel0_en_long := (others=>'0');
		channel1_en_long := (others=>'0');
		channel2_en_long := (others=>'0');
		channel3_en_long := (others=>'0');
		gtia_sound_long := (others=>'0');
		covox_0_long := (others=>'0');
		covox_1_long := (others=>'0');

		channel0_en_long(7 downto 4) := unsigned(channel_0);
		channel1_en_long(7 downto 4) := unsigned(channel_1);
		channel2_en_long(7 downto 4) := unsigned(channel_2);
		channel3_en_long(7 downto 4) := unsigned(channel_3);
		gtia_sound_long(7 downto 4) := gtia_sound&gtia_sound&gtia_sound&gtia_sound;
		covox_0_long(7 downto 0) := unsigned(covox_channel_0);
		covox_1_long(7 downto 0) := unsigned(covox_channel_1);

		volume_int_sum := ((channel0_en_long + channel1_en_long) + (channel2_en_long + channel3_en_long)) + (gtia_sound_long + (covox_0_long + covox_1_long));

		volume_sum(9 downto 0) <= std_logic_vector(volume_int_sum(9 downto 0)) or volume_int_sum(10)&volume_int_sum(10)&volume_int_sum(10)&volume_int_sum(10)&volume_int_sum(10)&volume_int_sum(10)&volume_int_sum(10)&volume_int_sum(10)&volume_int_sum(10)&volume_int_sum(10);
	end process;
	
 	process (volume_sum, volume_next)
	begin
		case volume_sum(9 downto 0) is 
			when "0000000000" =>
				volume_next <= X"8001";
			when "0000000001" =>
				volume_next <= X"80ce";
			when "0000000010" =>
				volume_next <= X"819a";
			when "0000000011" =>
				volume_next <= X"8266";
			when "0000000100" =>
				volume_next <= X"8331";
			when "0000000101" =>
				volume_next <= X"83fc";
			when "0000000110" =>
				volume_next <= X"84c6";
			when "0000000111" =>
				volume_next <= X"8590";
			when "0000001000" =>
				volume_next <= X"8659";
			when "0000001001" =>
				volume_next <= X"8722";
			when "0000001010" =>
				volume_next <= X"87ea";
			when "0000001011" =>
				volume_next <= X"88b2";
			when "0000001100" =>
				volume_next <= X"8979";
			when "0000001101" =>
				volume_next <= X"8a40";
			when "0000001110" =>
				volume_next <= X"8b07";
			when "0000001111" =>
				volume_next <= X"8bcd";
			when "0000010000" =>
				volume_next <= X"8c93";
			when "0000010001" =>
				volume_next <= X"8d58";
			when "0000010010" =>
				volume_next <= X"8e1c";
			when "0000010011" =>
				volume_next <= X"8ee1";
			when "0000010100" =>
				volume_next <= X"8fa4";
			when "0000010101" =>
				volume_next <= X"9068";
			when "0000010110" =>
				volume_next <= X"912a";
			when "0000010111" =>
				volume_next <= X"91ed";
			when "0000011000" =>
				volume_next <= X"92af";
			when "0000011001" =>
				volume_next <= X"9370";
			when "0000011010" =>
				volume_next <= X"9431";
			when "0000011011" =>
				volume_next <= X"94f2";
			when "0000011100" =>
				volume_next <= X"95b2";
			when "0000011101" =>
				volume_next <= X"9672";
			when "0000011110" =>
				volume_next <= X"9731";
			when "0000011111" =>
				volume_next <= X"97ef";
			when "0000100000" =>
				volume_next <= X"98ae";
			when "0000100001" =>
				volume_next <= X"996c";
			when "0000100010" =>
				volume_next <= X"9a29";
			when "0000100011" =>
				volume_next <= X"9ae6";
			when "0000100100" =>
				volume_next <= X"9ba2";
			when "0000100101" =>
				volume_next <= X"9c5e";
			when "0000100110" =>
				volume_next <= X"9d1a";
			when "0000100111" =>
				volume_next <= X"9dd5";
			when "0000101000" =>
				volume_next <= X"9e90";
			when "0000101001" =>
				volume_next <= X"9f4a";
			when "0000101010" =>
				volume_next <= X"a004";
			when "0000101011" =>
				volume_next <= X"a0bd";
			when "0000101100" =>
				volume_next <= X"a176";
			when "0000101101" =>
				volume_next <= X"a22f";
			when "0000101110" =>
				volume_next <= X"a2e7";
			when "0000101111" =>
				volume_next <= X"a39e";
			when "0000110000" =>
				volume_next <= X"a456";
			when "0000110001" =>
				volume_next <= X"a50c";
			when "0000110010" =>
				volume_next <= X"a5c3";
			when "0000110011" =>
				volume_next <= X"a678";
			when "0000110100" =>
				volume_next <= X"a72e";
			when "0000110101" =>
				volume_next <= X"a7e3";
			when "0000110110" =>
				volume_next <= X"a897";
			when "0000110111" =>
				volume_next <= X"a94b";
			when "0000111000" =>
				volume_next <= X"a9ff";
			when "0000111001" =>
				volume_next <= X"aab2";
			when "0000111010" =>
				volume_next <= X"ab65";
			when "0000111011" =>
				volume_next <= X"ac17";
			when "0000111100" =>
				volume_next <= X"acc9";
			when "0000111101" =>
				volume_next <= X"ad7b";
			when "0000111110" =>
				volume_next <= X"ae2c";
			when "0000111111" =>
				volume_next <= X"aedc";
			when "0001000000" =>
				volume_next <= X"af8c";
			when "0001000001" =>
				volume_next <= X"b03c";
			when "0001000010" =>
				volume_next <= X"b0eb";
			when "0001000011" =>
				volume_next <= X"b19a";
			when "0001000100" =>
				volume_next <= X"b249";
			when "0001000101" =>
				volume_next <= X"b2f7";
			when "0001000110" =>
				volume_next <= X"b3a4";
			when "0001000111" =>
				volume_next <= X"b451";
			when "0001001000" =>
				volume_next <= X"b4fe";
			when "0001001001" =>
				volume_next <= X"b5aa";
			when "0001001010" =>
				volume_next <= X"b656";
			when "0001001011" =>
				volume_next <= X"b702";
			when "0001001100" =>
				volume_next <= X"b7ad";
			when "0001001101" =>
				volume_next <= X"b857";
			when "0001001110" =>
				volume_next <= X"b901";
			when "0001001111" =>
				volume_next <= X"b9ab";
			when "0001010000" =>
				volume_next <= X"ba54";
			when "0001010001" =>
				volume_next <= X"bafd";
			when "0001010010" =>
				volume_next <= X"bba6";
			when "0001010011" =>
				volume_next <= X"bc4e";
			when "0001010100" =>
				volume_next <= X"bcf5";
			when "0001010101" =>
				volume_next <= X"bd9d";
			when "0001010110" =>
				volume_next <= X"be43";
			when "0001010111" =>
				volume_next <= X"beea";
			when "0001011000" =>
				volume_next <= X"bf90";
			when "0001011001" =>
				volume_next <= X"c035";
			when "0001011010" =>
				volume_next <= X"c0da";
			when "0001011011" =>
				volume_next <= X"c17f";
			when "0001011100" =>
				volume_next <= X"c223";
			when "0001011101" =>
				volume_next <= X"c2c7";
			when "0001011110" =>
				volume_next <= X"c36b";
			when "0001011111" =>
				volume_next <= X"c40e";
			when "0001100000" =>
				volume_next <= X"c4b0";
			when "0001100001" =>
				volume_next <= X"c552";
			when "0001100010" =>
				volume_next <= X"c5f4";
			when "0001100011" =>
				volume_next <= X"c696";
			when "0001100100" =>
				volume_next <= X"c737";
			when "0001100101" =>
				volume_next <= X"c7d7";
			when "0001100110" =>
				volume_next <= X"c877";
			when "0001100111" =>
				volume_next <= X"c917";
			when "0001101000" =>
				volume_next <= X"c9b6";
			when "0001101001" =>
				volume_next <= X"ca55";
			when "0001101010" =>
				volume_next <= X"caf4";
			when "0001101011" =>
				volume_next <= X"cb92";
			when "0001101100" =>
				volume_next <= X"cc2f";
			when "0001101101" =>
				volume_next <= X"cccd";
			when "0001101110" =>
				volume_next <= X"cd6a";
			when "0001101111" =>
				volume_next <= X"ce06";
			when "0001110000" =>
				volume_next <= X"cea2";
			when "0001110001" =>
				volume_next <= X"cf3e";
			when "0001110010" =>
				volume_next <= X"cfd9";
			when "0001110011" =>
				volume_next <= X"d074";
			when "0001110100" =>
				volume_next <= X"d10e";
			when "0001110101" =>
				volume_next <= X"d1a8";
			when "0001110110" =>
				volume_next <= X"d242";
			when "0001110111" =>
				volume_next <= X"d2db";
			when "0001111000" =>
				volume_next <= X"d374";
			when "0001111001" =>
				volume_next <= X"d40c";
			when "0001111010" =>
				volume_next <= X"d4a5";
			when "0001111011" =>
				volume_next <= X"d53c";
			when "0001111100" =>
				volume_next <= X"d5d3";
			when "0001111101" =>
				volume_next <= X"d66a";
			when "0001111110" =>
				volume_next <= X"d701";
			when "0001111111" =>
				volume_next <= X"d797";
			when "0010000000" =>
				volume_next <= X"d82c";
			when "0010000001" =>
				volume_next <= X"d8c2";
			when "0010000010" =>
				volume_next <= X"d956";
			when "0010000011" =>
				volume_next <= X"d9eb";
			when "0010000100" =>
				volume_next <= X"da7f";
			when "0010000101" =>
				volume_next <= X"db13";
			when "0010000110" =>
				volume_next <= X"dba6";
			when "0010000111" =>
				volume_next <= X"dc39";
			when "0010001000" =>
				volume_next <= X"dccb";
			when "0010001001" =>
				volume_next <= X"dd5e";
			when "0010001010" =>
				volume_next <= X"ddef";
			when "0010001011" =>
				volume_next <= X"de81";
			when "0010001100" =>
				volume_next <= X"df12";
			when "0010001101" =>
				volume_next <= X"dfa2";
			when "0010001110" =>
				volume_next <= X"e032";
			when "0010001111" =>
				volume_next <= X"e0c2";
			when "0010010000" =>
				volume_next <= X"e151";
			when "0010010001" =>
				volume_next <= X"e1e0";
			when "0010010010" =>
				volume_next <= X"e26f";
			when "0010010011" =>
				volume_next <= X"e2fd";
			when "0010010100" =>
				volume_next <= X"e38b";
			when "0010010101" =>
				volume_next <= X"e419";
			when "0010010110" =>
				volume_next <= X"e4a6";
			when "0010010111" =>
				volume_next <= X"e532";
			when "0010011000" =>
				volume_next <= X"e5bf";
			when "0010011001" =>
				volume_next <= X"e64b";
			when "0010011010" =>
				volume_next <= X"e6d6";
			when "0010011011" =>
				volume_next <= X"e761";
			when "0010011100" =>
				volume_next <= X"e7ec";
			when "0010011101" =>
				volume_next <= X"e877";
			when "0010011110" =>
				volume_next <= X"e901";
			when "0010011111" =>
				volume_next <= X"e98a";
			when "0010100000" =>
				volume_next <= X"ea14";
			when "0010100001" =>
				volume_next <= X"ea9d";
			when "0010100010" =>
				volume_next <= X"eb25";
			when "0010100011" =>
				volume_next <= X"ebad";
			when "0010100100" =>
				volume_next <= X"ec35";
			when "0010100101" =>
				volume_next <= X"ecbc";
			when "0010100110" =>
				volume_next <= X"ed43";
			when "0010100111" =>
				volume_next <= X"edca";
			when "0010101000" =>
				volume_next <= X"ee50";
			when "0010101001" =>
				volume_next <= X"eed6";
			when "0010101010" =>
				volume_next <= X"ef5c";
			when "0010101011" =>
				volume_next <= X"efe1";
			when "0010101100" =>
				volume_next <= X"f066";
			when "0010101101" =>
				volume_next <= X"f0ea";
			when "0010101110" =>
				volume_next <= X"f16e";
			when "0010101111" =>
				volume_next <= X"f1f2";
			when "0010110000" =>
				volume_next <= X"f275";
			when "0010110001" =>
				volume_next <= X"f2f8";
			when "0010110010" =>
				volume_next <= X"f37b";
			when "0010110011" =>
				volume_next <= X"f3fd";
			when "0010110100" =>
				volume_next <= X"f47f";
			when "0010110101" =>
				volume_next <= X"f500";
			when "0010110110" =>
				volume_next <= X"f582";
			when "0010110111" =>
				volume_next <= X"f602";
			when "0010111000" =>
				volume_next <= X"f683";
			when "0010111001" =>
				volume_next <= X"f703";
			when "0010111010" =>
				volume_next <= X"f782";
			when "0010111011" =>
				volume_next <= X"f802";
			when "0010111100" =>
				volume_next <= X"f881";
			when "0010111101" =>
				volume_next <= X"f8ff";
			when "0010111110" =>
				volume_next <= X"f97e";
			when "0010111111" =>
				volume_next <= X"f9fb";
			when "0011000000" =>
				volume_next <= X"fa79";
			when "0011000001" =>
				volume_next <= X"faf6";
			when "0011000010" =>
				volume_next <= X"fb73";
			when "0011000011" =>
				volume_next <= X"fbef";
			when "0011000100" =>
				volume_next <= X"fc6b";
			when "0011000101" =>
				volume_next <= X"fce7";
			when "0011000110" =>
				volume_next <= X"fd63";
			when "0011000111" =>
				volume_next <= X"fdde";
			when "0011001000" =>
				volume_next <= X"fe58";
			when "0011001001" =>
				volume_next <= X"fed3";
			when "0011001010" =>
				volume_next <= X"ff4c";
			when "0011001011" =>
				volume_next <= X"ffc6";
			when "0011001100" =>
				volume_next <= X"003e";
			when "0011001101" =>
				volume_next <= X"00b7";
			when "0011001110" =>
				volume_next <= X"0130";
			when "0011001111" =>
				volume_next <= X"01a8";
			when "0011010000" =>
				volume_next <= X"0220";
			when "0011010001" =>
				volume_next <= X"0297";
			when "0011010010" =>
				volume_next <= X"030e";
			when "0011010011" =>
				volume_next <= X"0385";
			when "0011010100" =>
				volume_next <= X"03fc";
			when "0011010101" =>
				volume_next <= X"0472";
			when "0011010110" =>
				volume_next <= X"04e8";
			when "0011010111" =>
				volume_next <= X"055d";
			when "0011011000" =>
				volume_next <= X"05d2";
			when "0011011001" =>
				volume_next <= X"0647";
			when "0011011010" =>
				volume_next <= X"06bb";
			when "0011011011" =>
				volume_next <= X"072f";
			when "0011011100" =>
				volume_next <= X"07a3";
			when "0011011101" =>
				volume_next <= X"0816";
			when "0011011110" =>
				volume_next <= X"0889";
			when "0011011111" =>
				volume_next <= X"08fc";
			when "0011100000" =>
				volume_next <= X"096e";
			when "0011100001" =>
				volume_next <= X"09e0";
			when "0011100010" =>
				volume_next <= X"0a52";
			when "0011100011" =>
				volume_next <= X"0ac3";
			when "0011100100" =>
				volume_next <= X"0b34";
			when "0011100101" =>
				volume_next <= X"0ba5";
			when "0011100110" =>
				volume_next <= X"0c15";
			when "0011100111" =>
				volume_next <= X"0c85";
			when "0011101000" =>
				volume_next <= X"0cf5";
			when "0011101001" =>
				volume_next <= X"0d64";
			when "0011101010" =>
				volume_next <= X"0dd3";
			when "0011101011" =>
				volume_next <= X"0e42";
			when "0011101100" =>
				volume_next <= X"0eb0";
			when "0011101101" =>
				volume_next <= X"0f1e";
			when "0011101110" =>
				volume_next <= X"0f8c";
			when "0011101111" =>
				volume_next <= X"0ff9";
			when "0011110000" =>
				volume_next <= X"1066";
			when "0011110001" =>
				volume_next <= X"10d2";
			when "0011110010" =>
				volume_next <= X"113f";
			when "0011110011" =>
				volume_next <= X"11ab";
			when "0011110100" =>
				volume_next <= X"1216";
			when "0011110101" =>
				volume_next <= X"1282";
			when "0011110110" =>
				volume_next <= X"12ed";
			when "0011110111" =>
				volume_next <= X"1357";
			when "0011111000" =>
				volume_next <= X"13c2";
			when "0011111001" =>
				volume_next <= X"142c";
			when "0011111010" =>
				volume_next <= X"1495";
			when "0011111011" =>
				volume_next <= X"14ff";
			when "0011111100" =>
				volume_next <= X"1568";
			when "0011111101" =>
				volume_next <= X"15d0";
			when "0011111110" =>
				volume_next <= X"1639";
			when "0011111111" =>
				volume_next <= X"16a1";
			when "0100000000" =>
				volume_next <= X"1709";
			when "0100000001" =>
				volume_next <= X"1770";
			when "0100000010" =>
				volume_next <= X"17d7";
			when "0100000011" =>
				volume_next <= X"183e";
			when "0100000100" =>
				volume_next <= X"18a4";
			when "0100000101" =>
				volume_next <= X"190a";
			when "0100000110" =>
				volume_next <= X"1970";
			when "0100000111" =>
				volume_next <= X"19d6";
			when "0100001000" =>
				volume_next <= X"1a3b";
			when "0100001001" =>
				volume_next <= X"1aa0";
			when "0100001010" =>
				volume_next <= X"1b04";
			when "0100001011" =>
				volume_next <= X"1b69";
			when "0100001100" =>
				volume_next <= X"1bcd";
			when "0100001101" =>
				volume_next <= X"1c30";
			when "0100001110" =>
				volume_next <= X"1c93";
			when "0100001111" =>
				volume_next <= X"1cf6";
			when "0100010000" =>
				volume_next <= X"1d59";
			when "0100010001" =>
				volume_next <= X"1dbb";
			when "0100010010" =>
				volume_next <= X"1e1e";
			when "0100010011" =>
				volume_next <= X"1e7f";
			when "0100010100" =>
				volume_next <= X"1ee1";
			when "0100010101" =>
				volume_next <= X"1f42";
			when "0100010110" =>
				volume_next <= X"1fa3";
			when "0100010111" =>
				volume_next <= X"2003";
			when "0100011000" =>
				volume_next <= X"2063";
			when "0100011001" =>
				volume_next <= X"20c3";
			when "0100011010" =>
				volume_next <= X"2123";
			when "0100011011" =>
				volume_next <= X"2182";
			when "0100011100" =>
				volume_next <= X"21e1";
			when "0100011101" =>
				volume_next <= X"2240";
			when "0100011110" =>
				volume_next <= X"229e";
			when "0100011111" =>
				volume_next <= X"22fc";
			when "0100100000" =>
				volume_next <= X"235a";
			when "0100100001" =>
				volume_next <= X"23b7";
			when "0100100010" =>
				volume_next <= X"2414";
			when "0100100011" =>
				volume_next <= X"2471";
			when "0100100100" =>
				volume_next <= X"24ce";
			when "0100100101" =>
				volume_next <= X"252a";
			when "0100100110" =>
				volume_next <= X"2586";
			when "0100100111" =>
				volume_next <= X"25e1";
			when "0100101000" =>
				volume_next <= X"263d";
			when "0100101001" =>
				volume_next <= X"2698";
			when "0100101010" =>
				volume_next <= X"26f3";
			when "0100101011" =>
				volume_next <= X"274d";
			when "0100101100" =>
				volume_next <= X"27a7";
			when "0100101101" =>
				volume_next <= X"2801";
			when "0100101110" =>
				volume_next <= X"285b";
			when "0100101111" =>
				volume_next <= X"28b4";
			when "0100110000" =>
				volume_next <= X"290d";
			when "0100110001" =>
				volume_next <= X"2965";
			when "0100110010" =>
				volume_next <= X"29be";
			when "0100110011" =>
				volume_next <= X"2a16";
			when "0100110100" =>
				volume_next <= X"2a6e";
			when "0100110101" =>
				volume_next <= X"2ac5";
			when "0100110110" =>
				volume_next <= X"2b1c";
			when "0100110111" =>
				volume_next <= X"2b73";
			when "0100111000" =>
				volume_next <= X"2bca";
			when "0100111001" =>
				volume_next <= X"2c20";
			when "0100111010" =>
				volume_next <= X"2c76";
			when "0100111011" =>
				volume_next <= X"2ccc";
			when "0100111100" =>
				volume_next <= X"2d22";
			when "0100111101" =>
				volume_next <= X"2d77";
			when "0100111110" =>
				volume_next <= X"2dcc";
			when "0100111111" =>
				volume_next <= X"2e20";
			when "0101000000" =>
				volume_next <= X"2e75";
			when "0101000001" =>
				volume_next <= X"2ec9";
			when "0101000010" =>
				volume_next <= X"2f1d";
			when "0101000011" =>
				volume_next <= X"2f70";
			when "0101000100" =>
				volume_next <= X"2fc3";
			when "0101000101" =>
				volume_next <= X"3016";
			when "0101000110" =>
				volume_next <= X"3069";
			when "0101000111" =>
				volume_next <= X"30bb";
			when "0101001000" =>
				volume_next <= X"310d";
			when "0101001001" =>
				volume_next <= X"315f";
			when "0101001010" =>
				volume_next <= X"31b1";
			when "0101001011" =>
				volume_next <= X"3202";
			when "0101001100" =>
				volume_next <= X"3253";
			when "0101001101" =>
				volume_next <= X"32a3";
			when "0101001110" =>
				volume_next <= X"32f4";
			when "0101001111" =>
				volume_next <= X"3344";
			when "0101010000" =>
				volume_next <= X"3394";
			when "0101010001" =>
				volume_next <= X"33e3";
			when "0101010010" =>
				volume_next <= X"3433";
			when "0101010011" =>
				volume_next <= X"3482";
			when "0101010100" =>
				volume_next <= X"34d0";
			when "0101010101" =>
				volume_next <= X"351f";
			when "0101010110" =>
				volume_next <= X"356d";
			when "0101010111" =>
				volume_next <= X"35bb";
			when "0101011000" =>
				volume_next <= X"3609";
			when "0101011001" =>
				volume_next <= X"3656";
			when "0101011010" =>
				volume_next <= X"36a3";
			when "0101011011" =>
				volume_next <= X"36f0";
			when "0101011100" =>
				volume_next <= X"373d";
			when "0101011101" =>
				volume_next <= X"3789";
			when "0101011110" =>
				volume_next <= X"37d5";
			when "0101011111" =>
				volume_next <= X"3821";
			when "0101100000" =>
				volume_next <= X"386c";
			when "0101100001" =>
				volume_next <= X"38b8";
			when "0101100010" =>
				volume_next <= X"3903";
			when "0101100011" =>
				volume_next <= X"394d";
			when "0101100100" =>
				volume_next <= X"3998";
			when "0101100101" =>
				volume_next <= X"39e2";
			when "0101100110" =>
				volume_next <= X"3a2c";
			when "0101100111" =>
				volume_next <= X"3a76";
			when "0101101000" =>
				volume_next <= X"3abf";
			when "0101101001" =>
				volume_next <= X"3b08";
			when "0101101010" =>
				volume_next <= X"3b51";
			when "0101101011" =>
				volume_next <= X"3b9a";
			when "0101101100" =>
				volume_next <= X"3be2";
			when "0101101101" =>
				volume_next <= X"3c2a";
			when "0101101110" =>
				volume_next <= X"3c72";
			when "0101101111" =>
				volume_next <= X"3cba";
			when "0101110000" =>
				volume_next <= X"3d01";
			when "0101110001" =>
				volume_next <= X"3d48";
			when "0101110010" =>
				volume_next <= X"3d8f";
			when "0101110011" =>
				volume_next <= X"3dd5";
			when "0101110100" =>
				volume_next <= X"3e1c";
			when "0101110101" =>
				volume_next <= X"3e62";
			when "0101110110" =>
				volume_next <= X"3ea8";
			when "0101110111" =>
				volume_next <= X"3eed";
			when "0101111000" =>
				volume_next <= X"3f32";
			when "0101111001" =>
				volume_next <= X"3f77";
			when "0101111010" =>
				volume_next <= X"3fbc";
			when "0101111011" =>
				volume_next <= X"4001";
			when "0101111100" =>
				volume_next <= X"4045";
			when "0101111101" =>
				volume_next <= X"4089";
			when "0101111110" =>
				volume_next <= X"40cd";
			when "0101111111" =>
				volume_next <= X"4110";
			when "0110000000" =>
				volume_next <= X"4154";
			when "0110000001" =>
				volume_next <= X"4197";
			when "0110000010" =>
				volume_next <= X"41da";
			when "0110000011" =>
				volume_next <= X"421c";
			when "0110000100" =>
				volume_next <= X"425e";
			when "0110000101" =>
				volume_next <= X"42a1";
			when "0110000110" =>
				volume_next <= X"42e2";
			when "0110000111" =>
				volume_next <= X"4324";
			when "0110001000" =>
				volume_next <= X"4365";
			when "0110001001" =>
				volume_next <= X"43a6";
			when "0110001010" =>
				volume_next <= X"43e7";
			when "0110001011" =>
				volume_next <= X"4428";
			when "0110001100" =>
				volume_next <= X"4468";
			when "0110001101" =>
				volume_next <= X"44a8";
			when "0110001110" =>
				volume_next <= X"44e8";
			when "0110001111" =>
				volume_next <= X"4528";
			when "0110010000" =>
				volume_next <= X"4567";
			when "0110010001" =>
				volume_next <= X"45a6";
			when "0110010010" =>
				volume_next <= X"45e5";
			when "0110010011" =>
				volume_next <= X"4624";
			when "0110010100" =>
				volume_next <= X"4663";
			when "0110010101" =>
				volume_next <= X"46a1";
			when "0110010110" =>
				volume_next <= X"46df";
			when "0110010111" =>
				volume_next <= X"471c";
			when "0110011000" =>
				volume_next <= X"475a";
			when "0110011001" =>
				volume_next <= X"4797";
			when "0110011010" =>
				volume_next <= X"47d4";
			when "0110011011" =>
				volume_next <= X"4811";
			when "0110011100" =>
				volume_next <= X"484e";
			when "0110011101" =>
				volume_next <= X"488a";
			when "0110011110" =>
				volume_next <= X"48c6";
			when "0110011111" =>
				volume_next <= X"4902";
			when "0110100000" =>
				volume_next <= X"493e";
			when "0110100001" =>
				volume_next <= X"4979";
			when "0110100010" =>
				volume_next <= X"49b4";
			when "0110100011" =>
				volume_next <= X"49ef";
			when "0110100100" =>
				volume_next <= X"4a2a";
			when "0110100101" =>
				volume_next <= X"4a65";
			when "0110100110" =>
				volume_next <= X"4a9f";
			when "0110100111" =>
				volume_next <= X"4ad9";
			when "0110101000" =>
				volume_next <= X"4b13";
			when "0110101001" =>
				volume_next <= X"4b4c";
			when "0110101010" =>
				volume_next <= X"4b86";
			when "0110101011" =>
				volume_next <= X"4bbf";
			when "0110101100" =>
				volume_next <= X"4bf8";
			when "0110101101" =>
				volume_next <= X"4c31";
			when "0110101110" =>
				volume_next <= X"4c69";
			when "0110101111" =>
				volume_next <= X"4ca2";
			when "0110110000" =>
				volume_next <= X"4cda";
			when "0110110001" =>
				volume_next <= X"4d11";
			when "0110110010" =>
				volume_next <= X"4d49";
			when "0110110011" =>
				volume_next <= X"4d81";
			when "0110110100" =>
				volume_next <= X"4db8";
			when "0110110101" =>
				volume_next <= X"4def";
			when "0110110110" =>
				volume_next <= X"4e25";
			when "0110110111" =>
				volume_next <= X"4e5c";
			when "0110111000" =>
				volume_next <= X"4e92";
			when "0110111001" =>
				volume_next <= X"4ec8";
			when "0110111010" =>
				volume_next <= X"4efe";
			when "0110111011" =>
				volume_next <= X"4f34";
			when "0110111100" =>
				volume_next <= X"4f69";
			when "0110111101" =>
				volume_next <= X"4f9f";
			when "0110111110" =>
				volume_next <= X"4fd4";
			when "0110111111" =>
				volume_next <= X"5009";
			when "0111000000" =>
				volume_next <= X"503d";
			when "0111000001" =>
				volume_next <= X"5072";
			when "0111000010" =>
				volume_next <= X"50a6";
			when "0111000011" =>
				volume_next <= X"50da";
			when "0111000100" =>
				volume_next <= X"510e";
			when "0111000101" =>
				volume_next <= X"5141";
			when "0111000110" =>
				volume_next <= X"5175";
			when "0111000111" =>
				volume_next <= X"51a8";
			when "0111001000" =>
				volume_next <= X"51db";
			when "0111001001" =>
				volume_next <= X"520d";
			when "0111001010" =>
				volume_next <= X"5240";
			when "0111001011" =>
				volume_next <= X"5272";
			when "0111001100" =>
				volume_next <= X"52a4";
			when "0111001101" =>
				volume_next <= X"52d6";
			when "0111001110" =>
				volume_next <= X"5308";
			when "0111001111" =>
				volume_next <= X"533a";
			when "0111010000" =>
				volume_next <= X"536b";
			when "0111010001" =>
				volume_next <= X"539c";
			when "0111010010" =>
				volume_next <= X"53cd";
			when "0111010011" =>
				volume_next <= X"53fe";
			when "0111010100" =>
				volume_next <= X"542e";
			when "0111010101" =>
				volume_next <= X"545f";
			when "0111010110" =>
				volume_next <= X"548f";
			when "0111010111" =>
				volume_next <= X"54bf";
			when "0111011000" =>
				volume_next <= X"54ee";
			when "0111011001" =>
				volume_next <= X"551e";
			when "0111011010" =>
				volume_next <= X"554d";
			when "0111011011" =>
				volume_next <= X"557c";
			when "0111011100" =>
				volume_next <= X"55ab";
			when "0111011101" =>
				volume_next <= X"55da";
			when "0111011110" =>
				volume_next <= X"5609";
			when "0111011111" =>
				volume_next <= X"5637";
			when "0111100000" =>
				volume_next <= X"5665";
			when "0111100001" =>
				volume_next <= X"5693";
			when "0111100010" =>
				volume_next <= X"56c1";
			when "0111100011" =>
				volume_next <= X"56ef";
			when "0111100100" =>
				volume_next <= X"571c";
			when "0111100101" =>
				volume_next <= X"5749";
			when "0111100110" =>
				volume_next <= X"5776";
			when "0111100111" =>
				volume_next <= X"57a3";
			when "0111101000" =>
				volume_next <= X"57d0";
			when "0111101001" =>
				volume_next <= X"57fc";
			when "0111101010" =>
				volume_next <= X"5829";
			when "0111101011" =>
				volume_next <= X"5855";
			when "0111101100" =>
				volume_next <= X"5881";
			when "0111101101" =>
				volume_next <= X"58ac";
			when "0111101110" =>
				volume_next <= X"58d8";
			when "0111101111" =>
				volume_next <= X"5903";
			when "0111110000" =>
				volume_next <= X"592e";
			when "0111110001" =>
				volume_next <= X"5959";
			when "0111110010" =>
				volume_next <= X"5984";
			when "0111110011" =>
				volume_next <= X"59af";
			when "0111110100" =>
				volume_next <= X"59d9";
			when "0111110101" =>
				volume_next <= X"5a03";
			when "0111110110" =>
				volume_next <= X"5a2e";
			when "0111110111" =>
				volume_next <= X"5a57";
			when "0111111000" =>
				volume_next <= X"5a81";
			when "0111111001" =>
				volume_next <= X"5aab";
			when "0111111010" =>
				volume_next <= X"5ad4";
			when "0111111011" =>
				volume_next <= X"5afd";
			when "0111111100" =>
				volume_next <= X"5b26";
			when "0111111101" =>
				volume_next <= X"5b4f";
			when "0111111110" =>
				volume_next <= X"5b78";
			when "0111111111" =>
				volume_next <= X"5ba0";
			when "1000000000" =>
				volume_next <= X"5bc9";
			when "1000000001" =>
				volume_next <= X"5bf1";
			when "1000000010" =>
				volume_next <= X"5c19";
			when "1000000011" =>
				volume_next <= X"5c41";
			when "1000000100" =>
				volume_next <= X"5c68";
			when "1000000101" =>
				volume_next <= X"5c90";
			when "1000000110" =>
				volume_next <= X"5cb7";
			when "1000000111" =>
				volume_next <= X"5cde";
			when "1000001000" =>
				volume_next <= X"5d05";
			when "1000001001" =>
				volume_next <= X"5d2c";
			when "1000001010" =>
				volume_next <= X"5d52";
			when "1000001011" =>
				volume_next <= X"5d79";
			when "1000001100" =>
				volume_next <= X"5d9f";
			when "1000001101" =>
				volume_next <= X"5dc5";
			when "1000001110" =>
				volume_next <= X"5deb";
			when "1000001111" =>
				volume_next <= X"5e11";
			when "1000010000" =>
				volume_next <= X"5e36";
			when "1000010001" =>
				volume_next <= X"5e5c";
			when "1000010010" =>
				volume_next <= X"5e81";
			when "1000010011" =>
				volume_next <= X"5ea6";
			when "1000010100" =>
				volume_next <= X"5ecb";
			when "1000010101" =>
				volume_next <= X"5ef0";
			when "1000010110" =>
				volume_next <= X"5f15";
			when "1000010111" =>
				volume_next <= X"5f39";
			when "1000011000" =>
				volume_next <= X"5f5d";
			when "1000011001" =>
				volume_next <= X"5f82";
			when "1000011010" =>
				volume_next <= X"5fa6";
			when "1000011011" =>
				volume_next <= X"5fc9";
			when "1000011100" =>
				volume_next <= X"5fed";
			when "1000011101" =>
				volume_next <= X"6011";
			when "1000011110" =>
				volume_next <= X"6034";
			when "1000011111" =>
				volume_next <= X"6057";
			when "1000100000" =>
				volume_next <= X"607a";
			when "1000100001" =>
				volume_next <= X"609d";
			when "1000100010" =>
				volume_next <= X"60c0";
			when "1000100011" =>
				volume_next <= X"60e3";
			when "1000100100" =>
				volume_next <= X"6105";
			when "1000100101" =>
				volume_next <= X"6127";
			when "1000100110" =>
				volume_next <= X"6149";
			when "1000100111" =>
				volume_next <= X"616b";
			when "1000101000" =>
				volume_next <= X"618d";
			when "1000101001" =>
				volume_next <= X"61af";
			when "1000101010" =>
				volume_next <= X"61d0";
			when "1000101011" =>
				volume_next <= X"61f2";
			when "1000101100" =>
				volume_next <= X"6213";
			when "1000101101" =>
				volume_next <= X"6234";
			when "1000101110" =>
				volume_next <= X"6255";
			when "1000101111" =>
				volume_next <= X"6276";
			when "1000110000" =>
				volume_next <= X"6296";
			when "1000110001" =>
				volume_next <= X"62b7";
			when "1000110010" =>
				volume_next <= X"62d7";
			when "1000110011" =>
				volume_next <= X"62f7";
			when "1000110100" =>
				volume_next <= X"6318";
			when "1000110101" =>
				volume_next <= X"6337";
			when "1000110110" =>
				volume_next <= X"6357";
			when "1000110111" =>
				volume_next <= X"6377";
			when "1000111000" =>
				volume_next <= X"6396";
			when "1000111001" =>
				volume_next <= X"63b6";
			when "1000111010" =>
				volume_next <= X"63d5";
			when "1000111011" =>
				volume_next <= X"63f4";
			when "1000111100" =>
				volume_next <= X"6413";
			when "1000111101" =>
				volume_next <= X"6432";
			when "1000111110" =>
				volume_next <= X"6450";
			when "1000111111" =>
				volume_next <= X"646f";
			when "1001000000" =>
				volume_next <= X"648d";
			when "1001000001" =>
				volume_next <= X"64ab";
			when "1001000010" =>
				volume_next <= X"64ca";
			when "1001000011" =>
				volume_next <= X"64e8";
			when "1001000100" =>
				volume_next <= X"6505";
			when "1001000101" =>
				volume_next <= X"6523";
			when "1001000110" =>
				volume_next <= X"6541";
			when "1001000111" =>
				volume_next <= X"655e";
			when "1001001000" =>
				volume_next <= X"657b";
			when "1001001001" =>
				volume_next <= X"6599";
			when "1001001010" =>
				volume_next <= X"65b6";
			when "1001001011" =>
				volume_next <= X"65d3";
			when "1001001100" =>
				volume_next <= X"65ef";
			when "1001001101" =>
				volume_next <= X"660c";
			when "1001001110" =>
				volume_next <= X"6628";
			when "1001001111" =>
				volume_next <= X"6645";
			when "1001010000" =>
				volume_next <= X"6661";
			when "1001010001" =>
				volume_next <= X"667d";
			when "1001010010" =>
				volume_next <= X"6699";
			when "1001010011" =>
				volume_next <= X"66b5";
			when "1001010100" =>
				volume_next <= X"66d1";
			when "1001010101" =>
				volume_next <= X"66ed";
			when "1001010110" =>
				volume_next <= X"6708";
			when "1001010111" =>
				volume_next <= X"6723";
			when "1001011000" =>
				volume_next <= X"673f";
			when "1001011001" =>
				volume_next <= X"675a";
			when "1001011010" =>
				volume_next <= X"6775";
			when "1001011011" =>
				volume_next <= X"6790";
			when "1001011100" =>
				volume_next <= X"67ab";
			when "1001011101" =>
				volume_next <= X"67c5";
			when "1001011110" =>
				volume_next <= X"67e0";
			when "1001011111" =>
				volume_next <= X"67fa";
			when "1001100000" =>
				volume_next <= X"6814";
			when "1001100001" =>
				volume_next <= X"682f";
			when "1001100010" =>
				volume_next <= X"6849";
			when "1001100011" =>
				volume_next <= X"6863";
			when "1001100100" =>
				volume_next <= X"687c";
			when "1001100101" =>
				volume_next <= X"6896";
			when "1001100110" =>
				volume_next <= X"68b0";
			when "1001100111" =>
				volume_next <= X"68c9";
			when "1001101000" =>
				volume_next <= X"68e3";
			when "1001101001" =>
				volume_next <= X"68fc";
			when "1001101010" =>
				volume_next <= X"6915";
			when "1001101011" =>
				volume_next <= X"692e";
			when "1001101100" =>
				volume_next <= X"6947";
			when "1001101101" =>
				volume_next <= X"6960";
			when "1001101110" =>
				volume_next <= X"6978";
			when "1001101111" =>
				volume_next <= X"6991";
			when "1001110000" =>
				volume_next <= X"69a9";
			when "1001110001" =>
				volume_next <= X"69c2";
			when "1001110010" =>
				volume_next <= X"69da";
			when "1001110011" =>
				volume_next <= X"69f2";
			when "1001110100" =>
				volume_next <= X"6a0a";
			when "1001110101" =>
				volume_next <= X"6a22";
			when "1001110110" =>
				volume_next <= X"6a3a";
			when "1001110111" =>
				volume_next <= X"6a52";
			when "1001111000" =>
				volume_next <= X"6a69";
			when "1001111001" =>
				volume_next <= X"6a81";
			when "1001111010" =>
				volume_next <= X"6a98";
			when "1001111011" =>
				volume_next <= X"6ab0";
			when "1001111100" =>
				volume_next <= X"6ac7";
			when "1001111101" =>
				volume_next <= X"6ade";
			when "1001111110" =>
				volume_next <= X"6af5";
			when "1001111111" =>
				volume_next <= X"6b0c";
			when "1010000000" =>
				volume_next <= X"6b23";
			when "1010000001" =>
				volume_next <= X"6b39";
			when "1010000010" =>
				volume_next <= X"6b50";
			when "1010000011" =>
				volume_next <= X"6b67";
			when "1010000100" =>
				volume_next <= X"6b7d";
			when "1010000101" =>
				volume_next <= X"6b93";
			when "1010000110" =>
				volume_next <= X"6ba9";
			when "1010000111" =>
				volume_next <= X"6bc0";
			when "1010001000" =>
				volume_next <= X"6bd6";
			when "1010001001" =>
				volume_next <= X"6bec";
			when "1010001010" =>
				volume_next <= X"6c01";
			when "1010001011" =>
				volume_next <= X"6c17";
			when "1010001100" =>
				volume_next <= X"6c2d";
			when "1010001101" =>
				volume_next <= X"6c42";
			when "1010001110" =>
				volume_next <= X"6c58";
			when "1010001111" =>
				volume_next <= X"6c6d";
			when "1010010000" =>
				volume_next <= X"6c82";
			when "1010010001" =>
				volume_next <= X"6c98";
			when "1010010010" =>
				volume_next <= X"6cad";
			when "1010010011" =>
				volume_next <= X"6cc2";
			when "1010010100" =>
				volume_next <= X"6cd7";
			when "1010010101" =>
				volume_next <= X"6ceb";
			when "1010010110" =>
				volume_next <= X"6d00";
			when "1010010111" =>
				volume_next <= X"6d15";
			when "1010011000" =>
				volume_next <= X"6d29";
			when "1010011001" =>
				volume_next <= X"6d3e";
			when "1010011010" =>
				volume_next <= X"6d52";
			when "1010011011" =>
				volume_next <= X"6d67";
			when "1010011100" =>
				volume_next <= X"6d7b";
			when "1010011101" =>
				volume_next <= X"6d8f";
			when "1010011110" =>
				volume_next <= X"6da3";
			when "1010011111" =>
				volume_next <= X"6db7";
			when "1010100000" =>
				volume_next <= X"6dcb";
			when "1010100001" =>
				volume_next <= X"6ddf";
			when "1010100010" =>
				volume_next <= X"6df3";
			when "1010100011" =>
				volume_next <= X"6e06";
			when "1010100100" =>
				volume_next <= X"6e1a";
			when "1010100101" =>
				volume_next <= X"6e2d";
			when "1010100110" =>
				volume_next <= X"6e41";
			when "1010100111" =>
				volume_next <= X"6e54";
			when "1010101000" =>
				volume_next <= X"6e67";
			when "1010101001" =>
				volume_next <= X"6e7b";
			when "1010101010" =>
				volume_next <= X"6e8e";
			when "1010101011" =>
				volume_next <= X"6ea1";
			when "1010101100" =>
				volume_next <= X"6eb4";
			when "1010101101" =>
				volume_next <= X"6ec7";
			when "1010101110" =>
				volume_next <= X"6ed9";
			when "1010101111" =>
				volume_next <= X"6eec";
			when "1010110000" =>
				volume_next <= X"6eff";
			when "1010110001" =>
				volume_next <= X"6f11";
			when "1010110010" =>
				volume_next <= X"6f24";
			when "1010110011" =>
				volume_next <= X"6f36";
			when "1010110100" =>
				volume_next <= X"6f49";
			when "1010110101" =>
				volume_next <= X"6f5b";
			when "1010110110" =>
				volume_next <= X"6f6d";
			when "1010110111" =>
				volume_next <= X"6f80";
			when "1010111000" =>
				volume_next <= X"6f92";
			when "1010111001" =>
				volume_next <= X"6fa4";
			when "1010111010" =>
				volume_next <= X"6fb6";
			when "1010111011" =>
				volume_next <= X"6fc8";
			when "1010111100" =>
				volume_next <= X"6fda";
			when "1010111101" =>
				volume_next <= X"6feb";
			when "1010111110" =>
				volume_next <= X"6ffd";
			when "1010111111" =>
				volume_next <= X"700f";
			when "1011000000" =>
				volume_next <= X"7020";
			when "1011000001" =>
				volume_next <= X"7032";
			when "1011000010" =>
				volume_next <= X"7043";
			when "1011000011" =>
				volume_next <= X"7055";
			when "1011000100" =>
				volume_next <= X"7066";
			when "1011000101" =>
				volume_next <= X"7077";
			when "1011000110" =>
				volume_next <= X"7089";
			when "1011000111" =>
				volume_next <= X"709a";
			when "1011001000" =>
				volume_next <= X"70ab";
			when "1011001001" =>
				volume_next <= X"70bc";
			when "1011001010" =>
				volume_next <= X"70cd";
			when "1011001011" =>
				volume_next <= X"70de";
			when "1011001100" =>
				volume_next <= X"70ef";
			when "1011001101" =>
				volume_next <= X"7100";
			when "1011001110" =>
				volume_next <= X"7110";
			when "1011001111" =>
				volume_next <= X"7121";
			when "1011010000" =>
				volume_next <= X"7132";
			when "1011010001" =>
				volume_next <= X"7142";
			when "1011010010" =>
				volume_next <= X"7153";
			when "1011010011" =>
				volume_next <= X"7163";
			when "1011010100" =>
				volume_next <= X"7174";
			when "1011010101" =>
				volume_next <= X"7184";
			when "1011010110" =>
				volume_next <= X"7195";
			when "1011010111" =>
				volume_next <= X"71a5";
			when "1011011000" =>
				volume_next <= X"71b5";
			when "1011011001" =>
				volume_next <= X"71c5";
			when "1011011010" =>
				volume_next <= X"71d6";
			when "1011011011" =>
				volume_next <= X"71e6";
			when "1011011100" =>
				volume_next <= X"71f6";
			when "1011011101" =>
				volume_next <= X"7206";
			when "1011011110" =>
				volume_next <= X"7216";
			when "1011011111" =>
				volume_next <= X"7226";
			when "1011100000" =>
				volume_next <= X"7236";
			when "1011100001" =>
				volume_next <= X"7245";
			when "1011100010" =>
				volume_next <= X"7255";
			when "1011100011" =>
				volume_next <= X"7265";
			when "1011100100" =>
				volume_next <= X"7275";
			when "1011100101" =>
				volume_next <= X"7284";
			when "1011100110" =>
				volume_next <= X"7294";
			when "1011100111" =>
				volume_next <= X"72a4";
			when "1011101000" =>
				volume_next <= X"72b3";
			when "1011101001" =>
				volume_next <= X"72c3";
			when "1011101010" =>
				volume_next <= X"72d2";
			when "1011101011" =>
				volume_next <= X"72e2";
			when "1011101100" =>
				volume_next <= X"72f1";
			when "1011101101" =>
				volume_next <= X"7300";
			when "1011101110" =>
				volume_next <= X"7310";
			when "1011101111" =>
				volume_next <= X"731f";
			when "1011110000" =>
				volume_next <= X"732e";
			when "1011110001" =>
				volume_next <= X"733d";
			when "1011110010" =>
				volume_next <= X"734d";
			when "1011110011" =>
				volume_next <= X"735c";
			when "1011110100" =>
				volume_next <= X"736b";
			when "1011110101" =>
				volume_next <= X"737a";
			when "1011110110" =>
				volume_next <= X"7389";
			when "1011110111" =>
				volume_next <= X"7398";
			when "1011111000" =>
				volume_next <= X"73a7";
			when "1011111001" =>
				volume_next <= X"73b6";
			when "1011111010" =>
				volume_next <= X"73c5";
			when "1011111011" =>
				volume_next <= X"73d4";
			when "1011111100" =>
				volume_next <= X"73e3";
			when "1011111101" =>
				volume_next <= X"73f1";
			when "1011111110" =>
				volume_next <= X"7400";
			when "1011111111" =>
				volume_next <= X"740f";
			when "1100000000" =>
				volume_next <= X"741e";
			when "1100000001" =>
				volume_next <= X"742c";
			when "1100000010" =>
				volume_next <= X"743b";
			when "1100000011" =>
				volume_next <= X"744a";
			when "1100000100" =>
				volume_next <= X"7459";
			when "1100000101" =>
				volume_next <= X"7467";
			when "1100000110" =>
				volume_next <= X"7476";
			when "1100000111" =>
				volume_next <= X"7484";
			when "1100001000" =>
				volume_next <= X"7493";
			when "1100001001" =>
				volume_next <= X"74a1";
			when "1100001010" =>
				volume_next <= X"74b0";
			when "1100001011" =>
				volume_next <= X"74be";
			when "1100001100" =>
				volume_next <= X"74cd";
			when "1100001101" =>
				volume_next <= X"74db";
			when "1100001110" =>
				volume_next <= X"74ea";
			when "1100001111" =>
				volume_next <= X"74f8";
			when "1100010000" =>
				volume_next <= X"7507";
			when "1100010001" =>
				volume_next <= X"7515";
			when "1100010010" =>
				volume_next <= X"7524";
			when "1100010011" =>
				volume_next <= X"7532";
			when "1100010100" =>
				volume_next <= X"7540";
			when "1100010101" =>
				volume_next <= X"754f";
			when "1100010110" =>
				volume_next <= X"755d";
			when "1100010111" =>
				volume_next <= X"756b";
			when "1100011000" =>
				volume_next <= X"757a";
			when "1100011001" =>
				volume_next <= X"7588";
			when "1100011010" =>
				volume_next <= X"7596";
			when "1100011011" =>
				volume_next <= X"75a4";
			when "1100011100" =>
				volume_next <= X"75b3";
			when "1100011101" =>
				volume_next <= X"75c1";
			when "1100011110" =>
				volume_next <= X"75cf";
			when "1100011111" =>
				volume_next <= X"75dd";
			when "1100100000" =>
				volume_next <= X"75ec";
			when "1100100001" =>
				volume_next <= X"75fa";
			when "1100100010" =>
				volume_next <= X"7608";
			when "1100100011" =>
				volume_next <= X"7616";
			when "1100100100" =>
				volume_next <= X"7624";
			when "1100100101" =>
				volume_next <= X"7633";
			when "1100100110" =>
				volume_next <= X"7641";
			when "1100100111" =>
				volume_next <= X"764f";
			when "1100101000" =>
				volume_next <= X"765d";
			when "1100101001" =>
				volume_next <= X"766b";
			when "1100101010" =>
				volume_next <= X"767a";
			when "1100101011" =>
				volume_next <= X"7688";
			when "1100101100" =>
				volume_next <= X"7696";
			when "1100101101" =>
				volume_next <= X"76a4";
			when "1100101110" =>
				volume_next <= X"76b2";
			when "1100101111" =>
				volume_next <= X"76c0";
			when "1100110000" =>
				volume_next <= X"76cf";
			when "1100110001" =>
				volume_next <= X"76dd";
			when "1100110010" =>
				volume_next <= X"76eb";
			when "1100110011" =>
				volume_next <= X"76f9";
			when "1100110100" =>
				volume_next <= X"7707";
			when "1100110101" =>
				volume_next <= X"7716";
			when "1100110110" =>
				volume_next <= X"7724";
			when "1100110111" =>
				volume_next <= X"7732";
			when "1100111000" =>
				volume_next <= X"7740";
			when "1100111001" =>
				volume_next <= X"774e";
			when "1100111010" =>
				volume_next <= X"775d";
			when "1100111011" =>
				volume_next <= X"776b";
			when "1100111100" =>
				volume_next <= X"7779";
			when "1100111101" =>
				volume_next <= X"7787";
			when "1100111110" =>
				volume_next <= X"7796";
			when "1100111111" =>
				volume_next <= X"77a4";
			when "1101000000" =>
				volume_next <= X"77b2";
			when "1101000001" =>
				volume_next <= X"77c1";
			when "1101000010" =>
				volume_next <= X"77cf";
			when "1101000011" =>
				volume_next <= X"77dd";
			when "1101000100" =>
				volume_next <= X"77eb";
			when "1101000101" =>
				volume_next <= X"77fa";
			when "1101000110" =>
				volume_next <= X"7808";
			when "1101000111" =>
				volume_next <= X"7817";
			when "1101001000" =>
				volume_next <= X"7825";
			when "1101001001" =>
				volume_next <= X"7833";
			when "1101001010" =>
				volume_next <= X"7842";
			when "1101001011" =>
				volume_next <= X"7850";
			when "1101001100" =>
				volume_next <= X"785f";
			when "1101001101" =>
				volume_next <= X"786d";
			when "1101001110" =>
				volume_next <= X"787c";
			when "1101001111" =>
				volume_next <= X"788a";
			when "1101010000" =>
				volume_next <= X"7899";
			when "1101010001" =>
				volume_next <= X"78a7";
			when "1101010010" =>
				volume_next <= X"78b6";
			when "1101010011" =>
				volume_next <= X"78c4";
			when "1101010100" =>
				volume_next <= X"78d3";
			when "1101010101" =>
				volume_next <= X"78e2";
			when "1101010110" =>
				volume_next <= X"78f0";
			when "1101010111" =>
				volume_next <= X"78ff";
			when "1101011000" =>
				volume_next <= X"790e";
			when "1101011001" =>
				volume_next <= X"791d";
			when "1101011010" =>
				volume_next <= X"792b";
			when "1101011011" =>
				volume_next <= X"793a";
			when "1101011100" =>
				volume_next <= X"7949";
			when "1101011101" =>
				volume_next <= X"7958";
			when "1101011110" =>
				volume_next <= X"7967";
			when "1101011111" =>
				volume_next <= X"7976";
			when "1101100000" =>
				volume_next <= X"7984";
			when "1101100001" =>
				volume_next <= X"7993";
			when "1101100010" =>
				volume_next <= X"79a2";
			when "1101100011" =>
				volume_next <= X"79b1";
			when "1101100100" =>
				volume_next <= X"79c1";
			when "1101100101" =>
				volume_next <= X"79d0";
			when "1101100110" =>
				volume_next <= X"79df";
			when "1101100111" =>
				volume_next <= X"79ee";
			when "1101101000" =>
				volume_next <= X"79fd";
			when "1101101001" =>
				volume_next <= X"7a0c";
			when "1101101010" =>
				volume_next <= X"7a1c";
			when "1101101011" =>
				volume_next <= X"7a2b";
			when "1101101100" =>
				volume_next <= X"7a3a";
			when "1101101101" =>
				volume_next <= X"7a4a";
			when "1101101110" =>
				volume_next <= X"7a59";
			when "1101101111" =>
				volume_next <= X"7a68";
			when "1101110000" =>
				volume_next <= X"7a78";
			when "1101110001" =>
				volume_next <= X"7a87";
			when "1101110010" =>
				volume_next <= X"7a97";
			when "1101110011" =>
				volume_next <= X"7aa7";
			when "1101110100" =>
				volume_next <= X"7ab6";
			when "1101110101" =>
				volume_next <= X"7ac6";
			when "1101110110" =>
				volume_next <= X"7ad6";
			when "1101110111" =>
				volume_next <= X"7ae5";
			when "1101111000" =>
				volume_next <= X"7af5";
			when "1101111001" =>
				volume_next <= X"7b05";
			when "1101111010" =>
				volume_next <= X"7b15";
			when "1101111011" =>
				volume_next <= X"7b25";
			when "1101111100" =>
				volume_next <= X"7b35";
			when "1101111101" =>
				volume_next <= X"7b45";
			when "1101111110" =>
				volume_next <= X"7b55";
			when "1101111111" =>
				volume_next <= X"7b65";
			when "1110000000" =>
				volume_next <= X"7b75";
			when "1110000001" =>
				volume_next <= X"7b86";
			when "1110000010" =>
				volume_next <= X"7b96";
			when "1110000011" =>
				volume_next <= X"7ba6";
			when "1110000100" =>
				volume_next <= X"7bb7";
			when "1110000101" =>
				volume_next <= X"7bc7";
			when "1110000110" =>
				volume_next <= X"7bd7";
			when "1110000111" =>
				volume_next <= X"7be8";
			when "1110001000" =>
				volume_next <= X"7bf9";
			when "1110001001" =>
				volume_next <= X"7c09";
			when "1110001010" =>
				volume_next <= X"7c1a";
			when "1110001011" =>
				volume_next <= X"7c2b";
			when "1110001100" =>
				volume_next <= X"7c3b";
			when "1110001101" =>
				volume_next <= X"7c4c";
			when "1110001110" =>
				volume_next <= X"7c5d";
			when "1110001111" =>
				volume_next <= X"7c6e";
			when "1110010000" =>
				volume_next <= X"7c7f";
			when "1110010001" =>
				volume_next <= X"7c90";
			when "1110010010" =>
				volume_next <= X"7ca1";
			when "1110010011" =>
				volume_next <= X"7cb3";
			when "1110010100" =>
				volume_next <= X"7cc4";
			when "1110010101" =>
				volume_next <= X"7cd5";
			when "1110010110" =>
				volume_next <= X"7ce6";
			when "1110010111" =>
				volume_next <= X"7cf8";
			when "1110011000" =>
				volume_next <= X"7d09";
			when "1110011001" =>
				volume_next <= X"7d1b";
			when "1110011010" =>
				volume_next <= X"7d2d";
			when "1110011011" =>
				volume_next <= X"7d3e";
			when "1110011100" =>
				volume_next <= X"7d50";
			when "1110011101" =>
				volume_next <= X"7d62";
			when "1110011110" =>
				volume_next <= X"7d74";
			when "1110011111" =>
				volume_next <= X"7d86";
			when "1110100000" =>
				volume_next <= X"7d98";
			when "1110100001" =>
				volume_next <= X"7daa";
			when "1110100010" =>
				volume_next <= X"7dbc";
			when "1110100011" =>
				volume_next <= X"7dce";
			when "1110100100" =>
				volume_next <= X"7de0";
			when "1110100101" =>
				volume_next <= X"7df3";
			when "1110100110" =>
				volume_next <= X"7e05";
			when "1110100111" =>
				volume_next <= X"7e18";
			when "1110101000" =>
				volume_next <= X"7e2a";
			when "1110101001" =>
				volume_next <= X"7e3d";
			when "1110101010" =>
				volume_next <= X"7e50";
			when "1110101011" =>
				volume_next <= X"7e62";
			when "1110101100" =>
				volume_next <= X"7e75";
			when "1110101101" =>
				volume_next <= X"7e88";
			when "1110101110" =>
				volume_next <= X"7e9b";
			when "1110101111" =>
				volume_next <= X"7eae";
			when "1110110000" =>
				volume_next <= X"7ec1";
			when "1110110001" =>
				volume_next <= X"7ed5";
			when "1110110010" =>
				volume_next <= X"7ee8";
			when "1110110011" =>
				volume_next <= X"7efb";
			when "1110110100" =>
				volume_next <= X"7f0f";
			when "1110110101" =>
				volume_next <= X"7f22";
			when "1110110110" =>
				volume_next <= X"7f36";
			when "1110110111" =>
				volume_next <= X"7f4a";
			when "1110111000" =>
				volume_next <= X"7f5d";
			when "1110111001" =>
				volume_next <= X"7f71";
			when "1110111010" =>
				volume_next <= X"7f85";
			when "1110111011" =>
				volume_next <= X"7f99";
			when "1110111100" =>
				volume_next <= X"7fad";
			when "1110111101" =>
				volume_next <= X"7fc1";
			when "1110111110" =>
				volume_next <= X"7fd6";
			when "1110111111" =>
				volume_next <= X"7fea";
			when "1111000000" =>
				volume_next <= X"7fff";
			when others =>
				volume_next <= X"7fff";
		end case;
        end process;

	-- output
	volume_out_next <= volume_next;
		
END vhdl;
