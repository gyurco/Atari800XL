
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80ef",
X"fc738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80f3",
X"d40c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580ea",
X"ac2d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580e8c0",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80d09c04",
X"fc3d0d76",
X"705255b3",
X"fa3f83e0",
X"800815ff",
X"05547375",
X"2e8e3873",
X"335372ae",
X"2e8638ff",
X"1454ef39",
X"77528114",
X"51b3923f",
X"83e08008",
X"307083e0",
X"80080780",
X"2583e080",
X"0c53863d",
X"0d04fc3d",
X"0d767052",
X"559ab13f",
X"83e08008",
X"54815383",
X"e0800880",
X"c7387451",
X"99f43f83",
X"e080080b",
X"0b80f1e0",
X"5383e080",
X"085253ff",
X"8f3f83e0",
X"8008a538",
X"0b0b80f1",
X"e4527251",
X"fefe3f83",
X"e0800894",
X"380b0b80",
X"f1e85272",
X"51feed3f",
X"83e08008",
X"802e8338",
X"81547353",
X"7283e080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"99ca3f81",
X"5383e080",
X"08993873",
X"5199933f",
X"0b0b80f1",
X"ec5283e0",
X"800851fe",
X"b33f83e0",
X"80085372",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"70525499",
X"973f8153",
X"83e08008",
X"99387351",
X"98e03f0b",
X"0b80f1f0",
X"5283e080",
X"0851fe80",
X"3f83e080",
X"08537283",
X"e0800c85",
X"3d0d04e0",
X"3d0da33d",
X"0870525e",
X"8f873f83",
X"e0800833",
X"943d5654",
X"73943880",
X"f6f05274",
X"5184c639",
X"7d527851",
X"92863f84",
X"d0397d51",
X"8eef3f83",
X"e0800852",
X"74518e9f",
X"3f83e09c",
X"0852933d",
X"70525d94",
X"f73f83e0",
X"80085980",
X"0b83e080",
X"08555b83",
X"e080087b",
X"2e943881",
X"1b74525b",
X"97f93f83",
X"e0800854",
X"83e08008",
X"ee38805a",
X"ff7a437a",
X"427a415f",
X"7909709f",
X"2c7b065b",
X"547a7a24",
X"8438ff1b",
X"5af61a70",
X"09709f2c",
X"72067bff",
X"125a5a52",
X"55558075",
X"25953876",
X"5197b83f",
X"83e08008",
X"76ff1858",
X"55577380",
X"24ed3874",
X"7f2e8638",
X"b9c63f74",
X"5f78ff1b",
X"70585d58",
X"807a2595",
X"38775197",
X"8e3f83e0",
X"800876ff",
X"18585558",
X"738024ed",
X"38800b83",
X"e3980c80",
X"0b83e3b8",
X"0c0b0b80",
X"f1f4518b",
X"e33f8180",
X"0b83e3b8",
X"0c0b0b80",
X"f1fc518b",
X"d33fa80b",
X"83e3980c",
X"76802e80",
X"e83883e3",
X"98087779",
X"32703070",
X"72078025",
X"70872b83",
X"e3b80c51",
X"56785356",
X"5696c13f",
X"83e08008",
X"802e8a38",
X"0b0b80f2",
X"84518b98",
X"3f765196",
X"813f83e0",
X"8008520b",
X"0b80f390",
X"518b853f",
X"76519687",
X"3f83e080",
X"0883e398",
X"08555775",
X"74258638",
X"a81656f7",
X"397583e3",
X"980c86f0",
X"7624ff94",
X"3887980b",
X"83e3980c",
X"77802eb7",
X"38775195",
X"bd3f83e0",
X"80087852",
X"5595dd3f",
X"0b0b80f2",
X"8c5483e0",
X"80088f38",
X"87398076",
X"34fd9639",
X"0b0b80f2",
X"88547453",
X"73520b0b",
X"80f1d451",
X"8a9e3f80",
X"540b0b80",
X"f3d0518a",
X"933f8114",
X"5473a82e",
X"098106ed",
X"38868da0",
X"51b5c53f",
X"8052903d",
X"70525480",
X"d5d83f83",
X"52735180",
X"d5d03f61",
X"802e80ff",
X"387b5473",
X"ff2e9638",
X"78802e81",
X"80387851",
X"94dd3f83",
X"e08008ff",
X"155559e7",
X"3978802e",
X"80eb3878",
X"5194d93f",
X"83e08008",
X"802efc84",
X"38785194",
X"a13f83e0",
X"8008520b",
X"0b80f1dc",
X"51ac813f",
X"83e08008",
X"a4387c51",
X"adb93f83",
X"e0800855",
X"74ff1656",
X"54807425",
X"fbef3874",
X"1d703355",
X"5673af2e",
X"fec838e8",
X"39785193",
X"df3f83e0",
X"8008527c",
X"51acf03f",
X"fbcf397f",
X"88296010",
X"057a0561",
X"055afc80",
X"39a23d0d",
X"04fe3d0d",
X"80f5f808",
X"70337081",
X"ff067084",
X"2a813281",
X"06555152",
X"5371802e",
X"8c38a873",
X"3480f5f8",
X"0851b871",
X"347183e0",
X"800c843d",
X"0d04fe3d",
X"0d80f5f8",
X"08703370",
X"81ff0670",
X"852a8132",
X"81065551",
X"52537180",
X"2e8c3898",
X"733480f5",
X"f80851b8",
X"71347183",
X"e0800c84",
X"3d0d0480",
X"3d0d80f5",
X"f4085193",
X"713480f6",
X"800851ff",
X"7134823d",
X"0d04fe3d",
X"0d029305",
X"3380f5f4",
X"08535380",
X"72348a51",
X"b38e3fd3",
X"3f80f684",
X"085280f8",
X"723480f6",
X"9c085280",
X"7234fa13",
X"80f6a408",
X"53537272",
X"3480f68c",
X"08528072",
X"3480f694",
X"08527272",
X"3480f5f8",
X"08528072",
X"3480f5f8",
X"0852b872",
X"34843d0d",
X"04ff3d0d",
X"028f0533",
X"80f5fc08",
X"52527171",
X"34fe9e3f",
X"83e08008",
X"802ef638",
X"833d0d04",
X"803d0d84",
X"39bbf33f",
X"feb83f83",
X"e0800880",
X"2ef33880",
X"f5fc0870",
X"337081ff",
X"0683e080",
X"0c515182",
X"3d0d0480",
X"3d0d80f5",
X"f40851a3",
X"713480f6",
X"800851ff",
X"713480f5",
X"f80851a8",
X"713480f5",
X"f80851b8",
X"7134823d",
X"0d04803d",
X"0d80f5f4",
X"08703370",
X"81c00670",
X"30708025",
X"83e0800c",
X"51515151",
X"823d0d04",
X"ff3d0d80",
X"f5f80870",
X"337081ff",
X"0670832a",
X"81327081",
X"06515151",
X"52527080",
X"2ee538b0",
X"723480f5",
X"f80851b8",
X"7134833d",
X"0d04803d",
X"0d80f6b0",
X"08700881",
X"0683e080",
X"0c51823d",
X"0d04fd3d",
X"0d757754",
X"54807325",
X"94387370",
X"81055533",
X"5280f290",
X"5185a13f",
X"ff1353e9",
X"39853d0d",
X"04f63d0d",
X"7c7e6062",
X"5a5d5b56",
X"80598155",
X"8539747a",
X"29557452",
X"755180d3",
X"bd3f83e0",
X"80087a27",
X"ed387480",
X"2e80e038",
X"74527551",
X"80d3a73f",
X"83e08008",
X"75537652",
X"5480d3cd",
X"3f83e080",
X"087a5375",
X"525680d3",
X"8d3f83e0",
X"80087930",
X"707b079f",
X"2a707780",
X"24075151",
X"54557287",
X"3883e080",
X"08c23876",
X"8118b016",
X"55585889",
X"74258b38",
X"b714537a",
X"853880d7",
X"14537278",
X"34811959",
X"ff9c3980",
X"77348c3d",
X"0d04f73d",
X"0d7b7d7f",
X"62029005",
X"bb053357",
X"59565a5a",
X"b0587283",
X"38a05875",
X"70708105",
X"52337159",
X"54559039",
X"8074258e",
X"38ff1477",
X"70810559",
X"33545472",
X"ef3873ff",
X"15555380",
X"73258938",
X"77527951",
X"782def39",
X"75337557",
X"5372802e",
X"90387252",
X"7951782d",
X"75708105",
X"573353ed",
X"398b3d0d",
X"04ee3d0d",
X"64666969",
X"70708105",
X"52335b4a",
X"5c5e5e76",
X"802e82f9",
X"3876a52e",
X"09810682",
X"e0388070",
X"41677070",
X"81055233",
X"714a5957",
X"5f76b02e",
X"0981068c",
X"38757081",
X"05573376",
X"4857815f",
X"d0175675",
X"892680da",
X"3876675c",
X"59805c93",
X"39778a24",
X"80c3387b",
X"8a29187b",
X"7081055d",
X"335a5cd0",
X"197081ff",
X"06585889",
X"7727a438",
X"ff9f1970",
X"81ff06ff",
X"a91b5a51",
X"56857627",
X"9238ffbf",
X"197081ff",
X"06515675",
X"85268a38",
X"c9195877",
X"8025ffb9",
X"387a477b",
X"407881ff",
X"06577680",
X"e42e80e5",
X"387680e4",
X"24a73876",
X"80d82e81",
X"86387680",
X"d8249038",
X"76802e81",
X"cc3876a5",
X"2e81b638",
X"81b93976",
X"80e32e81",
X"8c3881af",
X"397680f5",
X"2e9b3876",
X"80f5248b",
X"387680f3",
X"2e818138",
X"81993976",
X"80f82e80",
X"ca38818f",
X"39913d70",
X"55578053",
X"8a527984",
X"1b710853",
X"5b56fbfd",
X"3f7655ab",
X"3979841b",
X"7108943d",
X"705b5b52",
X"5b567580",
X"258c3875",
X"3056ad78",
X"340280c1",
X"05577654",
X"80538a52",
X"7551fbd1",
X"3f77557e",
X"54b83991",
X"3d705577",
X"80d83270",
X"30708025",
X"56515856",
X"90527984",
X"1b710853",
X"5b57fbad",
X"3f7555db",
X"3979841b",
X"83123354",
X"5b569839",
X"79841b71",
X"08575b56",
X"80547f53",
X"7c527d51",
X"fc9c3f87",
X"3976527d",
X"517c2d66",
X"70335881",
X"0547fd83",
X"39943d0d",
X"047283e0",
X"900c7183",
X"e0940c04",
X"fb3d0d88",
X"3d707084",
X"05520857",
X"54755383",
X"e0900852",
X"83e09408",
X"51fcc63f",
X"873d0d04",
X"ff3d0d73",
X"70085351",
X"02930533",
X"72347008",
X"8105710c",
X"833d0d04",
X"fc3d0d87",
X"3d881155",
X"785499b8",
X"5351fc99",
X"3f805287",
X"3d51d13f",
X"863d0d04",
X"fd3d0d75",
X"705254a3",
X"c23f83e0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83e0",
X"8008732e",
X"a13883e0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183e0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83e2c408",
X"248b3880",
X"cca53fff",
X"0b83e2c4",
X"0c800b83",
X"e0800c04",
X"ff3d0d73",
X"5283e0a0",
X"08722e8d",
X"38d83f71",
X"5196963f",
X"7183e0a0",
X"0c833d0d",
X"04f43d0d",
X"7e60625c",
X"5a558154",
X"bc150881",
X"92387451",
X"cf3f7958",
X"807a2580",
X"f83883e2",
X"f4087089",
X"2a5783ff",
X"06788480",
X"72315656",
X"57737825",
X"83387355",
X"7583e2c4",
X"082e8438",
X"ff883f83",
X"e2c40880",
X"25a63875",
X"892b5198",
X"d93f83e2",
X"f4088f3d",
X"fc11555c",
X"548152f8",
X"1b5196c3",
X"3f761483",
X"e2f40c75",
X"83e2c40c",
X"74537652",
X"785180ca",
X"b73f83e0",
X"800883e2",
X"f4081683",
X"e2f40c78",
X"7631761b",
X"5b595677",
X"8024ff8a",
X"38617a71",
X"0c547554",
X"75802e83",
X"38815473",
X"83e0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"993f7651",
X"feae3f86",
X"3dfc0553",
X"78527751",
X"95e53f79",
X"75710c54",
X"83e08008",
X"5483e080",
X"08802e83",
X"38815473",
X"83e0800c",
X"863d0d04",
X"fd3d0d76",
X"83e2c408",
X"53538072",
X"24893871",
X"732e8438",
X"fdd43f75",
X"51fde93f",
X"725197aa",
X"3f735273",
X"802e8338",
X"81527183",
X"e0800c85",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"e0800c51",
X"823d0d04",
X"80c40b83",
X"e0800c04",
X"fd3d0d75",
X"77715470",
X"5355539f",
X"9e3f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfcef3f",
X"735193ad",
X"3f7383e0",
X"a00c83e0",
X"80085383",
X"e0800880",
X"2e833881",
X"537283e0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcc33f",
X"72802ea5",
X"38bc1308",
X"5273519e",
X"a83f83e0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"e0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83e0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83e2c4",
X"0c7483e0",
X"a40c7583",
X"e2c00c80",
X"c7803f83",
X"e0800881",
X"ff065281",
X"53719938",
X"83e2dc51",
X"8e963f83",
X"e0800852",
X"83e08008",
X"802e8338",
X"72527153",
X"7283e080",
X"0c843d0d",
X"04fa3d0d",
X"787a82c4",
X"120882c4",
X"12087072",
X"24595656",
X"57577373",
X"2e098106",
X"913880c0",
X"165280c0",
X"17519c98",
X"3f83e080",
X"08557483",
X"e0800c88",
X"3d0d04f6",
X"3d0d7c5b",
X"807b715c",
X"54577a77",
X"2e8c3881",
X"1a82cc14",
X"08545a72",
X"f6388059",
X"80d9397a",
X"54815780",
X"707b7b31",
X"5a5755ff",
X"18537473",
X"2580c138",
X"82cc1408",
X"527351ff",
X"8c3f800b",
X"83e08008",
X"25a13882",
X"cc140882",
X"cc110882",
X"cc160c74",
X"82cc120c",
X"5375802e",
X"86387282",
X"cc170c72",
X"54805773",
X"82cc1508",
X"81175755",
X"56ffb839",
X"81195980",
X"0bff1b54",
X"54787325",
X"83388154",
X"76813270",
X"75065153",
X"72ff9038",
X"8c3d0d04",
X"f73d0d7b",
X"7d5a5a82",
X"d05283e2",
X"c0085180",
X"c6c83f83",
X"e0800857",
X"f9e43f79",
X"5283e2c8",
X"5195b63f",
X"83e08008",
X"54805383",
X"e0800873",
X"2e098106",
X"82833883",
X"e0a4080b",
X"0b80f1dc",
X"53705256",
X"9bd53f0b",
X"0b80f1dc",
X"5280c016",
X"519bc83f",
X"75bc170c",
X"7382c017",
X"0c810b82",
X"c4170c81",
X"0b82c817",
X"0c7382cc",
X"170cff17",
X"82d01755",
X"57819139",
X"83e0b033",
X"70822a70",
X"81065154",
X"55728180",
X"3874812a",
X"81065877",
X"80f63874",
X"842a8106",
X"82c4150c",
X"83e0b033",
X"810682c8",
X"150c7952",
X"73519aef",
X"3f73519b",
X"863f83e0",
X"80081453",
X"af737081",
X"05553472",
X"bc150c83",
X"e0b15272",
X"519ad03f",
X"83e0a808",
X"82c0150c",
X"83e0be52",
X"80c01451",
X"9abd3f78",
X"802e8d38",
X"7351782d",
X"83e08008",
X"802e9938",
X"7782cc15",
X"0c75802e",
X"86387382",
X"cc170c73",
X"82d015ff",
X"19595556",
X"76802e9b",
X"3883e0a8",
X"5283e2c8",
X"5194ac3f",
X"83e08008",
X"8a3883e0",
X"b1335372",
X"fed23878",
X"802e8938",
X"83e0a408",
X"51fcb83f",
X"83e0a408",
X"537283e0",
X"800c8b3d",
X"0d04ff3d",
X"0d805273",
X"51fdb53f",
X"833d0d04",
X"f03d0d62",
X"705254f6",
X"933f83e0",
X"80087453",
X"873d7053",
X"5555f6b3",
X"3ff7933f",
X"7351d33f",
X"63537452",
X"83e08008",
X"51fab73f",
X"923d0d04",
X"7183e080",
X"0c0480c0",
X"1283e080",
X"0c04803d",
X"0d7282c0",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"cc110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"82c41108",
X"83e0800c",
X"51823d0d",
X"04f93d0d",
X"7983e098",
X"08575781",
X"77278198",
X"38768817",
X"08278190",
X"38753355",
X"74822e89",
X"3874832e",
X"b4388180",
X"39745476",
X"1083fe06",
X"5376882a",
X"8c170805",
X"52893dfc",
X"055180c1",
X"9a3f83e0",
X"800880e0",
X"38029d05",
X"33893d33",
X"71882b07",
X"565680d2",
X"39845476",
X"822b83fc",
X"06537687",
X"2a8c1708",
X"0552893d",
X"fc055180",
X"c0e93f83",
X"e08008b0",
X"38029f05",
X"33028405",
X"9e053371",
X"982b7190",
X"2b07028c",
X"059d0533",
X"70882b72",
X"078d3d33",
X"7180ffff",
X"fe800607",
X"51525357",
X"58568339",
X"81557483",
X"e0800c89",
X"3d0d04fb",
X"3d0d83e0",
X"9808fe19",
X"881208fe",
X"05555654",
X"80567473",
X"278d3882",
X"14337571",
X"29941608",
X"05575375",
X"83e0800c",
X"873d0d04",
X"fc3d0d76",
X"52800b83",
X"e0980870",
X"33515253",
X"70832e09",
X"81069138",
X"95123394",
X"13337198",
X"2b71902b",
X"07555551",
X"9b12339a",
X"13337188",
X"2b077407",
X"83e0800c",
X"55863d0d",
X"04fc3d0d",
X"7683e098",
X"08555580",
X"75238815",
X"08537281",
X"2e883888",
X"14087326",
X"85388152",
X"b2397290",
X"38733352",
X"71832e09",
X"81068538",
X"90140853",
X"728c160c",
X"72802e8d",
X"387251fe",
X"d63f83e0",
X"80085285",
X"39901408",
X"52719016",
X"0c805271",
X"83e0800c",
X"863d0d04",
X"fa3d0d78",
X"83e09808",
X"71228105",
X"7083ffff",
X"06575457",
X"5573802e",
X"88389015",
X"08537286",
X"38835280",
X"e739738f",
X"06527180",
X"da388113",
X"90160c8c",
X"15085372",
X"9038830b",
X"84172257",
X"52737627",
X"80c638bf",
X"39821633",
X"ff057484",
X"2a065271",
X"b2387251",
X"fcaf3f81",
X"527183e0",
X"800827a8",
X"38835283",
X"e0800888",
X"1708279c",
X"3883e080",
X"088c160c",
X"83e08008",
X"51fdbc3f",
X"83e08008",
X"90160c73",
X"75238052",
X"7183e080",
X"0c883d0d",
X"04f23d0d",
X"60626458",
X"5e5b7533",
X"5574a02e",
X"09810688",
X"38811670",
X"4456ef39",
X"62703356",
X"5674af2e",
X"09810684",
X"38811643",
X"800b881c",
X"0c627033",
X"5155749f",
X"2691387a",
X"51fdd23f",
X"83e08008",
X"56807d34",
X"83813993",
X"3d841c08",
X"7058595f",
X"8a55a076",
X"70810558",
X"34ff1555",
X"74ff2e09",
X"8106ef38",
X"80705a5c",
X"887f085f",
X"5a7b811d",
X"7081ff06",
X"60137033",
X"70af3270",
X"30a07327",
X"71802507",
X"5151525b",
X"535e5755",
X"7480e738",
X"76ae2e09",
X"81068338",
X"8155787a",
X"27750755",
X"74802e9f",
X"38798832",
X"703078ae",
X"32703070",
X"73079f2a",
X"53515751",
X"5675bb38",
X"88598b5a",
X"ffab3976",
X"982b5574",
X"80258738",
X"80ef8c17",
X"3357ff9f",
X"17557499",
X"268938e0",
X"177081ff",
X"06585578",
X"811a7081",
X"ff06721b",
X"535b5755",
X"767534fe",
X"f8397b1e",
X"7f0c8055",
X"76a02683",
X"38815574",
X"8b19347a",
X"51fc823f",
X"83e08008",
X"80f538a0",
X"547a2270",
X"852b83e0",
X"06545590",
X"1b08527c",
X"51bba43f",
X"83e08008",
X"5783e080",
X"08818138",
X"7c335574",
X"802e80f4",
X"388b1d33",
X"70832a70",
X"81065156",
X"5674b438",
X"8b7d841d",
X"0883e080",
X"08595b5b",
X"58ff1858",
X"77ff2e9a",
X"38797081",
X"055b3379",
X"7081055b",
X"33717131",
X"52565675",
X"802ee238",
X"86397580",
X"2e96387a",
X"51fbe53f",
X"ff863983",
X"e0800856",
X"83e08008",
X"b6388339",
X"7656841b",
X"088b1133",
X"515574a7",
X"388b1d33",
X"70842a70",
X"81065156",
X"56748938",
X"83569439",
X"81569039",
X"7c51fa94",
X"3f83e080",
X"08881c0c",
X"fd813975",
X"83e0800c",
X"903d0d04",
X"f83d0d7a",
X"7c595782",
X"5483fe53",
X"77527651",
X"b9e93f83",
X"5683e080",
X"0880ec38",
X"81173377",
X"3371882b",
X"07565682",
X"567482d4",
X"d52e0981",
X"0680d438",
X"7554b653",
X"77527651",
X"b9bd3f83",
X"e0800898",
X"38811733",
X"77337188",
X"2b0783e0",
X"80085256",
X"56748182",
X"c62eac38",
X"825480d2",
X"53775276",
X"51b9943f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62e83",
X"38815675",
X"83e0800c",
X"8a3d0d04",
X"eb3d0d67",
X"5a800b83",
X"e0980cb8",
X"c93f83e0",
X"80088106",
X"55825674",
X"83ee3874",
X"75538f3d",
X"70535759",
X"feca3f83",
X"e0800881",
X"ff065776",
X"812e0981",
X"0680d438",
X"905483be",
X"53745275",
X"51b8a83f",
X"83e08008",
X"80c9388f",
X"3d335574",
X"802e80c9",
X"3802bf05",
X"33028405",
X"be053371",
X"982b7190",
X"2b07028c",
X"05bd0533",
X"70882b72",
X"07953d33",
X"71077058",
X"7b575e52",
X"5e575957",
X"fdee3f83",
X"e0800881",
X"ff065776",
X"832e0981",
X"06863881",
X"5682f139",
X"76802e86",
X"38865682",
X"e739a454",
X"8d537852",
X"7551b7bf",
X"3f815683",
X"e0800882",
X"d33802be",
X"05330284",
X"05bd0533",
X"71882b07",
X"595d77ab",
X"380280ce",
X"05330284",
X"0580cd05",
X"3371982b",
X"71902b07",
X"973d3370",
X"882b7207",
X"02940580",
X"cb053371",
X"0754525e",
X"57595602",
X"b7053378",
X"71290288",
X"05b60533",
X"028c05b5",
X"05337188",
X"2b07701d",
X"707f8c05",
X"0c5f5957",
X"595d8e3d",
X"33821b34",
X"02b90533",
X"903d3371",
X"882b075a",
X"5c78841b",
X"2302bb05",
X"33028405",
X"ba053371",
X"882b0756",
X"5c74ab38",
X"0280ca05",
X"33028405",
X"80c90533",
X"71982b71",
X"902b0796",
X"3d337088",
X"2b720702",
X"940580c7",
X"05337107",
X"51525357",
X"5e5c7476",
X"31783179",
X"842a903d",
X"33547171",
X"31535656",
X"b7ac3f83",
X"e0800882",
X"0570881c",
X"0c83e080",
X"08e08a05",
X"56567483",
X"dffe2683",
X"38825783",
X"fff67627",
X"85388357",
X"89398656",
X"76802e80",
X"db38767a",
X"3476832e",
X"098106b0",
X"380280d6",
X"05330284",
X"0580d505",
X"3371982b",
X"71902b07",
X"993d3370",
X"882b7207",
X"02940580",
X"d3053371",
X"077f9005",
X"0c525e57",
X"58568639",
X"771b901b",
X"0c841a22",
X"8c1b0819",
X"71842a05",
X"941c0c5d",
X"800b811b",
X"347983e0",
X"980c8056",
X"7583e080",
X"0c973d0d",
X"04e93d0d",
X"83e09808",
X"56855475",
X"802e8182",
X"38800b81",
X"1734993d",
X"e011466a",
X"548a3d70",
X"5458ec05",
X"51f6e63f",
X"83e08008",
X"5483e080",
X"0880df38",
X"893d3354",
X"73802e91",
X"3802ab05",
X"3370842a",
X"81065155",
X"74802e86",
X"38835480",
X"c1397651",
X"f48a3f83",
X"e08008a0",
X"170c02bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"3371079c",
X"1c0c5278",
X"981b0c53",
X"56595781",
X"0b811734",
X"74547383",
X"e0800c99",
X"3d0d04f5",
X"3d0d7d7f",
X"617283e0",
X"98085a5d",
X"5d595c80",
X"7b0c8557",
X"75802e81",
X"e0388116",
X"33810655",
X"84577480",
X"2e81d238",
X"91397481",
X"17348639",
X"800b8117",
X"34815781",
X"c0399c16",
X"08981708",
X"31557478",
X"27833874",
X"5877802e",
X"81a93898",
X"16087083",
X"ff065657",
X"7480cf38",
X"821633ff",
X"0577892a",
X"067081ff",
X"065a5578",
X"a0387687",
X"38a01608",
X"558d39a4",
X"160851f0",
X"e83f83e0",
X"80085581",
X"7527ffa8",
X"3874a417",
X"0ca41608",
X"51f2843f",
X"83e08008",
X"5583e080",
X"08802eff",
X"893883e0",
X"800819a8",
X"170c9816",
X"0883ff06",
X"84807131",
X"51557775",
X"27833877",
X"557483ff",
X"ff065498",
X"160883ff",
X"0653a816",
X"08527957",
X"7b83387b",
X"577651b1",
X"e63f83e0",
X"8008fed0",
X"38981608",
X"1598170c",
X"741a7876",
X"317c0817",
X"7d0c595a",
X"fed33980",
X"577683e0",
X"800c8d3d",
X"0d04fa3d",
X"0d7883e0",
X"98085556",
X"85557380",
X"2e81e138",
X"81143381",
X"06538455",
X"72802e81",
X"d3389c14",
X"08537276",
X"27833872",
X"56981408",
X"57800b98",
X"150c7580",
X"2e81b738",
X"82143370",
X"892b5653",
X"76802eb5",
X"387452ff",
X"1651b2ae",
X"3f83e080",
X"08ff1876",
X"54705358",
X"53b29f3f",
X"83e08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed73f83",
X"e0800853",
X"810b83e0",
X"8008278b",
X"38881408",
X"83e08008",
X"26883880",
X"0b811534",
X"b03983e0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc83f",
X"83e08008",
X"8c3883e0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683e0",
X"800805a8",
X"150c8055",
X"7483e080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83e09808",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1d23f",
X"83e08008",
X"5583e080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef8",
X"3f83e080",
X"0888170c",
X"7551efa9",
X"3f83e080",
X"08557483",
X"e0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683e0",
X"9808802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f83f83e0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"adf13f83",
X"e0800841",
X"83e08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"ede23f83",
X"e0800841",
X"83e08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"83a53f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f33f83e0",
X"80088332",
X"70307072",
X"079f2c83",
X"e0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"81b13f75",
X"83e0800c",
X"9e3d0d04",
X"fd3d0d75",
X"77535473",
X"33517089",
X"38713351",
X"70802ea1",
X"38733372",
X"33525372",
X"71278538",
X"ff519439",
X"70732785",
X"3881518b",
X"39811481",
X"135354d3",
X"39805170",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"77545472",
X"337081ff",
X"06525270",
X"802ea338",
X"7181ff06",
X"8114ffbf",
X"12535452",
X"70992689",
X"38a01270",
X"81ff0653",
X"51717470",
X"81055634",
X"d2398074",
X"34853d0d",
X"04ffbd3d",
X"0d80c63d",
X"0852a53d",
X"705254ff",
X"b33f80c7",
X"3d085285",
X"3d705253",
X"ffa63f72",
X"527351fe",
X"df3f80c5",
X"3d0d04fe",
X"3d0d7476",
X"53537170",
X"81055333",
X"51707370",
X"81055534",
X"70f03884",
X"3d0d04fe",
X"3d0d7452",
X"80723352",
X"5370732e",
X"8d388112",
X"81147133",
X"53545270",
X"f5387283",
X"e0800c84",
X"3d0d0471",
X"83e38c0c",
X"8880800b",
X"83e3880c",
X"8480800b",
X"83e3900c",
X"04f03d0d",
X"80f5c408",
X"54733383",
X"e3943483",
X"a0805683",
X"e38c0816",
X"83e38808",
X"17565474",
X"33743483",
X"e3900816",
X"54807434",
X"81165675",
X"83a0a02e",
X"098106db",
X"3883a480",
X"5683e38c",
X"081683e3",
X"88081756",
X"54743374",
X"3483e390",
X"08165480",
X"74348116",
X"567583a4",
X"a02e0981",
X"06db3883",
X"a8805683",
X"e38c0816",
X"83e38808",
X"17565474",
X"33743483",
X"e3900816",
X"54807434",
X"81165675",
X"83a8902e",
X"098106db",
X"3880f5c4",
X"0854ff74",
X"34805683",
X"e38c0816",
X"83e39008",
X"17555573",
X"33753481",
X"16567583",
X"a0802e09",
X"8106e438",
X"83b08056",
X"83e38c08",
X"1683e390",
X"08175555",
X"73337534",
X"81165675",
X"8480802e",
X"098106e4",
X"3886fd3f",
X"893d58a2",
X"5380f18c",
X"527751af",
X"8c3f8057",
X"8c805683",
X"e3900816",
X"77195555",
X"73337534",
X"81168118",
X"585676a2",
X"2e098106",
X"e63880f5",
X"e8085486",
X"743480f5",
X"ec085480",
X"743480f5",
X"e4085480",
X"743480f5",
X"d40854af",
X"743480f5",
X"e00854bf",
X"743480f5",
X"dc085480",
X"743480f5",
X"d808549f",
X"743480f5",
X"d0085480",
X"743480f5",
X"bc0854e0",
X"743480f5",
X"b4085476",
X"743480f5",
X"b0085483",
X"743480f5",
X"b8085482",
X"7434923d",
X"0d04fe3d",
X"0d805383",
X"e3900813",
X"83e38c08",
X"14525270",
X"33723481",
X"13537283",
X"a0802e09",
X"8106e438",
X"83b08053",
X"83e39008",
X"1383e38c",
X"08145252",
X"70337234",
X"81135372",
X"8480802e",
X"098106e4",
X"3883a080",
X"5383e390",
X"081383e3",
X"8c081452",
X"52703372",
X"34811353",
X"7283a0a0",
X"2e098106",
X"e43883a4",
X"805383e3",
X"90081383",
X"e38c0814",
X"52527033",
X"72348113",
X"537283a4",
X"a02e0981",
X"06e43883",
X"a8805383",
X"e3900813",
X"83e38c08",
X"14525270",
X"33723481",
X"13537283",
X"a8902e09",
X"8106e438",
X"80f5c408",
X"5183e394",
X"33713484",
X"3d0d0480",
X"3d0d80f6",
X"cc087008",
X"810683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d80f6",
X"cc087008",
X"70fe0676",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80f6cc08",
X"70087081",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80f6cc08",
X"700870fd",
X"06761007",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"f6cc0870",
X"0870822c",
X"bf0683e0",
X"800c5151",
X"823d0d04",
X"ff3d0d80",
X"f6cc0870",
X"0870fe83",
X"0676822b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80f6cc08",
X"70087088",
X"2c870683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80f6cc08",
X"700870f1",
X"ff067688",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d80f6cc",
X"08700870",
X"8b2cbf06",
X"83e0800c",
X"5151823d",
X"0d04ff3d",
X"0d80f6cc",
X"08700870",
X"f88fff06",
X"768b2b07",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"f6dc0870",
X"0870882c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"f6dc0870",
X"0870892c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"f6dc0870",
X"08708a2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"f6dc0870",
X"08708b2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"fd3d0d75",
X"81e62987",
X"2a80f6bc",
X"0854730c",
X"853d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d848080",
X"53805288",
X"800a51ff",
X"b33f8180",
X"80538052",
X"82800a51",
X"c63f843d",
X"0d04803d",
X"0d8151fc",
X"ce3f7280",
X"2e8338d2",
X"3f8151fc",
X"f03f8051",
X"fceb3f80",
X"51fcb83f",
X"823d0d04",
X"fd3d0d75",
X"52805480",
X"ff722588",
X"38810bff",
X"80135354",
X"ffbf1251",
X"70992686",
X"38e01252",
X"9e39ff9f",
X"12519971",
X"279538d0",
X"12e01370",
X"54545189",
X"71278838",
X"8f732783",
X"38805273",
X"802e8538",
X"81801252",
X"7181ff06",
X"83e0800c",
X"853d0d04",
X"803d0d84",
X"d8c05180",
X"71708105",
X"53347084",
X"e0c02e09",
X"8106f038",
X"823d0d04",
X"fe3d0d02",
X"97053351",
X"ff863f83",
X"e0800881",
X"ff0683e3",
X"98085452",
X"8073249b",
X"3883e3b4",
X"08137283",
X"e3b80807",
X"53537173",
X"3483e398",
X"08810583",
X"e3980c84",
X"3d0d04fa",
X"3d0d8280",
X"0a1b5580",
X"57883dfc",
X"05547953",
X"74527851",
X"d5ae3f88",
X"3d0d04fe",
X"3d0d83e3",
X"ac085274",
X"51dc8d3f",
X"83e08008",
X"8c387653",
X"755283e3",
X"ac0851c7",
X"3f843d0d",
X"04fe3d0d",
X"83e3ac08",
X"53755274",
X"51d6cb3f",
X"83e08008",
X"8d387753",
X"765283e3",
X"ac0851ff",
X"a23f843d",
X"0d04fe3d",
X"0d83e3b0",
X"0851d5bf",
X"3f83e080",
X"08818080",
X"2e098106",
X"883883c1",
X"8080539b",
X"3983e3b0",
X"0851d5a3",
X"3f83e080",
X"0880d080",
X"2e098106",
X"933883c1",
X"b0805383",
X"e0800852",
X"83e3b008",
X"51fed83f",
X"843d0d04",
X"803d0dfa",
X"cc3f83e0",
X"80088429",
X"80f3dc05",
X"700883e0",
X"800c5182",
X"3d0d04ee",
X"3d0d8043",
X"80428041",
X"80705a5b",
X"fdd23f80",
X"0b83e398",
X"0c800b83",
X"e3b80c80",
X"f2dc51d0",
X"933f8180",
X"0b83e3b8",
X"0c80f2e0",
X"51d0853f",
X"80d00b83",
X"e3980c78",
X"30707a07",
X"80257087",
X"2b83e3b8",
X"0c5155f9",
X"bb3f83e0",
X"80085280",
X"f2e851cf",
X"df3f80f8",
X"0b83e398",
X"0c788132",
X"70307072",
X"07802570",
X"872b83e3",
X"b80c5156",
X"56fef13f",
X"83e08008",
X"5280f2f4",
X"51cfb53f",
X"81a00b83",
X"e3980c78",
X"82327030",
X"70720780",
X"2570872b",
X"83e3b80c",
X"515683e3",
X"b0085256",
X"d0cf3f83",
X"e0800852",
X"80f2fc51",
X"cf863f81",
X"f00b83e3",
X"980c810b",
X"83e39c5b",
X"5883e398",
X"0882197a",
X"32703070",
X"72078025",
X"70872b83",
X"e3b80c51",
X"578e3d70",
X"55ff1b54",
X"57575798",
X"be3f7970",
X"84055b08",
X"51d0863f",
X"745483e0",
X"80085377",
X"5280f384",
X"51ceb93f",
X"a81783e3",
X"980c8118",
X"5877852e",
X"098106ff",
X"b0388390",
X"0b83e398",
X"0c788732",
X"70307072",
X"07802570",
X"872b83e3",
X"b80c5156",
X"80f39452",
X"56ce853f",
X"83e00b83",
X"e3980c78",
X"88327030",
X"70720780",
X"2570872b",
X"83e3b80c",
X"515680f3",
X"a85256cd",
X"e33f868d",
X"a051f9a0",
X"3f805291",
X"3d705255",
X"99b43f83",
X"52745199",
X"ad3f6119",
X"59788025",
X"85388059",
X"90398879",
X"25853888",
X"59873978",
X"882682b1",
X"3878822b",
X"5580f1b0",
X"150804f6",
X"f33f83e0",
X"80086157",
X"5575812e",
X"09810689",
X"3883e080",
X"08105590",
X"3975ff2e",
X"09810688",
X"3883e080",
X"08812c55",
X"90752585",
X"38905588",
X"39748024",
X"83388155",
X"7451f6d0",
X"3f81e639",
X"f6e33f83",
X"e0800861",
X"05557480",
X"25853880",
X"55883987",
X"75258338",
X"87557451",
X"f6df3f81",
X"c4396087",
X"3862802e",
X"81bb388a",
X"dd0b83e0",
X"9c0c83e3",
X"b00851ff",
X"bed53ffb",
X"8d3f81a5",
X"39605680",
X"76259938",
X"89f60b83",
X"e09c0c83",
X"e3901570",
X"085255ff",
X"beb53f74",
X"08529139",
X"75802591",
X"3883e390",
X"150851cd",
X"c63f8052",
X"fd1951b8",
X"3962802e",
X"80eb3883",
X"e3901570",
X"0883e39c",
X"08720c83",
X"e39c0cfd",
X"1a705351",
X"558ad53f",
X"83e08008",
X"5680518a",
X"cb3f83e0",
X"80085274",
X"5186e93f",
X"75528051",
X"86e23fb5",
X"3962802e",
X"b0388add",
X"0b83e09c",
X"0c83e3ac",
X"0851ffbd",
X"ca3f83e3",
X"ac0851cc",
X"d43f9c80",
X"0a5380c0",
X"805283e0",
X"800851f9",
X"a63f8155",
X"8c396287",
X"387a802e",
X"fad23880",
X"557483e0",
X"800c943d",
X"0d04fe3d",
X"0df5cd3f",
X"83e08008",
X"802e8638",
X"805180f7",
X"39f5d53f",
X"83e08008",
X"80eb38f5",
X"fb3f83e0",
X"8008802e",
X"aa388151",
X"f3cd3fef",
X"983f800b",
X"83e3980c",
X"fa813f83",
X"e0800853",
X"ff0b83e3",
X"980cf1ea",
X"3f72be38",
X"7251f3ab",
X"3fbc39f5",
X"af3f83e0",
X"8008802e",
X"b1388151",
X"f3993fee",
X"e43f89f6",
X"0b83e09c",
X"0c83e39c",
X"0851ffbc",
X"a63fff0b",
X"83e3980c",
X"f1b43f83",
X"e39c0852",
X"80518594",
X"3f8151f6",
X"993f843d",
X"0d04fc3d",
X"0d908080",
X"52868480",
X"8051cfa8",
X"3f83e080",
X"0880c338",
X"88df3f80",
X"f6e051d3",
X"e93f83e0",
X"800883e3",
X"b0085480",
X"f3b05383",
X"e0800852",
X"55cec33f",
X"83e08008",
X"8438f886",
X"3f9c800a",
X"5480c080",
X"5380f3bc",
X"527451f7",
X"d03f8151",
X"f5c03f92",
X"ea3f8151",
X"f5b83ffe",
X"913ffc39",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"0283e08c",
X"08fc050c",
X"800b83e3",
X"9c0b83e0",
X"8c08f805",
X"0c83e08c",
X"08f4050c",
X"cda23f83",
X"e0800886",
X"05fc0683",
X"e08c08f0",
X"050c0283",
X"e08c08f0",
X"0508310d",
X"833d7083",
X"e08c08f8",
X"05087084",
X"0583e08c",
X"08f8050c",
X"0c51c9ef",
X"3f83e08c",
X"08f40508",
X"810583e0",
X"8c08f405",
X"0c83e08c",
X"08f40508",
X"862e0981",
X"06ffad38",
X"86948080",
X"51ecbc3f",
X"ff0b83e3",
X"980c800b",
X"83e3b80c",
X"84d8c00b",
X"83e3b40c",
X"8151f0eb",
X"3f8151f1",
X"943f8051",
X"f18f3f81",
X"51f1b93f",
X"8151f296",
X"3f8251f1",
X"e03f80c6",
X"e0528051",
X"c7b33ffd",
X"dd3f83e0",
X"8c08fc05",
X"080d800b",
X"83e0800c",
X"873d0d83",
X"e08c0c04",
X"803d0d81",
X"ff51800b",
X"83e3c412",
X"34ff1151",
X"70f43882",
X"3d0d04ff",
X"3d0d7370",
X"33535181",
X"11337134",
X"71811234",
X"833d0d04",
X"fb3d0d77",
X"79565680",
X"70715555",
X"52717525",
X"ac387216",
X"70337014",
X"7081ff06",
X"55515151",
X"71742789",
X"38811270",
X"81ff0653",
X"51718114",
X"7083ffff",
X"06555254",
X"747324d6",
X"387183e0",
X"800c873d",
X"0d04fd3d",
X"0d7554c0",
X"dd3f83e0",
X"8008802e",
X"f63883e5",
X"e0088605",
X"7081ff06",
X"5253ffbe",
X"b53f8439",
X"fba03fc0",
X"bd3f83e0",
X"8008812e",
X"f338ffbf",
X"973f83e0",
X"80087434",
X"ffbf8d3f",
X"83e08008",
X"811534ff",
X"bf823f83",
X"e0800882",
X"1534ffbe",
X"f73f83e0",
X"80088315",
X"34ffbeec",
X"3f83e080",
X"08841534",
X"8439fada",
X"3fffbff6",
X"3f83e080",
X"08802ef2",
X"38733383",
X"e3c43481",
X"143383e3",
X"c5348214",
X"3383e3c6",
X"34831433",
X"83e3c734",
X"845283e3",
X"c451fea0",
X"3f83e080",
X"0881ff06",
X"84153355",
X"5372742e",
X"0981068d",
X"38ffbee6",
X"3f83e080",
X"08802e9a",
X"3883e5e0",
X"08a82e09",
X"81068938",
X"860b83e5",
X"e00c8739",
X"a80b83e5",
X"e00c80e4",
X"51f09d3f",
X"853d0d04",
X"f43d0d7e",
X"60595580",
X"5d807582",
X"2b7183e5",
X"e4120c83",
X"e5f8175b",
X"5b577679",
X"3477772e",
X"83b23876",
X"527751c8",
X"a73f8e3d",
X"fc055490",
X"5383e5cc",
X"527751c7",
X"e33f7c56",
X"75902e09",
X"81068390",
X"3883e5cc",
X"51fcfc3f",
X"83e5ce51",
X"fcf53f83",
X"e5d051fc",
X"ee3f7683",
X"e5dc0c77",
X"51c5ae3f",
X"80f1e452",
X"83e08008",
X"51ffb480",
X"3f83e080",
X"08812e09",
X"810680d3",
X"387683e5",
X"f40c820b",
X"83e5cc34",
X"ff960b83",
X"e5cd3477",
X"51c7f03f",
X"83e08008",
X"5583e080",
X"08772588",
X"3883e080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"e5ce3474",
X"83e5cf34",
X"7683e5d0",
X"34ff800b",
X"83e5d134",
X"818f3983",
X"e5cc3383",
X"e5cd3371",
X"882b0756",
X"5b7483ff",
X"ff2e0981",
X"0680e738",
X"fe800b83",
X"e5f40c81",
X"0b83e5dc",
X"0cff0b83",
X"e5cc34ff",
X"0b83e5cd",
X"347751c6",
X"fe3f83e0",
X"800883e5",
X"fc0c83e0",
X"80085583",
X"e0800880",
X"25883883",
X"e080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583e5ce",
X"347483e5",
X"cf347683",
X"e5d034ff",
X"800b83e5",
X"d134810b",
X"83e5db34",
X"a4397485",
X"962e0981",
X"0680fd38",
X"7583e5f4",
X"0c7751c6",
X"b33f83e5",
X"db3383e0",
X"80080755",
X"7483e5db",
X"3483e5db",
X"33810655",
X"74802e83",
X"38845783",
X"e5d03383",
X"e5d13371",
X"882b0756",
X"5c748180",
X"2e098106",
X"a13883e5",
X"ce3383e5",
X"cf337188",
X"2b07565b",
X"ad807527",
X"87387682",
X"07579c39",
X"76810757",
X"96397482",
X"802e0981",
X"06873876",
X"83075787",
X"397481ff",
X"268a3877",
X"83e5e41b",
X"0c767934",
X"8e3d0d04",
X"803d0d72",
X"842983e5",
X"e4057008",
X"83e0800c",
X"51823d0d",
X"04fe3d0d",
X"800b83e5",
X"c80c800b",
X"83e5c40c",
X"ff0b83e3",
X"c00ca80b",
X"83e5e00c",
X"ae51ffb8",
X"e93f800b",
X"83e5e454",
X"52807370",
X"8405550c",
X"81125271",
X"842e0981",
X"06ef3884",
X"3d0d04fe",
X"3d0d7402",
X"84059605",
X"22535371",
X"802e9738",
X"72708105",
X"543351ff",
X"b9873fff",
X"127083ff",
X"ff065152",
X"e639843d",
X"0d04fe3d",
X"0d029205",
X"225382ac",
X"51ebb53f",
X"80c351ff",
X"b8e33f81",
X"9651eba8",
X"3f725283",
X"e3c451ff",
X"b23f7252",
X"83e3c451",
X"f8da3f83",
X"e0800881",
X"ff0651ff",
X"b8bf3f84",
X"3d0d04ff",
X"b13d0d80",
X"d13df805",
X"51f9833f",
X"83e5c808",
X"810583e5",
X"c80c80cf",
X"3d33cf11",
X"7081ff06",
X"51565674",
X"832688ec",
X"38758f06",
X"ff055675",
X"83e3c008",
X"2e9b3875",
X"83269638",
X"7583e3c0",
X"0c758429",
X"83e5e405",
X"70085355",
X"7551fa9c",
X"3f807624",
X"88c83875",
X"842983e5",
X"e4055574",
X"08802e88",
X"b93883e3",
X"c0088429",
X"83e5e405",
X"70080288",
X"0582b905",
X"33525b55",
X"7480d22e",
X"84b03874",
X"80d22490",
X"3874bf2e",
X"9c387480",
X"d02e81d7",
X"3887f739",
X"7480d32e",
X"80d23874",
X"80d72e81",
X"c63887e6",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055656",
X"ffb7c03f",
X"80c151ff",
X"b6f33ff6",
X"d33f860b",
X"83e3c434",
X"815283e3",
X"c451ffb8",
X"ad3f8151",
X"fde43f74",
X"8938860b",
X"83e5e00c",
X"8739a80b",
X"83e5e00c",
X"ffb78c3f",
X"80c151ff",
X"b6bf3ff6",
X"9f3f900b",
X"83e5db33",
X"81065656",
X"74802e83",
X"38985683",
X"e5d03383",
X"e5d13371",
X"882b0756",
X"59748180",
X"2e098106",
X"9c3883e5",
X"ce3383e5",
X"cf337188",
X"2b075657",
X"ad807527",
X"8c387581",
X"80075685",
X"3975a007",
X"567583e3",
X"c434ff0b",
X"83e3c534",
X"e00b83e3",
X"c634800b",
X"83e3c734",
X"845283e3",
X"c451ffb7",
X"a13f8451",
X"869d3902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"5659ffb5",
X"fe3f7951",
X"c0fa3f83",
X"e0800880",
X"2e8b3880",
X"ce51ffb5",
X"a43f85f2",
X"3980c151",
X"ffb59a3f",
X"ffb6a13f",
X"ffb4a43f",
X"83e5f408",
X"58837525",
X"9b3883e5",
X"d03383e5",
X"d1337188",
X"2b07fc17",
X"71297a05",
X"8380055a",
X"51578d39",
X"74818029",
X"18ff8005",
X"58818057",
X"80567676",
X"2e9338ff",
X"b4f63f83",
X"e0800883",
X"e3c41734",
X"811656ea",
X"39ffb4e4",
X"3f83e080",
X"0881ff06",
X"775383e3",
X"c45256f4",
X"c33f83e0",
X"800881ff",
X"06557575",
X"2e098106",
X"818a38ff",
X"b4e53f80",
X"c151ffb4",
X"983fffb5",
X"9f3f7752",
X"7951ffbf",
X"8f3f805e",
X"80d13dfd",
X"f4055476",
X"5383e3c4",
X"527951ff",
X"bd9b3f02",
X"82b90533",
X"55815874",
X"80d72e09",
X"8106bd38",
X"80d13dfd",
X"f0055476",
X"538f3d70",
X"537a5259",
X"ffbea13f",
X"80567676",
X"2ea23875",
X"1983e3c4",
X"17337133",
X"70723270",
X"30708025",
X"70307e06",
X"811d5d5e",
X"51515152",
X"5b55db39",
X"82ac51e5",
X"ef3f7780",
X"2e863880",
X"c3518439",
X"80ce51ff",
X"b3933fff",
X"b49a3fff",
X"b29d3f83",
X"dd390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290559",
X"5580705d",
X"59ffb3b3",
X"3f80c151",
X"ffb2e63f",
X"83e5dc08",
X"792e82de",
X"3883e5fc",
X"0880fc05",
X"5580fd52",
X"74518896",
X"3f83e080",
X"085b7782",
X"24b238ff",
X"1870872b",
X"83ffff80",
X"0680f3fc",
X"0583e3c4",
X"59575581",
X"80557570",
X"81055733",
X"77708105",
X"5934ff15",
X"7081ff06",
X"515574ea",
X"38828d39",
X"7782e82e",
X"81ab3877",
X"82e92e09",
X"810681b2",
X"3880f3cc",
X"51ffb980",
X"3f785877",
X"87327030",
X"70720780",
X"257a8a32",
X"70307072",
X"07802573",
X"0753545a",
X"51575575",
X"802e9738",
X"78782692",
X"38a00b83",
X"e3c41a34",
X"81197081",
X"ff065a55",
X"eb398118",
X"7081ff06",
X"59558a78",
X"27ffbc38",
X"8f5883e3",
X"bf183383",
X"e3c41934",
X"ff187081",
X"ff065955",
X"778426ea",
X"38905880",
X"0b83e3c4",
X"19348118",
X"7081ff06",
X"70982b52",
X"59557480",
X"25e93880",
X"c6557a85",
X"8f248438",
X"80c25574",
X"83e3c434",
X"80f10b83",
X"e3c73481",
X"0b83e3c8",
X"347a83e3",
X"c5347a88",
X"2c557483",
X"e3c63480",
X"cb3982f0",
X"782580c4",
X"387780fd",
X"29fd97d3",
X"05527951",
X"ffbbbd3f",
X"80d13dfd",
X"ec055480",
X"fd5383e3",
X"c4527951",
X"ffbaf53f",
X"7b811959",
X"567580fc",
X"24833878",
X"5877882c",
X"557483e4",
X"c1347783",
X"e4c23475",
X"83e4c334",
X"81805980",
X"cc3983e5",
X"f4085783",
X"78259b38",
X"83e5d033",
X"83e5d133",
X"71882b07",
X"fc1a7129",
X"79058380",
X"05595159",
X"8d397781",
X"802917ff",
X"80055781",
X"80597652",
X"7951ffba",
X"cb3f80d1",
X"3dfdec05",
X"54785383",
X"e3c45279",
X"51ffba84",
X"3f7851f6",
X"b93fffb0",
X"b73fffae",
X"ba3f8b39",
X"83e5c408",
X"810583e5",
X"c40c80d1",
X"3d0d04f6",
X"da3febaa",
X"3ff939fc",
X"3d0d7678",
X"71842983",
X"e5e40570",
X"08515353",
X"53709e38",
X"80ce7234",
X"80cf0b81",
X"133480ce",
X"0b821334",
X"80c50b83",
X"13347084",
X"133480e7",
X"3983e5f8",
X"13335480",
X"d2723473",
X"822a7081",
X"06515180",
X"cf537084",
X"3880d753",
X"72811334",
X"a00b8213",
X"34738306",
X"5170812e",
X"9e387081",
X"24883870",
X"802e8f38",
X"9f397082",
X"2e923870",
X"832e9238",
X"933980d8",
X"558e3980",
X"d3558939",
X"80cd5584",
X"3980c455",
X"74831334",
X"80c40b84",
X"1334800b",
X"85133486",
X"3d0d04fd",
X"3d0d7554",
X"80740c80",
X"0b84150c",
X"800b8815",
X"0c80f5c8",
X"08703370",
X"81ff0670",
X"812a8132",
X"71813271",
X"81067181",
X"0631841a",
X"0c565670",
X"832a8132",
X"71822a81",
X"32718106",
X"71810631",
X"790c5255",
X"51515180",
X"f5c00870",
X"33700981",
X"0688170c",
X"5151853d",
X"0d04fe3d",
X"0d747654",
X"527151ff",
X"9a3f7281",
X"2ea23881",
X"73268d38",
X"72822eab",
X"3872832e",
X"9f38e639",
X"7108e238",
X"841208dd",
X"38881208",
X"d838a039",
X"88120881",
X"2e098106",
X"cc389439",
X"88120881",
X"2e8d3871",
X"08893884",
X"1208802e",
X"ffb73884",
X"3d0d04fd",
X"3d0d7554",
X"7383e684",
X"082ea738",
X"80f6c008",
X"74a00a07",
X"710c80f6",
X"d0085353",
X"71085170",
X"802ef938",
X"80730c71",
X"085170fb",
X"387383e6",
X"840c853d",
X"0d04ff0b",
X"83e6840c",
X"8180800b",
X"83e6800c",
X"800b83e0",
X"800c04fc",
X"3d0d7602",
X"8405a205",
X"22028805",
X"a605227a",
X"54555555",
X"ff9d3f72",
X"802ea338",
X"83e68008",
X"14527133",
X"75708105",
X"57348114",
X"7083ffff",
X"06ff1570",
X"83ffff06",
X"56525552",
X"da39800b",
X"83e0800c",
X"863d0d04",
X"f73d0d7b",
X"7d7f1158",
X"55598055",
X"73762eb1",
X"3883e680",
X"088b3d59",
X"57741970",
X"3375fc06",
X"1970085d",
X"7683067b",
X"07535454",
X"51727134",
X"79720c81",
X"14811656",
X"5473762e",
X"098106d9",
X"38800b83",
X"e0800c8b",
X"3d0d04fe",
X"3d0d80f6",
X"c00883e6",
X"8408900a",
X"07710c80",
X"f6d00853",
X"53710851",
X"70802ef9",
X"3880730c",
X"71085170",
X"fb38843d",
X"0d0483e0",
X"8c080283",
X"e08c0cfd",
X"3d0d8053",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"83d43f83",
X"e0800870",
X"83e0800c",
X"54853d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cfd3d",
X"0d815383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"05085183",
X"a13f83e0",
X"80087083",
X"e0800c54",
X"853d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cf93d0d",
X"800b83e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"8025b938",
X"83e08c08",
X"88050830",
X"83e08c08",
X"88050c80",
X"0b83e08c",
X"08f4050c",
X"83e08c08",
X"fc05088a",
X"38810b83",
X"e08c08f4",
X"050c83e0",
X"8c08f405",
X"0883e08c",
X"08fc050c",
X"83e08c08",
X"8c050880",
X"25b93883",
X"e08c088c",
X"05083083",
X"e08c088c",
X"050c800b",
X"83e08c08",
X"f0050c83",
X"e08c08fc",
X"05088a38",
X"810b83e0",
X"8c08f005",
X"0c83e08c",
X"08f00508",
X"83e08c08",
X"fc050c80",
X"5383e08c",
X"088c0508",
X"5283e08c",
X"08880508",
X"5181df3f",
X"83e08008",
X"7083e08c",
X"08f8050c",
X"5483e08c",
X"08fc0508",
X"802e9038",
X"83e08c08",
X"f8050830",
X"83e08c08",
X"f8050c83",
X"e08c08f8",
X"05087083",
X"e0800c54",
X"893d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"800b83e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"80259938",
X"83e08c08",
X"88050830",
X"83e08c08",
X"88050c81",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"8c050880",
X"25903883",
X"e08c088c",
X"05083083",
X"e08c088c",
X"050c8153",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"bd3f83e0",
X"80087083",
X"e08c08f8",
X"050c5483",
X"e08c08fc",
X"0508802e",
X"903883e0",
X"8c08f805",
X"083083e0",
X"8c08f805",
X"0c83e08c",
X"08f80508",
X"7083e080",
X"0c54873d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cfd",
X"3d0d810b",
X"83e08c08",
X"fc050c80",
X"0b83e08c",
X"08f8050c",
X"83e08c08",
X"8c050883",
X"e08c0888",
X"050827b9",
X"3883e08c",
X"08fc0508",
X"802eae38",
X"800b83e0",
X"8c088c05",
X"0824a238",
X"83e08c08",
X"8c050810",
X"83e08c08",
X"8c050c83",
X"e08c08fc",
X"05081083",
X"e08c08fc",
X"050cffb8",
X"3983e08c",
X"08fc0508",
X"802e80e1",
X"3883e08c",
X"088c0508",
X"83e08c08",
X"88050826",
X"ad3883e0",
X"8c088805",
X"0883e08c",
X"088c0508",
X"3183e08c",
X"0888050c",
X"83e08c08",
X"f8050883",
X"e08c08fc",
X"05080783",
X"e08c08f8",
X"050c83e0",
X"8c08fc05",
X"08812a83",
X"e08c08fc",
X"050c83e0",
X"8c088c05",
X"08812a83",
X"e08c088c",
X"050cff95",
X"3983e08c",
X"08900508",
X"802e9338",
X"83e08c08",
X"88050870",
X"83e08c08",
X"f4050c51",
X"913983e0",
X"8c08f805",
X"087083e0",
X"8c08f405",
X"0c5183e0",
X"8c08f405",
X"0883e080",
X"0c853d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cff3d",
X"0d800b83",
X"e08c08fc",
X"050c83e0",
X"8c088805",
X"088106ff",
X"11700970",
X"83e08c08",
X"8c050806",
X"83e08c08",
X"fc050811",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"0508812a",
X"83e08c08",
X"88050c83",
X"e08c088c",
X"05081083",
X"e08c088c",
X"050c5151",
X"515183e0",
X"8c088805",
X"08802e84",
X"38ffab39",
X"83e08c08",
X"fc050870",
X"83e0800c",
X"51833d0d",
X"83e08c0c",
X"04fc3d0d",
X"7670797b",
X"55555555",
X"8f72278c",
X"38727507",
X"83065170",
X"802ea938",
X"ff125271",
X"ff2e9838",
X"72708105",
X"54337470",
X"81055634",
X"ff125271",
X"ff2e0981",
X"06ea3874",
X"83e0800c",
X"863d0d04",
X"74517270",
X"84055408",
X"71708405",
X"530c7270",
X"84055408",
X"71708405",
X"530c7270",
X"84055408",
X"71708405",
X"530c7270",
X"84055408",
X"71708405",
X"530cf012",
X"52718f26",
X"c9388372",
X"27953872",
X"70840554",
X"08717084",
X"05530cfc",
X"12527183",
X"26ed3870",
X"54ff8139",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"000025f3",
X"00002634",
X"00002656",
X"00002675",
X"00002675",
X"00002675",
X"00002675",
X"000026e5",
X"00002716",
X"25732025",
X"73000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"524f4d00",
X"42494e00",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"43617274",
X"72696467",
X"6520386b",
X"2073696d",
X"706c6500",
X"45786974",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"6e616d65",
X"20000000",
X"00000000",
X"00000000",
X"00003918",
X"0000391c",
X"00003924",
X"00003930",
X"0000393c",
X"00003948",
X"00003954",
X"00003958",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"0001d20f",
X"0001d400",
X"0001d401",
X"0001d409",
X"0001d010",
X"0001d301",
X"0001d300",
X"0001d20a",
X"0001d01b",
X"0001d016",
X"0001d019",
X"0001d018",
X"0001d017",
X"0001d01a",
X"0001d403",
X"0001d402",
X"0001d40e",
X"0004007c",
X"00040078",
X"00040074",
X"00040068",
X"00040060",
X"0004005c",
X"00040058",
X"00040054",
X"00040050",
X"0004004c",
X"00040048",
X"00040044",
X"00040040",
X"00040034",
X"00040030",
X"0004002c",
X"00040028",
X"00040024",
X"00040020",
X"0004001c",
X"00040018",
X"00040014",
X"00040010",
X"0004000c",
X"00040008",
X"00040004",
X"00040000",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
