
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f7",
X"f8738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80fb",
X"b00c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f3",
X"c32d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580f1d7",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80dbb204",
X"f23d0d60",
X"913dec11",
X"56565990",
X"53f01552",
X"7851948a",
X"3f83e080",
X"0880e538",
X"7a902e09",
X"810680dc",
X"3802b305",
X"3380fbb8",
X"0b80fbb8",
X"33575757",
X"8c397477",
X"2e8a3884",
X"16703356",
X"5674f338",
X"75337058",
X"5574802e",
X"80cf3880",
X"0b821722",
X"70832a57",
X"58587775",
X"27bb3896",
X"800a5790",
X"3dec0554",
X"80c08053",
X"76527851",
X"93ac3f83",
X"e0800888",
X"387a80c0",
X"802e8538",
X"80579a39",
X"811880c0",
X"80188218",
X"2270832a",
X"585c5858",
X"747826cb",
X"38811633",
X"577683e0",
X"800c903d",
X"0d04fc3d",
X"0d767052",
X"55b3c93f",
X"83e08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"811451b2",
X"e13f83e0",
X"80083070",
X"83e08008",
X"07802583",
X"e0800c53",
X"863d0d04",
X"fc3d0d76",
X"7052559a",
X"823f83e0",
X"80085481",
X"5383e080",
X"0880c738",
X"745199c5",
X"3f83e080",
X"080b0b80",
X"f9b85383",
X"e0800852",
X"53ff8f3f",
X"83e08008",
X"a5380b0b",
X"80f9bc52",
X"7251fefe",
X"3f83e080",
X"0894380b",
X"0b80f9c0",
X"527251fe",
X"ed3f83e0",
X"8008802e",
X"83388154",
X"73537283",
X"e0800c86",
X"3d0d04fd",
X"3d0d7570",
X"5254999b",
X"3f815383",
X"e0800898",
X"38735198",
X"e43f83e0",
X"a0085283",
X"e0800851",
X"feb43f83",
X"e0800853",
X"7283e080",
X"0c853d0d",
X"04e03d0d",
X"a33d0870",
X"525e8f89",
X"3f83e080",
X"0833943d",
X"56547394",
X"3880ffec",
X"52745184",
X"c7397d52",
X"7851928c",
X"3f84d139",
X"7d518ef1",
X"3f83e080",
X"08527451",
X"8ea13f83",
X"e0a80852",
X"933d7052",
X"5d94fc3f",
X"83e08008",
X"59800b83",
X"e0800855",
X"5b83e080",
X"087b2e94",
X"38811b74",
X"525b97fe",
X"3f83e080",
X"085483e0",
X"8008ee38",
X"805aff7a",
X"437a427a",
X"415f7909",
X"709f2c7b",
X"065b547a",
X"7a248438",
X"ff1b5af6",
X"1a700970",
X"9f2c7206",
X"7bff125a",
X"5a525555",
X"80752595",
X"38765197",
X"bd3f83e0",
X"800876ff",
X"18585557",
X"738024ed",
X"38747f2e",
X"873880c3",
X"a13f745f",
X"78ff1b70",
X"585d5880",
X"7a259538",
X"77519792",
X"3f83e080",
X"0876ff18",
X"58555873",
X"8024ed38",
X"800b83e7",
X"bc0c800b",
X"83e7dc0c",
X"0b0b80f9",
X"c4518be4",
X"3f81800b",
X"83e7dc0c",
X"0b0b80f9",
X"cc518bd4",
X"3fa80b83",
X"e7bc0c76",
X"802e80e8",
X"3883e7bc",
X"08777932",
X"70307072",
X"07802570",
X"872b83e7",
X"dc0c5156",
X"78535656",
X"96c53f83",
X"e0800880",
X"2e8a380b",
X"0b80f9d4",
X"518b993f",
X"76519685",
X"3f83e080",
X"08520b0b",
X"80fae051",
X"8b863f76",
X"51968b3f",
X"83e08008",
X"83e7bc08",
X"55577574",
X"258638a8",
X"1656f739",
X"7583e7bc",
X"0c86f076",
X"24ff9438",
X"87980b83",
X"e7bc0c77",
X"802eb738",
X"775195c1",
X"3f83e080",
X"08785255",
X"95e13f0b",
X"0b80f9dc",
X"5483e080",
X"088f3887",
X"39807634",
X"fd95390b",
X"0b80f9d8",
X"54745373",
X"520b0b80",
X"f9ac518a",
X"9f3f8054",
X"0b0b80fb",
X"ac518a94",
X"3f811454",
X"73a82e09",
X"8106ed38",
X"868da051",
X"bfa03f80",
X"52903d70",
X"525480e0",
X"873f8352",
X"735180df",
X"ff3f6180",
X"2e80ff38",
X"7b5473ff",
X"2e963878",
X"802e8180",
X"38785194",
X"e13f83e0",
X"8008ff15",
X"5559e739",
X"78802e80",
X"eb387851",
X"94dd3f83",
X"e0800880",
X"2efc8338",
X"785194a5",
X"3f83e080",
X"08520b0b",
X"80f9b451",
X"ac833f83",
X"e08008a4",
X"387c51ad",
X"bb3f83e0",
X"80085574",
X"ff165654",
X"807425fb",
X"ee38741d",
X"70335556",
X"73af2efe",
X"c838e839",
X"785193e3",
X"3f83e080",
X"08527c51",
X"acf23ffb",
X"ce397f88",
X"29601005",
X"7a056105",
X"5afbff39",
X"a23d0d04",
X"fe3d0d80",
X"feec0870",
X"337081ff",
X"0670842a",
X"81328106",
X"55515253",
X"71802e8c",
X"38a87334",
X"80feec08",
X"51b87134",
X"7183e080",
X"0c843d0d",
X"04fe3d0d",
X"80feec08",
X"70337081",
X"ff067085",
X"2a813281",
X"06555152",
X"5371802e",
X"8c389873",
X"3480feec",
X"0851b871",
X"347183e0",
X"800c843d",
X"0d04803d",
X"0d80fee8",
X"08519371",
X"3480fef4",
X"0851ff71",
X"34823d0d",
X"04fe3d0d",
X"02930533",
X"80fee808",
X"53538072",
X"348a51bc",
X"e93fd33f",
X"80fef808",
X"5280f872",
X"3480ff90",
X"08528072",
X"34fa1380",
X"ff980853",
X"53727234",
X"80ff8008",
X"52807234",
X"80ff8808",
X"52727234",
X"80feec08",
X"52807234",
X"80feec08",
X"52b87234",
X"843d0d04",
X"ff3d0d02",
X"8f053380",
X"fef00852",
X"52717134",
X"fe9e3f83",
X"e0800880",
X"2ef63883",
X"3d0d0480",
X"3d0d8539",
X"80c6953f",
X"feb73f83",
X"e0800880",
X"2ef23880",
X"fef00870",
X"337081ff",
X"0683e080",
X"0c515182",
X"3d0d0480",
X"3d0d80fe",
X"e80851a3",
X"713480fe",
X"f40851ff",
X"713480fe",
X"ec0851a8",
X"713480fe",
X"ec0851b8",
X"7134823d",
X"0d04803d",
X"0d80fee8",
X"08703370",
X"81c00670",
X"30708025",
X"83e0800c",
X"51515151",
X"823d0d04",
X"ff3d0d80",
X"feec0870",
X"337081ff",
X"0670832a",
X"81327081",
X"06515151",
X"52527080",
X"2ee538b0",
X"723480fe",
X"ec0851b8",
X"7134833d",
X"0d04803d",
X"0d80ffa4",
X"08700881",
X"0683e080",
X"0c51823d",
X"0d04fd3d",
X"0d757754",
X"54807325",
X"94387370",
X"81055533",
X"5280f9e0",
X"5185a13f",
X"ff1353e9",
X"39853d0d",
X"04f63d0d",
X"7c7e6062",
X"5a5d5b56",
X"80598155",
X"8539747a",
X"29557452",
X"755180db",
X"e03f83e0",
X"80087a27",
X"ed387480",
X"2e80e038",
X"74527551",
X"80dbca3f",
X"83e08008",
X"75537652",
X"5480dbf0",
X"3f83e080",
X"087a5375",
X"525680db",
X"b03f83e0",
X"80087930",
X"707b079f",
X"2a707780",
X"24075151",
X"54557287",
X"3883e080",
X"08c23876",
X"8118b016",
X"55585889",
X"74258b38",
X"b714537a",
X"853880d7",
X"14537278",
X"34811959",
X"ff9c3980",
X"77348c3d",
X"0d04f73d",
X"0d7b7d7f",
X"62029005",
X"bb053357",
X"59565a5a",
X"b0587283",
X"38a05875",
X"70708105",
X"52337159",
X"54559039",
X"8074258e",
X"38ff1477",
X"70810559",
X"33545472",
X"ef3873ff",
X"15555380",
X"73258938",
X"77527951",
X"782def39",
X"75337557",
X"5372802e",
X"90387252",
X"7951782d",
X"75708105",
X"573353ed",
X"398b3d0d",
X"04ee3d0d",
X"64666969",
X"70708105",
X"52335b4a",
X"5c5e5e76",
X"802e82f9",
X"3876a52e",
X"09810682",
X"e0388070",
X"41677070",
X"81055233",
X"714a5957",
X"5f76b02e",
X"0981068c",
X"38757081",
X"05573376",
X"4857815f",
X"d0175675",
X"892680da",
X"3876675c",
X"59805c93",
X"39778a24",
X"80c3387b",
X"8a29187b",
X"7081055d",
X"335a5cd0",
X"197081ff",
X"06585889",
X"7727a438",
X"ff9f1970",
X"81ff06ff",
X"a91b5a51",
X"56857627",
X"9238ffbf",
X"197081ff",
X"06515675",
X"85268a38",
X"c9195877",
X"8025ffb9",
X"387a477b",
X"407881ff",
X"06577680",
X"e42e80e5",
X"387680e4",
X"24a73876",
X"80d82e81",
X"86387680",
X"d8249038",
X"76802e81",
X"cc3876a5",
X"2e81b638",
X"81b93976",
X"80e32e81",
X"8c3881af",
X"397680f5",
X"2e9b3876",
X"80f5248b",
X"387680f3",
X"2e818138",
X"81993976",
X"80f82e80",
X"ca38818f",
X"39913d70",
X"55578053",
X"8a527984",
X"1b710853",
X"5b56fbfd",
X"3f7655ab",
X"3979841b",
X"7108943d",
X"705b5b52",
X"5b567580",
X"258c3875",
X"3056ad78",
X"340280c1",
X"05577654",
X"80538a52",
X"7551fbd1",
X"3f77557e",
X"54b83991",
X"3d705577",
X"80d83270",
X"30708025",
X"56515856",
X"90527984",
X"1b710853",
X"5b57fbad",
X"3f7555db",
X"3979841b",
X"83123354",
X"5b569839",
X"79841b71",
X"08575b56",
X"80547f53",
X"7c527d51",
X"fc9c3f87",
X"3976527d",
X"517c2d66",
X"70335881",
X"0547fd83",
X"39943d0d",
X"047283e0",
X"900c7183",
X"e0940c04",
X"fb3d0d88",
X"3d707084",
X"05520857",
X"54755383",
X"e0900852",
X"83e09408",
X"51fcc63f",
X"873d0d04",
X"ff3d0d73",
X"70085351",
X"02930533",
X"72347008",
X"8105710c",
X"833d0d04",
X"fc3d0d87",
X"3d881155",
X"78549aac",
X"5351fc99",
X"3f805287",
X"3d51d13f",
X"863d0d04",
X"fd3d0d75",
X"705254a3",
X"c33f83e0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83e0",
X"8008732e",
X"a13883e0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183e0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83e2d408",
X"248a38a4",
X"ad3fff0b",
X"83e2d40c",
X"800b83e0",
X"800c04ff",
X"3d0d7352",
X"83e0b008",
X"722e8d38",
X"d93f7151",
X"96983f71",
X"83e0b00c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"558154bc",
X"15088191",
X"387451cf",
X"3f795880",
X"7a2580f7",
X"3883e384",
X"0870892a",
X"5783ff06",
X"78848072",
X"31565657",
X"73782583",
X"38735575",
X"83e2d408",
X"2e8438ff",
X"893f83e2",
X"d4088025",
X"a6387589",
X"2b5198db",
X"3f83e384",
X"088f3dfc",
X"11555c54",
X"8152f81b",
X"5196c53f",
X"761483e3",
X"840c7583",
X"e2d40c74",
X"53765278",
X"51a2de3f",
X"83e08008",
X"83e38408",
X"1683e384",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8b3861",
X"7a710c54",
X"75547580",
X"2e833881",
X"547383e0",
X"800c8e3d",
X"0d04fc3d",
X"0dfe9b3f",
X"7651feaf",
X"3f863dfc",
X"05537852",
X"775195e8",
X"3f797571",
X"0c5483e0",
X"80085483",
X"e0800880",
X"2e833881",
X"547383e0",
X"800c863d",
X"0d04fe3d",
X"0d7583e2",
X"d4085353",
X"80722489",
X"3871732e",
X"8438fdd6",
X"3f7451fd",
X"ea3f7251",
X"97ad3f83",
X"e0800852",
X"83e08008",
X"802e8338",
X"81527183",
X"e0800c84",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"e0800c51",
X"823d0d04",
X"80c40b83",
X"e0800c04",
X"fd3d0d75",
X"77715470",
X"5355539f",
X"9b3f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfceb3f",
X"735193aa",
X"3f7383e0",
X"b00c83e0",
X"80085383",
X"e0800880",
X"2e833881",
X"537283e0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcbf3f",
X"72802ea5",
X"38bc1308",
X"5273519e",
X"a53f83e0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"e0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83e0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83e2d4",
X"0c7483e0",
X"b40c7583",
X"e2d00c9f",
X"923f83e0",
X"800881ff",
X"06528153",
X"71993883",
X"e2ec518e",
X"943f83e0",
X"80085283",
X"e0800880",
X"2e833872",
X"52715372",
X"83e0800c",
X"843d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"519c963f",
X"83e08008",
X"557483e0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"e0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283e2d0",
X"085180ce",
X"e83f83e0",
X"800857f9",
X"e13f7952",
X"83e2d851",
X"95b43f83",
X"e0800854",
X"805383e0",
X"8008732e",
X"09810682",
X"833883e0",
X"b4080b0b",
X"80f9b453",
X"7052569b",
X"d33f0b0b",
X"80f9b452",
X"80c01651",
X"9bc63f75",
X"bc170c73",
X"82c0170c",
X"810b82c4",
X"170c810b",
X"82c8170c",
X"7382cc17",
X"0cff1782",
X"d0175557",
X"81913983",
X"e0c03370",
X"822a7081",
X"06515455",
X"72818038",
X"74812a81",
X"06587780",
X"f6387484",
X"2a810682",
X"c4150c83",
X"e0c03381",
X"0682c815",
X"0c795273",
X"519aed3f",
X"73519b84",
X"3f83e080",
X"081453af",
X"73708105",
X"553472bc",
X"150c83e0",
X"c1527251",
X"9ace3f83",
X"e0b80882",
X"c0150c83",
X"e0ce5280",
X"c014519a",
X"bb3f7880",
X"2e8d3873",
X"51782d83",
X"e0800880",
X"2e993877",
X"82cc150c",
X"75802e86",
X"387382cc",
X"170c7382",
X"d015ff19",
X"59555676",
X"802e9b38",
X"83e0b852",
X"83e2d851",
X"94aa3f83",
X"e080088a",
X"3883e0c1",
X"335372fe",
X"d2387880",
X"2e893883",
X"e0b40851",
X"fcb83f83",
X"e0b40853",
X"7283e080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb53f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f690",
X"3f83e080",
X"08745387",
X"3d705355",
X"55f6b03f",
X"f7903f73",
X"51d33f63",
X"53745283",
X"e0800851",
X"fab83f92",
X"3d0d0471",
X"83e0800c",
X"0480c012",
X"83e0800c",
X"04803d0d",
X"7282c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"e0800c51",
X"823d0d04",
X"f93d0d79",
X"83e09808",
X"57578177",
X"27819638",
X"76881708",
X"27818e38",
X"75335574",
X"822e8938",
X"74832eb3",
X"3880fe39",
X"74547610",
X"83fe0653",
X"76882a8c",
X"17080552",
X"893dfc05",
X"5199c03f",
X"83e08008",
X"80df3802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d13984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"5199903f",
X"83e08008",
X"b038029f",
X"05330284",
X"059e0533",
X"71982b71",
X"902b0702",
X"8c059d05",
X"3370882b",
X"72078d3d",
X"337180ff",
X"fffe8006",
X"07515253",
X"57585683",
X"39815574",
X"83e0800c",
X"893d0d04",
X"fb3d0d83",
X"e09808fe",
X"19881208",
X"fe055556",
X"54805674",
X"73278d38",
X"82143375",
X"71299416",
X"08055753",
X"7583e080",
X"0c873d0d",
X"04fc3d0d",
X"7652800b",
X"83e09808",
X"70335152",
X"5370832e",
X"09810691",
X"38951233",
X"94133371",
X"982b7190",
X"2b075555",
X"519b1233",
X"9a133371",
X"882b0774",
X"0783e080",
X"0c55863d",
X"0d04fc3d",
X"0d7683e0",
X"98085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"fed63f83",
X"e0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183e080",
X"0c863d0d",
X"04fa3d0d",
X"7883e098",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fcb13f",
X"81527183",
X"e0800827",
X"a8388352",
X"83e08008",
X"88170827",
X"9c3883e0",
X"80088c16",
X"0c83e080",
X"0851fdbc",
X"3f83e080",
X"0890160c",
X"73752380",
X"527183e0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585e5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"9f269138",
X"7a51fdd2",
X"3f83e080",
X"0856807d",
X"34838139",
X"933d841c",
X"08705859",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"3880705a",
X"5c887f08",
X"5f5a7b81",
X"1d7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535e57",
X"557480e7",
X"3876ae2e",
X"09810683",
X"38815578",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675bb",
X"3888598b",
X"5affab39",
X"76982b55",
X"74802587",
X"3880f788",
X"173357ff",
X"9f175574",
X"99268938",
X"e0177081",
X"ff065855",
X"78811a70",
X"81ff0672",
X"1b535b57",
X"55767534",
X"fef8397b",
X"1e7f0c80",
X"5576a026",
X"83388155",
X"748b1934",
X"7a51fc82",
X"3f83e080",
X"0880f538",
X"a0547a22",
X"70852b83",
X"e0065455",
X"901b0852",
X"7c5193cb",
X"3f83e080",
X"085783e0",
X"80088181",
X"387c3355",
X"74802e80",
X"f4388b1d",
X"3370832a",
X"70810651",
X"565674b4",
X"388b7d84",
X"1d0883e0",
X"8008595b",
X"5b58ff18",
X"5877ff2e",
X"9a387970",
X"81055b33",
X"79708105",
X"5b337171",
X"31525656",
X"75802ee2",
X"38863975",
X"802e9638",
X"7a51fbe5",
X"3fff8639",
X"83e08008",
X"5683e080",
X"08b63883",
X"39765684",
X"1b088b11",
X"33515574",
X"a7388b1d",
X"3370842a",
X"70810651",
X"56567489",
X"38835694",
X"39815690",
X"397c51fa",
X"943f83e0",
X"8008881c",
X"0cfd8139",
X"7583e080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"5192903f",
X"835683e0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"5191e43f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"765191bb",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583e080",
X"0c8a3d0d",
X"04eb3d0d",
X"675a800b",
X"83e0980c",
X"90dd3f83",
X"e0800881",
X"06558256",
X"7483ee38",
X"7475538f",
X"3d705357",
X"59feca3f",
X"83e08008",
X"81ff0657",
X"76812e09",
X"810680d4",
X"38905483",
X"be537452",
X"755190cf",
X"3f83e080",
X"0880c938",
X"8f3d3355",
X"74802e80",
X"c93802bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"33710770",
X"587b575e",
X"525e5759",
X"57fdee3f",
X"83e08008",
X"81ff0657",
X"76832e09",
X"81068638",
X"815682f1",
X"3976802e",
X"86388656",
X"82e739a4",
X"548d5378",
X"5275518f",
X"e63f8156",
X"83e08008",
X"82d33802",
X"be053302",
X"8405bd05",
X"3371882b",
X"07595d77",
X"ab380280",
X"ce053302",
X"840580cd",
X"05337198",
X"2b71902b",
X"07973d33",
X"70882b72",
X"07029405",
X"80cb0533",
X"71075452",
X"5e575956",
X"02b70533",
X"78712902",
X"8805b605",
X"33028c05",
X"b5053371",
X"882b0770",
X"1d707f8c",
X"050c5f59",
X"57595d8e",
X"3d33821b",
X"3402b905",
X"33903d33",
X"71882b07",
X"5a5c7884",
X"1b2302bb",
X"05330284",
X"05ba0533",
X"71882b07",
X"565c74ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"07515253",
X"575e5c74",
X"76317831",
X"79842a90",
X"3d335471",
X"71315356",
X"56bfce3f",
X"83e08008",
X"82057088",
X"1c0c83e0",
X"8008e08a",
X"05565674",
X"83dffe26",
X"83388257",
X"83fff676",
X"27853883",
X"57893986",
X"5676802e",
X"80db3876",
X"7a347683",
X"2e098106",
X"b0380280",
X"d6053302",
X"840580d5",
X"05337198",
X"2b71902b",
X"07993d33",
X"70882b72",
X"07029405",
X"80d30533",
X"71077f90",
X"050c525e",
X"57585686",
X"39771b90",
X"1b0c841a",
X"228c1b08",
X"1971842a",
X"05941c0c",
X"5d800b81",
X"1b347983",
X"e0980c80",
X"567583e0",
X"800c973d",
X"0d04e93d",
X"0d83e098",
X"08568554",
X"75802e81",
X"8238800b",
X"81173499",
X"3de01146",
X"6a548a3d",
X"705458ec",
X"0551f6e6",
X"3f83e080",
X"085483e0",
X"800880df",
X"38893d33",
X"5473802e",
X"913802ab",
X"05337084",
X"2a810651",
X"5574802e",
X"86388354",
X"80c13976",
X"51f48a3f",
X"83e08008",
X"a0170c02",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"9c1c0c52",
X"78981b0c",
X"53565957",
X"810b8117",
X"34745473",
X"83e0800c",
X"993d0d04",
X"f53d0d7d",
X"7f617283",
X"e098085a",
X"5d5d595c",
X"807b0c85",
X"5775802e",
X"81e03881",
X"16338106",
X"55845774",
X"802e81d2",
X"38913974",
X"81173486",
X"39800b81",
X"17348157",
X"81c0399c",
X"16089817",
X"08315574",
X"78278338",
X"74587780",
X"2e81a938",
X"98160870",
X"83ff0656",
X"577480cf",
X"38821633",
X"ff057789",
X"2a067081",
X"ff065a55",
X"78a03876",
X"8738a016",
X"08558d39",
X"a4160851",
X"f0ea3f83",
X"e0800855",
X"817527ff",
X"a83874a4",
X"170ca416",
X"0851f284",
X"3f83e080",
X"085583e0",
X"8008802e",
X"ff893883",
X"e0800819",
X"a8170c98",
X"160883ff",
X"06848071",
X"31515577",
X"75278338",
X"77557483",
X"ffff0654",
X"98160883",
X"ff0653a8",
X"16085279",
X"577b8338",
X"7b577651",
X"8a8d3f83",
X"e08008fe",
X"d0389816",
X"08159817",
X"0c741a78",
X"76317c08",
X"177d0c59",
X"5afed339",
X"80577683",
X"e0800c8d",
X"3d0d04fa",
X"3d0d7883",
X"e0980855",
X"56855573",
X"802e81e1",
X"38811433",
X"81065384",
X"5572802e",
X"81d3389c",
X"14085372",
X"76278338",
X"72569814",
X"0857800b",
X"98150c75",
X"802e81b7",
X"38821433",
X"70892b56",
X"5376802e",
X"b5387452",
X"ff1651ba",
X"d03f83e0",
X"8008ff18",
X"76547053",
X"5853bac1",
X"3f83e080",
X"08732696",
X"38743070",
X"78067098",
X"170c7771",
X"31a41708",
X"52585153",
X"8939a014",
X"0870a416",
X"0c537476",
X"27b93872",
X"51eed93f",
X"83e08008",
X"53810b83",
X"e0800827",
X"8b388814",
X"0883e080",
X"08268838",
X"800b8115",
X"34b03983",
X"e08008a4",
X"150c9814",
X"08159815",
X"0c757531",
X"56c43998",
X"14081670",
X"98160c73",
X"5256efc8",
X"3f83e080",
X"088c3883",
X"e0800881",
X"15348155",
X"94398214",
X"33ff0576",
X"892a0683",
X"e0800805",
X"a8150c80",
X"557483e0",
X"800c883d",
X"0d04ef3d",
X"0d635685",
X"5583e098",
X"08802e80",
X"d238933d",
X"f4058417",
X"0c645388",
X"3d705376",
X"5257f1d2",
X"3f83e080",
X"085583e0",
X"8008b438",
X"883d3354",
X"73802ea1",
X"3802a705",
X"3370842a",
X"70810651",
X"55558355",
X"73802e97",
X"387651ee",
X"f83f83e0",
X"80088817",
X"0c7551ef",
X"a93f83e0",
X"80085574",
X"83e0800c",
X"933d0d04",
X"e43d0d6e",
X"a13d0840",
X"5e855683",
X"e0980880",
X"2e848538",
X"9e3df405",
X"841f0c7e",
X"98387d51",
X"eef83f83",
X"e0800856",
X"83ee3981",
X"4181f639",
X"834181f1",
X"39933d7f",
X"96054159",
X"807f8295",
X"055e5675",
X"6081ff05",
X"34834190",
X"1e08762e",
X"81d338a0",
X"547d2270",
X"852b83e0",
X"06545890",
X"1e085278",
X"5186983f",
X"83e08008",
X"4183e080",
X"08ffb838",
X"78335c7b",
X"802effb4",
X"388b1933",
X"70bf0671",
X"81065243",
X"5574802e",
X"80de387b",
X"81bf0655",
X"748f2480",
X"d3389a19",
X"33557480",
X"cb38f31d",
X"70585d81",
X"56758b2e",
X"09810685",
X"388e568b",
X"39759a2e",
X"09810683",
X"389c5675",
X"19707081",
X"05523371",
X"33811a82",
X"1a5f5b52",
X"5b557486",
X"38797734",
X"853980df",
X"7734777b",
X"57577aa0",
X"2e098106",
X"c0388156",
X"7b81e532",
X"7030709f",
X"2a515155",
X"7bae2e93",
X"3874802e",
X"8e386183",
X"2a708106",
X"51557480",
X"2e97387d",
X"51ede23f",
X"83e08008",
X"4183e080",
X"08873890",
X"1e08feaf",
X"38806034",
X"75802e88",
X"387c527f",
X"5183a53f",
X"60802e86",
X"38800b90",
X"1f0c6056",
X"60832e85",
X"386081d0",
X"38891f57",
X"901e0880",
X"2e81a838",
X"80567519",
X"70335155",
X"74a02ea0",
X"3874852e",
X"09810684",
X"3881e555",
X"74777081",
X"05593481",
X"167081ff",
X"06575587",
X"7627d738",
X"88193355",
X"74a02ea9",
X"38ae7770",
X"81055934",
X"88567519",
X"70335155",
X"74a02e95",
X"38747770",
X"81055934",
X"81167081",
X"ff065755",
X"8a7627e2",
X"388b1933",
X"7f880534",
X"9f19339e",
X"1a337198",
X"2b71902b",
X"079d1c33",
X"70882b72",
X"079c1e33",
X"7107640c",
X"52991d33",
X"981e3371",
X"882b0753",
X"51535759",
X"56747f84",
X"05239719",
X"33961a33",
X"71882b07",
X"5656747f",
X"86052380",
X"77347d51",
X"ebf33f83",
X"e0800883",
X"32703070",
X"72079f2c",
X"83e08008",
X"06525656",
X"961f3355",
X"748a3889",
X"1f52961f",
X"5181b13f",
X"7583e080",
X"0c9e3d0d",
X"04fd3d0d",
X"75775354",
X"73335170",
X"89387133",
X"5170802e",
X"a1387333",
X"72335253",
X"72712785",
X"38ff5194",
X"39707327",
X"85388151",
X"8b398114",
X"81135354",
X"d3398051",
X"7083e080",
X"0c853d0d",
X"04fd3d0d",
X"75775454",
X"72337081",
X"ff065252",
X"70802ea3",
X"387181ff",
X"068114ff",
X"bf125354",
X"52709926",
X"8938a012",
X"7081ff06",
X"53517174",
X"70810556",
X"34d23980",
X"7434853d",
X"0d04ffbd",
X"3d0d80c6",
X"3d0852a5",
X"3d705254",
X"ffb33f80",
X"c73d0852",
X"853d7052",
X"53ffa63f",
X"72527351",
X"fedf3f80",
X"c53d0d04",
X"fe3d0d74",
X"76535371",
X"70810553",
X"33517073",
X"70810555",
X"3470f038",
X"843d0d04",
X"fe3d0d74",
X"52807233",
X"52537073",
X"2e8d3881",
X"12811471",
X"33535452",
X"70f53872",
X"83e0800c",
X"843d0d04",
X"fc3d0d76",
X"557483e3",
X"98082eaf",
X"38805374",
X"5187cb3f",
X"83e08008",
X"81ff06ff",
X"147081ff",
X"06723070",
X"9f2a5152",
X"55535472",
X"802e8438",
X"71dd3873",
X"fe387483",
X"e3980c86",
X"3d0d04ff",
X"3d0dff0b",
X"83e3980c",
X"84af3f81",
X"51878f3f",
X"83e08008",
X"81ff0652",
X"71ee3881",
X"d63f7183",
X"e0800c83",
X"3d0d04fc",
X"3d0d7602",
X"8405a205",
X"22028805",
X"a605227a",
X"54555555",
X"ff823f72",
X"802ea038",
X"83e3ac14",
X"33757081",
X"05573481",
X"147083ff",
X"ff06ff15",
X"7083ffff",
X"06565255",
X"52dd3980",
X"0b83e080",
X"0c863d0d",
X"04fc3d0d",
X"76787a11",
X"56535580",
X"5371742e",
X"93387215",
X"51703383",
X"e3ac1334",
X"81128114",
X"5452ea39",
X"800b83e0",
X"800c863d",
X"0d04fd3d",
X"0d905483",
X"e3980851",
X"86fe3f83",
X"e0800881",
X"ff06ff15",
X"71307130",
X"7073079f",
X"2a729f2a",
X"06525552",
X"555372db",
X"38853d0d",
X"04ff3d0d",
X"83e3a408",
X"1083e39c",
X"080780ff",
X"a8085271",
X"0c833d0d",
X"04800b83",
X"e3a40ce1",
X"3f04810b",
X"83e3a40c",
X"d83f04ed",
X"3f047183",
X"e3a00c04",
X"803d0d80",
X"51f43f81",
X"0b83e3a4",
X"0c810b83",
X"e39c0cff",
X"b83f823d",
X"0d04803d",
X"0d723070",
X"74078025",
X"83e39c0c",
X"51ffa23f",
X"823d0d04",
X"fe3d0d02",
X"93053380",
X"ffac0854",
X"730c80ff",
X"a8085271",
X"08708106",
X"515170f7",
X"38720870",
X"81ff0683",
X"e0800c51",
X"843d0d04",
X"803d0d81",
X"ff51cd3f",
X"83e08008",
X"81ff0683",
X"e0800c82",
X"3d0d04ff",
X"3d0d7490",
X"2b740780",
X"ff9c0852",
X"710c833d",
X"0d0404fb",
X"3d0d7802",
X"84059f05",
X"3370982b",
X"55575572",
X"80259b38",
X"7580ff06",
X"56805280",
X"f751e03f",
X"83e08008",
X"81ff0654",
X"73812680",
X"ff388051",
X"fee03fff",
X"9f3f8151",
X"fed83fff",
X"973f7551",
X"fee63f74",
X"982a51fe",
X"df3f7490",
X"2a7081ff",
X"065253fe",
X"d33f7488",
X"2a7081ff",
X"065253fe",
X"c73f7481",
X"ff0651fe",
X"bf3f8155",
X"7580c02e",
X"09810686",
X"38819555",
X"8d397580",
X"c82e0981",
X"06843881",
X"87557451",
X"fe9e3f8a",
X"55fec53f",
X"83e08008",
X"81ff0670",
X"982b5454",
X"7280258c",
X"38ff1570",
X"81ff0656",
X"5374e238",
X"7383e080",
X"0c873d0d",
X"04fa3d0d",
X"fdbe3f80",
X"51fdd33f",
X"8a54fe90",
X"3fff1470",
X"81ff0655",
X"5373f338",
X"73745355",
X"80c051fe",
X"a63f83e0",
X"800881ff",
X"06547381",
X"2e098106",
X"829f3883",
X"aa5280c8",
X"51fe8c3f",
X"83e08008",
X"81ff0653",
X"72812e09",
X"810681a8",
X"38745487",
X"3d741154",
X"56fdc53f",
X"83e08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e53802",
X"9a053353",
X"72812e09",
X"810681d9",
X"38029b05",
X"335380ce",
X"90547281",
X"aa2e8d38",
X"81c73980",
X"e4518ace",
X"3fff1454",
X"73802e81",
X"b838820a",
X"5281e951",
X"fda53f83",
X"e0800881",
X"ff065372",
X"de387252",
X"80fa51fd",
X"923f83e0",
X"800881ff",
X"06537281",
X"90387254",
X"731653fc",
X"d33f83e0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e8",
X"38873d33",
X"70862a70",
X"81065154",
X"548c5572",
X"80e33884",
X"5580de39",
X"745281e9",
X"51fccc3f",
X"83e08008",
X"81ff0653",
X"825581e9",
X"56817327",
X"86387355",
X"80c15680",
X"ce90548a",
X"3980e451",
X"89c03fff",
X"14547380",
X"2ea93880",
X"527551fc",
X"9a3f83e0",
X"800881ff",
X"065372e1",
X"38848052",
X"80d051fc",
X"863f83e0",
X"800881ff",
X"06537280",
X"2e833880",
X"557483e3",
X"a8348051",
X"fb803ffb",
X"bf3f883d",
X"0d04fb3d",
X"0d775480",
X"0b83e3a8",
X"3370832a",
X"70810651",
X"55575572",
X"752e0981",
X"06853873",
X"892b5473",
X"5280d151",
X"fbbd3f83",
X"e0800881",
X"ff065372",
X"bd3882b8",
X"c054fb80",
X"3f83e080",
X"0881ff06",
X"537281ff",
X"2e098106",
X"8938ff14",
X"5473e738",
X"9f397281",
X"fe2e0981",
X"06963883",
X"e7ac5283",
X"e3ac51fa",
X"ea3ffad0",
X"3ffacd3f",
X"83398155",
X"8051fa82",
X"3ffac13f",
X"7481ff06",
X"83e0800c",
X"873d0d04",
X"fb3d0d77",
X"83e3ac56",
X"548151f9",
X"e53f83e3",
X"a8337083",
X"2a708106",
X"51545672",
X"85387389",
X"2b547352",
X"80d851fa",
X"b63f83e0",
X"800881ff",
X"06537280",
X"e43881ff",
X"51f9cd3f",
X"81fe51f9",
X"c73f8480",
X"53747081",
X"05563351",
X"f9ba3fff",
X"137083ff",
X"ff065153",
X"72eb3872",
X"51f9a93f",
X"7251f9a4",
X"3ff9cd3f",
X"83e08008",
X"9f0653a7",
X"88547285",
X"2e8c3899",
X"3980e451",
X"86f83fff",
X"1454f9b0",
X"3f83e080",
X"0881ff2e",
X"843873e9",
X"388051f8",
X"dd3ff99c",
X"3f800b83",
X"e0800c87",
X"3d0d0471",
X"83e7b00c",
X"8880800b",
X"83e7ac0c",
X"8480800b",
X"83e7b40c",
X"04fd3d0d",
X"77701755",
X"7705ff1a",
X"535371ff",
X"2e943873",
X"70810555",
X"33517073",
X"70810555",
X"34ff1252",
X"e939853d",
X"0d04fc3d",
X"0d80feb8",
X"08557433",
X"83e7b834",
X"a05483a0",
X"805383e7",
X"b0085283",
X"e7ac0851",
X"ffb73fa0",
X"5483a480",
X"5383e7b0",
X"085283e7",
X"ac0851ff",
X"a43f9054",
X"83a88053",
X"83e7b008",
X"5283e7ac",
X"0851ff91",
X"3fa05380",
X"5283e7b4",
X"0883a080",
X"055185d2",
X"3fa05380",
X"5283e7b4",
X"0883a480",
X"055185c2",
X"3f905380",
X"5283e7b4",
X"0883a880",
X"055185b2",
X"3f80feb8",
X"0855ff75",
X"3483a080",
X"54805383",
X"e7b00852",
X"83e7b408",
X"51fec63f",
X"80d08054",
X"83b08053",
X"83e7b008",
X"5283e7b4",
X"0851feb1",
X"3f86d33f",
X"a2548053",
X"83e7b408",
X"8c800552",
X"80fcac51",
X"fe9b3f80",
X"fedc0855",
X"86753480",
X"fee00855",
X"80753480",
X"fed80855",
X"80753480",
X"fec80855",
X"af753480",
X"fed40855",
X"bf753480",
X"fed00855",
X"80753480",
X"fecc0855",
X"9f753480",
X"fec40855",
X"80753480",
X"feb00855",
X"e0753480",
X"fea80855",
X"a2753480",
X"fea40855",
X"83753480",
X"feac0855",
X"82753486",
X"3d0d04fc",
X"3d0d83a0",
X"80548053",
X"83e7b408",
X"5283e7b0",
X"0851fda1",
X"3f80d080",
X"5483b080",
X"5383e7b4",
X"085283e7",
X"b00851fd",
X"8c3fa054",
X"83a08053",
X"83e7b408",
X"5283e7b0",
X"0851fcf9",
X"3fa05483",
X"a4805383",
X"e7b40852",
X"83e7b008",
X"51fce63f",
X"905483a8",
X"805383e7",
X"b4085283",
X"e7b00851",
X"fcd33f80",
X"feb80855",
X"83e7b833",
X"7534863d",
X"0d04803d",
X"0d80ffc0",
X"08700881",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d80ffc0",
X"08700870",
X"fe067607",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"ffc00870",
X"0870812c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"ff3d0d80",
X"ffc00870",
X"0870fd06",
X"76100772",
X"0c525283",
X"3d0d0480",
X"3d0d80ff",
X"c0087008",
X"70822cbf",
X"0683e080",
X"0c515182",
X"3d0d04ff",
X"3d0d80ff",
X"c0087008",
X"70fe8306",
X"76822b07",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"ffc00870",
X"0870882c",
X"870683e0",
X"800c5151",
X"823d0d04",
X"ff3d0d80",
X"ffc00870",
X"0870f1ff",
X"0676882b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80ffc008",
X"7008708b",
X"2cbf0683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80ffc008",
X"700870f8",
X"8fff0676",
X"8b2b0772",
X"0c525283",
X"3d0d0480",
X"3d0d80ff",
X"c0087008",
X"70912cbf",
X"0683e080",
X"0c515182",
X"3d0d04ff",
X"3d0d80ff",
X"c0087008",
X"70fc87ff",
X"ff067691",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d80ffd0",
X"08700870",
X"882c8106",
X"83e0800c",
X"5151823d",
X"0d04803d",
X"0d80ffd0",
X"08700870",
X"892c8106",
X"83e0800c",
X"5151823d",
X"0d04803d",
X"0d80ffd0",
X"08700870",
X"8a2c8106",
X"83e0800c",
X"5151823d",
X"0d04803d",
X"0d80ffd0",
X"08700870",
X"8b2c8106",
X"83e0800c",
X"5151823d",
X"0d04fd3d",
X"0d7581e6",
X"29872a80",
X"ffb00854",
X"730c853d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"81055434",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727084",
X"05540cff",
X"1151f039",
X"843d0d04",
X"fe3d0d84",
X"80805380",
X"5288800a",
X"51ffb33f",
X"81808053",
X"80528280",
X"0a51c63f",
X"843d0d04",
X"803d0d81",
X"51fc9b3f",
X"72802e83",
X"38d23f81",
X"51fcbd3f",
X"8051fcb8",
X"3f8051fc",
X"853f823d",
X"0d04fd3d",
X"0d755280",
X"5480ff72",
X"25883881",
X"0bff8013",
X"5354ffbf",
X"12517099",
X"268638e0",
X"12529e39",
X"ff9f1251",
X"99712795",
X"38d012e0",
X"13705454",
X"51897127",
X"88388f73",
X"27833880",
X"5273802e",
X"85388180",
X"12527181",
X"ff0683e0",
X"800c853d",
X"0d04803d",
X"0d84d8c0",
X"51807170",
X"81055334",
X"7084e0c0",
X"2e098106",
X"f038823d",
X"0d04fe3d",
X"0d029705",
X"3351ff86",
X"3f83e080",
X"0881ff06",
X"83e7bc08",
X"54528073",
X"249b3883",
X"e7d80813",
X"7283e7dc",
X"08075353",
X"71733483",
X"e7bc0881",
X"0583e7bc",
X"0c843d0d",
X"04fa3d0d",
X"82800a1b",
X"55805788",
X"3dfc0554",
X"79537452",
X"7851cbd2",
X"3f883d0d",
X"04fe3d0d",
X"83e7d408",
X"527451d2",
X"b63f83e0",
X"80088c38",
X"76537552",
X"83e7d408",
X"51c73f84",
X"3d0d04fe",
X"3d0d83e7",
X"d4085375",
X"527451cc",
X"f53f83e0",
X"80088d38",
X"77537652",
X"83e7d408",
X"51ffa23f",
X"843d0d04",
X"fe3d0d83",
X"e7d40851",
X"cbe93f83",
X"e0800881",
X"80802e09",
X"81068838",
X"83c18080",
X"539b3983",
X"e7d40851",
X"cbcd3f83",
X"e0800880",
X"d0802e09",
X"81069338",
X"83c1b080",
X"5383e080",
X"085283e7",
X"d40851fe",
X"d83f843d",
X"0d04803d",
X"0dfa993f",
X"83e08008",
X"842980fc",
X"d0057008",
X"83e0800c",
X"51823d0d",
X"04ee3d0d",
X"80438042",
X"80418070",
X"5a5bfdd2",
X"3f800b83",
X"e7bc0c80",
X"0b83e7dc",
X"0c80faac",
X"51c6b93f",
X"81800b83",
X"e7dc0c80",
X"fab051c6",
X"ab3f80d0",
X"0b83e7bc",
X"0c783070",
X"7a078025",
X"70872b83",
X"e7dc0c51",
X"55f9883f",
X"83e08008",
X"5280fab8",
X"51c6853f",
X"80f80b83",
X"e7bc0c78",
X"81327030",
X"70720780",
X"2570872b",
X"83e7dc0c",
X"515656fe",
X"f13f83e0",
X"80085280",
X"fac451c5",
X"db3f81a0",
X"0b83e7bc",
X"0c788232",
X"70307072",
X"07802570",
X"872b83e7",
X"dc0c5156",
X"83e7d408",
X"5256c6f5",
X"3f83e080",
X"085280fa",
X"cc51c5ac",
X"3f81f00b",
X"83e7bc0c",
X"810b83e7",
X"c05b5883",
X"e7bc0882",
X"197a3270",
X"30707207",
X"80257087",
X"2b83e7dc",
X"0c51578e",
X"3d7055ff",
X"1b545757",
X"5799923f",
X"79708405",
X"5b0851c6",
X"ac3f7454",
X"83e08008",
X"53775280",
X"fad451c4",
X"df3fa817",
X"83e7bc0c",
X"81185877",
X"852e0981",
X"06ffb038",
X"83900b83",
X"e7bc0c78",
X"87327030",
X"70720780",
X"2570872b",
X"83e7dc0c",
X"515656f8",
X"ba3f80fa",
X"e45583e0",
X"8008802e",
X"8e3883e7",
X"d00851c5",
X"d83f83e0",
X"80085574",
X"5280faec",
X"51c48d3f",
X"83e00b83",
X"e7bc0c78",
X"88327030",
X"70720780",
X"2570872b",
X"83e7dc0c",
X"515780fa",
X"f85255c3",
X"eb3f868d",
X"a051f982",
X"3f805291",
X"3d705255",
X"99ea3f83",
X"52745199",
X"e33f6119",
X"59788025",
X"85388059",
X"90398879",
X"25853888",
X"59873978",
X"882682db",
X"3878822b",
X"5580f988",
X"150804f6",
X"a23f83e0",
X"80086157",
X"5575812e",
X"09810689",
X"3883e080",
X"08105590",
X"3975ff2e",
X"09810688",
X"3883e080",
X"08812c55",
X"90752585",
X"38905588",
X"39748024",
X"83388155",
X"7451f5ff",
X"3f829039",
X"f6923f83",
X"e0800861",
X"05557480",
X"25853880",
X"55883987",
X"75258338",
X"87557451",
X"f68e3f81",
X"ee396087",
X"3862802e",
X"81e53883",
X"e0a40883",
X"e0a00c8c",
X"830b83e0",
X"a80c83e7",
X"d40851ff",
X"b4d33ffa",
X"e73f81c7",
X"39605680",
X"76259938",
X"8b9c0b83",
X"e0a80c83",
X"e7b41570",
X"085255ff",
X"b4b33f74",
X"08529139",
X"75802591",
X"3883e7b4",
X"150851c3",
X"c63f8052",
X"fd1951b8",
X"3962802e",
X"818d3883",
X"e7b41570",
X"0883e7c0",
X"08720c83",
X"e7c00cfd",
X"1a705351",
X"558b823f",
X"83e08008",
X"5680518a",
X"f83f83e0",
X"80085274",
X"5187903f",
X"75528051",
X"87893f80",
X"d6396055",
X"807525b8",
X"3883e0ac",
X"0883e0a0",
X"0c8c830b",
X"83e0a80c",
X"83e7d008",
X"51ffb3bd",
X"3f83e7d0",
X"0851ffb0",
X"b33f83e0",
X"800881ff",
X"06705255",
X"f5a13f74",
X"802e9c38",
X"8155a039",
X"74802593",
X"3883e7d0",
X"0851c2b7",
X"3f8051f5",
X"863f8439",
X"6287387a",
X"802efa8a",
X"38805574",
X"83e0800c",
X"943d0d04",
X"fe3d0df5",
X"853f83e0",
X"8008802e",
X"86388051",
X"80f739f5",
X"8d3f83e0",
X"800880eb",
X"38f5b33f",
X"83e08008",
X"802eaa38",
X"8151f2d2",
X"3fefa73f",
X"800b83e7",
X"bc0cf9b9",
X"3f83e080",
X"0853ff0b",
X"83e7bc0c",
X"f1b13f72",
X"be387251",
X"f2b03fbc",
X"39f4e73f",
X"83e08008",
X"802eb138",
X"8151f29e",
X"3feef33f",
X"8b9c0b83",
X"e0a80c83",
X"e7c00851",
X"ffb2823f",
X"ff0b83e7",
X"bc0cf0fb",
X"3f83e7c0",
X"08528051",
X"85993f81",
X"51f5d13f",
X"843d0d04",
X"fc3d0d90",
X"80805286",
X"84808051",
X"c58a3f83",
X"e0800880",
X"c33888ea",
X"3f80ffd4",
X"51c9ca3f",
X"83e08008",
X"559c800a",
X"5480c080",
X"5380fb80",
X"5283e080",
X"0851f79f",
X"3f83e7d4",
X"085380fb",
X"90527451",
X"c4943f83",
X"e0800884",
X"38f7ad3f",
X"8151f4f8",
X"3f92f63f",
X"8151f4f0",
X"3ffe913f",
X"fc3983e0",
X"8c080283",
X"e08c0cfb",
X"3d0d0280",
X"fb9c0b83",
X"e0a40c80",
X"fba00b83",
X"e09c0c80",
X"fba40b83",
X"e0ac0c83",
X"e08c08fc",
X"050c800b",
X"83e7c00b",
X"83e08c08",
X"f8050c83",
X"e08c08f4",
X"050cc2ec",
X"3f83e080",
X"088605fc",
X"0683e08c",
X"08f0050c",
X"0283e08c",
X"08f00508",
X"310d833d",
X"7083e08c",
X"08f80508",
X"70840583",
X"e08c08f8",
X"050c0c51",
X"ffbfb43f",
X"83e08c08",
X"f4050881",
X"0583e08c",
X"08f4050c",
X"83e08c08",
X"f4050886",
X"2e098106",
X"ffac3886",
X"94808051",
X"ec893fff",
X"0b83e7bc",
X"0c800b83",
X"e7dc0c84",
X"d8c00b83",
X"e7d80c81",
X"51efd73f",
X"8151f080",
X"3f8051ef",
X"fb3f8151",
X"f0a53f81",
X"51f1823f",
X"8251f0cc",
X"3f8051f1",
X"aa3f80d1",
X"ae528051",
X"ffbcf23f",
X"fdbe3f83",
X"e08c08fc",
X"05080d80",
X"0b83e080",
X"0c873d0d",
X"83e08c0c",
X"04803d0d",
X"81ff5180",
X"0b83e7e8",
X"1234ff11",
X"5170f438",
X"823d0d04",
X"ff3d0d73",
X"70335351",
X"81113371",
X"34718112",
X"34833d0d",
X"04fb3d0d",
X"77795656",
X"80707155",
X"55527175",
X"25ac3872",
X"16703370",
X"147081ff",
X"06555151",
X"51717427",
X"89388112",
X"7081ff06",
X"53517181",
X"147083ff",
X"ff065552",
X"54747324",
X"d6387183",
X"e0800c87",
X"3d0d04fc",
X"3d0d7655",
X"ffb69b3f",
X"83e08008",
X"802ef538",
X"83ea8408",
X"86057081",
X"ff065253",
X"ffb3f23f",
X"8439fb80",
X"3fffb5fa",
X"3f83e080",
X"08812ef2",
X"38805473",
X"1553ffb4",
X"ce3f83e0",
X"80087334",
X"81145473",
X"852e0981",
X"06e93884",
X"39fad53f",
X"ffb5cf3f",
X"83e08008",
X"802ef238",
X"743383e7",
X"e8348115",
X"3383e7e9",
X"34821533",
X"83e7ea34",
X"83153383",
X"e7eb3484",
X"5283e7e8",
X"51feba3f",
X"83e08008",
X"81ff0684",
X"16335653",
X"72752e09",
X"81068d38",
X"ffb4bf3f",
X"83e08008",
X"802e9a38",
X"83ea8408",
X"a82e0981",
X"06893886",
X"0b83ea84",
X"0c8739a8",
X"0b83ea84",
X"0c80e451",
X"efd03f86",
X"3d0d04f4",
X"3d0d7e60",
X"5955805d",
X"8075822b",
X"7183ea88",
X"120c83ea",
X"9c175b5b",
X"57767934",
X"77772e83",
X"b8387652",
X"7751ffbd",
X"fd3f8e3d",
X"fc055490",
X"5383e9f0",
X"527751ff",
X"bdb83f7c",
X"5675902e",
X"09810683",
X"943883e9",
X"f051fd94",
X"3f83e9f2",
X"51fd8d3f",
X"83e9f451",
X"fd863f76",
X"83ea800c",
X"7751ffbb",
X"843f80f9",
X"bc5283e0",
X"800851ff",
X"aa883f83",
X"e0800881",
X"2e098106",
X"80d43876",
X"83ea980c",
X"820b83e9",
X"f034ff96",
X"0b83e9f1",
X"347751ff",
X"bdc93f83",
X"e0800855",
X"83e08008",
X"77258838",
X"83e08008",
X"8f055574",
X"842c7083",
X"ffff0670",
X"882a5851",
X"557583e9",
X"f2347483",
X"e9f33476",
X"83e9f434",
X"ff800b83",
X"e9f53481",
X"903983e9",
X"f03383e9",
X"f1337188",
X"2b07565b",
X"7483ffff",
X"2e098106",
X"80e838fe",
X"800b83ea",
X"980c810b",
X"83ea800c",
X"ff0b83e9",
X"f034ff0b",
X"83e9f134",
X"7751ffbc",
X"d63f83e0",
X"800883ea",
X"a00c83e0",
X"80085583",
X"e0800880",
X"25883883",
X"e080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583e9f2",
X"347483e9",
X"f3347683",
X"e9f434ff",
X"800b83e9",
X"f534810b",
X"83e9ff34",
X"a5397485",
X"962e0981",
X"0680fe38",
X"7583ea98",
X"0c7751ff",
X"bc8a3f83",
X"e9ff3383",
X"e0800807",
X"557483e9",
X"ff3483e9",
X"ff338106",
X"5574802e",
X"83388457",
X"83e9f433",
X"83e9f533",
X"71882b07",
X"565c7481",
X"802e0981",
X"06a13883",
X"e9f23383",
X"e9f33371",
X"882b0756",
X"5bad8075",
X"27873876",
X"8207579c",
X"39768107",
X"57963974",
X"82802e09",
X"81068738",
X"76830757",
X"87397481",
X"ff268a38",
X"7783ea88",
X"1b0c7679",
X"348e3d0d",
X"04803d0d",
X"72842983",
X"ea880570",
X"0883e080",
X"0c51823d",
X"0d04fe3d",
X"0d800b83",
X"e9ec0c80",
X"0b83e9e8",
X"0cff0b83",
X"e7e40ca8",
X"0b83ea84",
X"0cae51ff",
X"aebb3f80",
X"0b83ea88",
X"54528073",
X"70840555",
X"0c811252",
X"71842e09",
X"8106ef38",
X"843d0d04",
X"fe3d0d74",
X"02840596",
X"05225353",
X"71802e97",
X"38727081",
X"05543351",
X"ffaed93f",
X"ff127083",
X"ffff0651",
X"52e63984",
X"3d0d04fe",
X"3d0d0292",
X"05225382",
X"ac51eae2",
X"3f80c351",
X"ffaeb53f",
X"819651ea",
X"d53f7252",
X"83e7e851",
X"ffb23f72",
X"5283e7e8",
X"51f8ee3f",
X"83e08008",
X"81ff0651",
X"ffae913f",
X"843d0d04",
X"ffb13d0d",
X"80d13df8",
X"0551f997",
X"3f83e9ec",
X"08810583",
X"e9ec0c80",
X"cf3d33cf",
X"117081ff",
X"06515656",
X"74832688",
X"ed38758f",
X"06ff0556",
X"7583e7e4",
X"082e9b38",
X"75832696",
X"387583e7",
X"e40c7584",
X"2983ea88",
X"05700853",
X"557551fa",
X"963f8076",
X"2488c938",
X"75842983",
X"ea880555",
X"7408802e",
X"88ba3883",
X"e7e40884",
X"2983ea88",
X"05700802",
X"880582b9",
X"0533525b",
X"557480d2",
X"2e84b138",
X"7480d224",
X"903874bf",
X"2e9c3874",
X"80d02e81",
X"d73887f8",
X"397480d3",
X"2e80d238",
X"7480d72e",
X"81c63887",
X"e7390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290556",
X"56ffad93",
X"3f80c151",
X"ffacc53f",
X"f6e73f86",
X"0b83e7e8",
X"34815283",
X"e7e851ff",
X"ae803f81",
X"51fde43f",
X"74893886",
X"0b83ea84",
X"0c8739a8",
X"0b83ea84",
X"0cffacdf",
X"3f80c151",
X"ffac913f",
X"f6b33f90",
X"0b83e9ff",
X"33810656",
X"5674802e",
X"83389856",
X"83e9f433",
X"83e9f533",
X"71882b07",
X"56597481",
X"802e0981",
X"069c3883",
X"e9f23383",
X"e9f33371",
X"882b0756",
X"57ad8075",
X"278c3875",
X"81800756",
X"853975a0",
X"07567583",
X"e7e834ff",
X"0b83e7e9",
X"34e00b83",
X"e7ea3480",
X"0b83e7eb",
X"34845283",
X"e7e851ff",
X"acf43f84",
X"51869e39",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"055659ff",
X"abd13f79",
X"51ffb6d0",
X"3f83e080",
X"08802e8b",
X"3880ce51",
X"ffaaf53f",
X"85f23980",
X"c151ffaa",
X"eb3fffab",
X"f33fffa9",
X"f53f83ea",
X"98085883",
X"75259b38",
X"83e9f433",
X"83e9f533",
X"71882b07",
X"fc177129",
X"7a058380",
X"055a5157",
X"8d397481",
X"802918ff",
X"80055881",
X"80578056",
X"76762e93",
X"38ffaac7",
X"3f83e080",
X"0883e7e8",
X"17348116",
X"56ea39ff",
X"aab53f83",
X"e0800881",
X"ff067753",
X"83e7e852",
X"56f4d63f",
X"83e08008",
X"81ff0655",
X"75752e09",
X"8106818a",
X"38ffaab7",
X"3f80c151",
X"ffa9e93f",
X"ffaaf13f",
X"77527951",
X"ffb4df3f",
X"805e80d1",
X"3dfdf405",
X"54765383",
X"e7e85279",
X"51ffb2ec",
X"3f0282b9",
X"05335581",
X"587480d7",
X"2e098106",
X"bd3880d1",
X"3dfdf005",
X"5476538f",
X"3d70537a",
X"5259ffb3",
X"f13f8056",
X"76762ea2",
X"38751983",
X"e7e81733",
X"71337072",
X"32703070",
X"80257030",
X"7e06811d",
X"5d5e5151",
X"51525b55",
X"db3982ac",
X"51e59b3f",
X"77802e86",
X"3880c351",
X"843980ce",
X"51ffa8e4",
X"3fffa9ec",
X"3fffa7ee",
X"3f83dd39",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"05595580",
X"705d59ff",
X"a9853f80",
X"c151ffa8",
X"b73f83ea",
X"8008792e",
X"82de3883",
X"eaa00880",
X"fc055580",
X"fd527451",
X"868b3f83",
X"e080085b",
X"778224b2",
X"38ff1870",
X"872b83ff",
X"ff800680",
X"fcf00583",
X"e7e85957",
X"55818055",
X"75708105",
X"57337770",
X"81055934",
X"ff157081",
X"ff065155",
X"74ea3882",
X"8d397782",
X"e82e81ab",
X"387782e9",
X"2e098106",
X"81b23880",
X"fba851ff",
X"aed23f78",
X"58778732",
X"70307072",
X"0780257a",
X"8a327030",
X"70720780",
X"25730753",
X"545a5157",
X"5575802e",
X"97387878",
X"269238a0",
X"0b83e7e8",
X"1a348119",
X"7081ff06",
X"5a55eb39",
X"81187081",
X"ff065955",
X"8a7827ff",
X"bc388f58",
X"83e7e318",
X"3383e7e8",
X"1934ff18",
X"7081ff06",
X"59557784",
X"26ea3890",
X"58800b83",
X"e7e81934",
X"81187081",
X"ff067098",
X"2b525955",
X"748025e9",
X"3880c655",
X"7a858f24",
X"843880c2",
X"557483e7",
X"e83480f1",
X"0b83e7eb",
X"34810b83",
X"e7ec347a",
X"83e7e934",
X"7a882c55",
X"7483e7ea",
X"3480cb39",
X"82f07825",
X"80c43877",
X"80fd29fd",
X"97d30552",
X"7951ffb1",
X"8d3f80d1",
X"3dfdec05",
X"5480fd53",
X"83e7e852",
X"7951ffb0",
X"c53f7b81",
X"19595675",
X"80fc2483",
X"38785877",
X"882c5574",
X"83e8e534",
X"7783e8e6",
X"347583e8",
X"e7348180",
X"5980cc39",
X"83ea9808",
X"57837825",
X"9b3883e9",
X"f43383e9",
X"f5337188",
X"2b07fc1a",
X"71297905",
X"83800559",
X"51598d39",
X"77818029",
X"17ff8005",
X"57818059",
X"76527951",
X"ffb09b3f",
X"80d13dfd",
X"ec055478",
X"5383e7e8",
X"527951ff",
X"afd43f78",
X"51f6b83f",
X"ffa6893f",
X"ffa48b3f",
X"8b3983e9",
X"e8088105",
X"83e9e80c",
X"80d13d0d",
X"04f6d93f",
X"eb9e3ff9",
X"39fc3d0d",
X"76787184",
X"2983ea88",
X"05700851",
X"53535370",
X"9e3880ce",
X"723480cf",
X"0b811334",
X"80ce0b82",
X"133480c5",
X"0b831334",
X"70841334",
X"80e73983",
X"ea9c1333",
X"5480d272",
X"3473822a",
X"70810651",
X"5180cf53",
X"70843880",
X"d7537281",
X"1334a00b",
X"82133473",
X"83065170",
X"812e9e38",
X"70812488",
X"3870802e",
X"8f389f39",
X"70822e92",
X"3870832e",
X"92389339",
X"80d8558e",
X"3980d355",
X"893980cd",
X"55843980",
X"c4557483",
X"133480c4",
X"0b841334",
X"800b8513",
X"34863d0d",
X"04fd3d0d",
X"75548074",
X"0c800b84",
X"150c800b",
X"88150c80",
X"febc0870",
X"337081ff",
X"0670812a",
X"81327181",
X"32718106",
X"71810631",
X"841a0c56",
X"5670832a",
X"81327182",
X"2a813271",
X"81067181",
X"0631790c",
X"52555151",
X"5180feb4",
X"08703370",
X"09810688",
X"170c5151",
X"853d0d04",
X"fe3d0d74",
X"76545271",
X"51ff9a3f",
X"72812ea2",
X"38817326",
X"8d387282",
X"2eab3872",
X"832e9f38",
X"e6397108",
X"e2388412",
X"08dd3888",
X"1208d838",
X"a0398812",
X"08812e09",
X"8106cc38",
X"94398812",
X"08812e8d",
X"38710889",
X"38841208",
X"802effb7",
X"38843d0d",
X"0483e08c",
X"080283e0",
X"8c0cfd3d",
X"0d805383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"05085183",
X"d43f83e0",
X"80087083",
X"e0800c54",
X"853d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cfd3d0d",
X"815383e0",
X"8c088c05",
X"085283e0",
X"8c088805",
X"085183a1",
X"3f83e080",
X"087083e0",
X"800c5485",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"f93d0d80",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"88050880",
X"25b93883",
X"e08c0888",
X"05083083",
X"e08c0888",
X"050c800b",
X"83e08c08",
X"f4050c83",
X"e08c08fc",
X"05088a38",
X"810b83e0",
X"8c08f405",
X"0c83e08c",
X"08f40508",
X"83e08c08",
X"fc050c83",
X"e08c088c",
X"05088025",
X"b93883e0",
X"8c088c05",
X"083083e0",
X"8c088c05",
X"0c800b83",
X"e08c08f0",
X"050c83e0",
X"8c08fc05",
X"088a3881",
X"0b83e08c",
X"08f0050c",
X"83e08c08",
X"f0050883",
X"e08c08fc",
X"050c8053",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"81df3f83",
X"e0800870",
X"83e08c08",
X"f8050c54",
X"83e08c08",
X"fc050880",
X"2e903883",
X"e08c08f8",
X"05083083",
X"e08c08f8",
X"050c83e0",
X"8c08f805",
X"087083e0",
X"800c5489",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"fb3d0d80",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"88050880",
X"25993883",
X"e08c0888",
X"05083083",
X"e08c0888",
X"050c810b",
X"83e08c08",
X"fc050c83",
X"e08c088c",
X"05088025",
X"903883e0",
X"8c088c05",
X"083083e0",
X"8c088c05",
X"0c815383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"050851bd",
X"3f83e080",
X"087083e0",
X"8c08f805",
X"0c5483e0",
X"8c08fc05",
X"08802e90",
X"3883e08c",
X"08f80508",
X"3083e08c",
X"08f8050c",
X"83e08c08",
X"f8050870",
X"83e0800c",
X"54873d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cfd3d",
X"0d810b83",
X"e08c08fc",
X"050c800b",
X"83e08c08",
X"f8050c83",
X"e08c088c",
X"050883e0",
X"8c088805",
X"0827b938",
X"83e08c08",
X"fc050880",
X"2eae3880",
X"0b83e08c",
X"088c0508",
X"24a23883",
X"e08c088c",
X"05081083",
X"e08c088c",
X"050c83e0",
X"8c08fc05",
X"081083e0",
X"8c08fc05",
X"0cffb839",
X"83e08c08",
X"fc050880",
X"2e80e138",
X"83e08c08",
X"8c050883",
X"e08c0888",
X"050826ad",
X"3883e08c",
X"08880508",
X"83e08c08",
X"8c050831",
X"83e08c08",
X"88050c83",
X"e08c08f8",
X"050883e0",
X"8c08fc05",
X"080783e0",
X"8c08f805",
X"0c83e08c",
X"08fc0508",
X"812a83e0",
X"8c08fc05",
X"0c83e08c",
X"088c0508",
X"812a83e0",
X"8c088c05",
X"0cff9539",
X"83e08c08",
X"90050880",
X"2e933883",
X"e08c0888",
X"05087083",
X"e08c08f4",
X"050c5191",
X"3983e08c",
X"08f80508",
X"7083e08c",
X"08f4050c",
X"5183e08c",
X"08f40508",
X"83e0800c",
X"853d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cff3d0d",
X"800b83e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"8106ff11",
X"70097083",
X"e08c088c",
X"05080683",
X"e08c08fc",
X"05081183",
X"e08c08fc",
X"050c83e0",
X"8c088805",
X"08812a83",
X"e08c0888",
X"050c83e0",
X"8c088c05",
X"081083e0",
X"8c088c05",
X"0c515151",
X"5183e08c",
X"08880508",
X"802e8438",
X"ffab3983",
X"e08c08fc",
X"05087083",
X"e0800c51",
X"833d0d83",
X"e08c0c04",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002b5f",
X"00002ba0",
X"00002bc2",
X"00002be9",
X"00002be9",
X"00002be9",
X"00002be9",
X"00002c5a",
X"00002cac",
X"25732025",
X"73000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"6e616d65",
X"20000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00003ce8",
X"00003cec",
X"00003cf4",
X"00003d00",
X"00003d0c",
X"00003d18",
X"00003d24",
X"00003d28",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"0001d20f",
X"0001d400",
X"0001d401",
X"0001d409",
X"0001d010",
X"0001d301",
X"0001d300",
X"0001d20a",
X"0001d01b",
X"0001d016",
X"0001d019",
X"0001d018",
X"0001d017",
X"0001d01a",
X"0001d403",
X"0001d402",
X"0001d40e",
X"0004007c",
X"00040078",
X"00040074",
X"00040068",
X"00040060",
X"0004005c",
X"00040058",
X"00040054",
X"00040050",
X"0004004c",
X"00040048",
X"00040044",
X"00040040",
X"00040034",
X"00040030",
X"0004002c",
X"00040028",
X"00040024",
X"00040020",
X"0004001c",
X"00040018",
X"00040014",
X"00040010",
X"0004000c",
X"00040008",
X"00040004",
X"00040000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"69383030",
X"00000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
