
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80db",
X"9c738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80e0",
X"ac0c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580d6",
X"e72d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580d4fb",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"8d9f0480",
X"3d0d80e1",
X"c4087008",
X"810683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d80e1",
X"c4087008",
X"70fe0676",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80e1c408",
X"70087081",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80e1c408",
X"700870fd",
X"06761007",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"e1c40870",
X"0870822c",
X"bf0683e0",
X"800c5151",
X"823d0d04",
X"ff3d0d80",
X"e1c40870",
X"0870fe83",
X"0676822b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80e1c408",
X"70087088",
X"2c870683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80e1c408",
X"700870f1",
X"ff067688",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d80e1c4",
X"08700870",
X"8b2cbf06",
X"83e0800c",
X"5151823d",
X"0d04ff3d",
X"0d80e1c4",
X"08700870",
X"f88fff06",
X"768b2b07",
X"720c5252",
X"833d0d04",
X"fd3d0d75",
X"81e62987",
X"2a80e1b4",
X"0854730c",
X"853d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d848080",
X"53805288",
X"800a51ff",
X"b33f8180",
X"80538052",
X"82800a51",
X"c63f843d",
X"0d04803d",
X"0d8151fd",
X"dc3f7280",
X"2e8338d2",
X"3f8051fd",
X"d03f8051",
X"fd9d3f82",
X"3d0d04fd",
X"3d0d7552",
X"805480ff",
X"72258838",
X"810bff80",
X"135354ff",
X"bf125170",
X"99268638",
X"e012529e",
X"39ff9f12",
X"51997127",
X"9538d012",
X"e0137054",
X"54518971",
X"2788388f",
X"73278338",
X"80527380",
X"2e853881",
X"80125271",
X"81ff0683",
X"e0800c85",
X"3d0d0480",
X"3d0d823d",
X"0d04ff3d",
X"0d80e0d0",
X"0880e0e0",
X"08525271",
X"33713483",
X"3d0d0483",
X"e08c0802",
X"83e08c0c",
X"fd3d0d80",
X"0b83e09c",
X"0c86b8c0",
X"0b83e0a0",
X"0c8151fc",
X"b83f8151",
X"fce23f8d",
X"83528051",
X"9b803f80",
X"0b83e09c",
X"0c0b0b80",
X"dbac519a",
X"fc3f8480",
X"80528684",
X"8080519e",
X"a83f83e0",
X"8008818b",
X"380b0b80",
X"dbcc519a",
X"e03f9de2",
X"3f83e080",
X"088605fc",
X"0683e08c",
X"08f8050c",
X"0283e08c",
X"08f80508",
X"310d833d",
X"0b0b80db",
X"dc5283e0",
X"8c08fc05",
X"0c9ab23f",
X"83e08c08",
X"fc050852",
X"0b0b80db",
X"ec51a0de",
X"3f83e080",
X"0883e08c",
X"08f8050c",
X"83e08008",
X"aa380b0b",
X"80dbfc51",
X"9a873f88",
X"913f83e0",
X"8c08fc05",
X"085283e0",
X"8c08f805",
X"085184b1",
X"3f8151fd",
X"a93f918e",
X"3f92390b",
X"0b80dc8c",
X"5187390b",
X"0b80dca0",
X"5199d63f",
X"fe883ffc",
X"39803d0d",
X"81ff5180",
X"0b83e0a8",
X"1234ff11",
X"5170f438",
X"823d0d04",
X"ff3d0d73",
X"70335351",
X"81113371",
X"34718112",
X"34833d0d",
X"04fb3d0d",
X"77028405",
X"a2052255",
X"56807071",
X"55565271",
X"7427ac38",
X"72167033",
X"70147081",
X"ff065551",
X"51517175",
X"27893881",
X"127081ff",
X"06535171",
X"81147083",
X"ffff0655",
X"52557373",
X"26d63871",
X"83e0800c",
X"873d0d04",
X"fd3d0d75",
X"5493883f",
X"83e08008",
X"802ef638",
X"83e2c008",
X"86057081",
X"ff065253",
X"90e13f84",
X"39fceb3f",
X"92e93f83",
X"e0800881",
X"2ef33891",
X"c43f83e0",
X"80087434",
X"91bb3f83",
X"e0800881",
X"153491b1",
X"3f83e080",
X"08821534",
X"91a73f83",
X"e0800883",
X"1534919d",
X"3f83e080",
X"08841534",
X"8439fcaa",
X"3f92a83f",
X"83e08008",
X"802ef338",
X"80dcb451",
X"97e33f73",
X"3383e0a8",
X"34811433",
X"83e0a934",
X"82143383",
X"e0aa3483",
X"143383e0",
X"ab348452",
X"83e0a851",
X"fe9b3f83",
X"e0800881",
X"ff067433",
X"5380dcbc",
X"525397ad",
X"3f811433",
X"5280dcbc",
X"5197a23f",
X"82143352",
X"80dcbc51",
X"97973f83",
X"14335280",
X"dcbc5197",
X"8c3f8414",
X"335280dc",
X"bc519781",
X"3f725280",
X"dcbc5196",
X"f83f8414",
X"33547274",
X"2e098106",
X"8c3890d3",
X"3f83e080",
X"08802eb8",
X"3880dcc0",
X"5196da3f",
X"83e2c008",
X"a82e0981",
X"068d3886",
X"0b83e2c0",
X"0c80dcc8",
X"518b39a8",
X"0b83e2c0",
X"0c80dcd0",
X"5196b63f",
X"83e2c008",
X"5280dcbc",
X"5196aa3f",
X"80dc9c51",
X"96a33f80",
X"e451f8e8",
X"3f853d0d",
X"04fc3d0d",
X"76785555",
X"80537215",
X"70335351",
X"71802eba",
X"3871ae2e",
X"86388113",
X"53ec3973",
X"33811233",
X"54527173",
X"2e098106",
X"a1388114",
X"33821233",
X"54527173",
X"2e098106",
X"9138810b",
X"82153383",
X"13335355",
X"5273712e",
X"83388052",
X"7183e080",
X"0c863d0d",
X"04f63d0d",
X"7d57805b",
X"7c822b58",
X"800b83e2",
X"c4190c76",
X"802e83b2",
X"38805276",
X"5198813f",
X"8c3dfc05",
X"54905383",
X"e2b05276",
X"51979e3f",
X"7a567590",
X"2e883880",
X"dcd85182",
X"e33983e2",
X"b051fbc4",
X"3f83e2b2",
X"51fbbd3f",
X"83e2b451",
X"fbb63f80",
X"0b83e2bc",
X"0c765196",
X"c93f80dc",
X"f05283e0",
X"800851fe",
X"c03f83e0",
X"80089a38",
X"765196b2",
X"3f80dcf4",
X"5283e080",
X"0851fea9",
X"3f83e080",
X"08802ea3",
X"3880dcf8",
X"5194b23f",
X"800b83e2",
X"d40c820b",
X"83e2b034",
X"ff960b83",
X"e2b13476",
X"51978f3f",
X"80c73983",
X"e2b03383",
X"e2b13371",
X"882b0756",
X"597483ff",
X"ff2e0981",
X"0680e938",
X"80dd8051",
X"93f73ffe",
X"800b83e2",
X"d40c810b",
X"83e2bc0c",
X"ff0b83e2",
X"b034ff0b",
X"83e2b134",
X"765196ce",
X"3f83e080",
X"0883e2d8",
X"0c83e080",
X"085583e0",
X"80088025",
X"883883e0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83e2b234",
X"7483e2b3",
X"34800b83",
X"e2b434ff",
X"800b83e2",
X"b5349f39",
X"7485962e",
X"0981068f",
X"3880dd88",
X"5193863f",
X"7583e2d4",
X"0c883980",
X"dd905180",
X"d73983e2",
X"b43383e2",
X"b5337188",
X"2b075656",
X"7481802e",
X"098106a1",
X"3883e2b2",
X"3383e2b3",
X"3371882b",
X"07565aad",
X"80752787",
X"3880dda4",
X"51ab3980",
X"dda851a5",
X"39748280",
X"2e098106",
X"873880dd",
X"ac519639",
X"7481ff26",
X"873880dd",
X"b0518a39",
X"80ddb451",
X"929f3fa6",
X"39929a3f",
X"83e2b233",
X"83e2b333",
X"71882b07",
X"535980dc",
X"bc519285",
X"3f80ddc4",
X"5191fe3f",
X"7683e2c4",
X"190c8c3d",
X"0d04fe3d",
X"0d800b83",
X"e2ac0c80",
X"0b83e2a8",
X"0cff0b83",
X"e0a40ca8",
X"0b83e2c0",
X"0cae5189",
X"fa3f800b",
X"83e2c454",
X"52807370",
X"8405550c",
X"81125271",
X"842e0981",
X"06ef3884",
X"3d0d04fe",
X"3d0d7402",
X"84059605",
X"22535371",
X"802e9638",
X"72708105",
X"5433518a",
X"993fff12",
X"7083ffff",
X"065152e7",
X"39843d0d",
X"04fe3d0d",
X"02920522",
X"80ddc852",
X"5390fe3f",
X"725280dc",
X"bc5190f5",
X"3f82ac51",
X"f3ba3f80",
X"c35189e6",
X"3f819651",
X"f3ae3f72",
X"5283e0a8",
X"51ffa43f",
X"725283e0",
X"a851f7ad",
X"3f83e080",
X"0881ff06",
X"70525389",
X"c13f80dd",
X"d05190bd",
X"3f725280",
X"dcbc5190",
X"b43f80dd",
X"d85190ad",
X"3f843d0d",
X"04f33d0d",
X"8f3df805",
X"51f7c53f",
X"83e2ac08",
X"810583e2",
X"ac0c8d3d",
X"33cf1170",
X"81ff0651",
X"56567482",
X"26879938",
X"758e0680",
X"dddc5255",
X"8ff73f74",
X"5280dcbc",
X"518fee3f",
X"7483e0a4",
X"082e8b38",
X"74832486",
X"387483e0",
X"a40c8075",
X"248d3874",
X"842983e2",
X"c4055574",
X"088b3880",
X"dde4518f",
X"c43f86e2",
X"3983e0a4",
X"08842983",
X"e2c40570",
X"08028805",
X"b1053352",
X"5b557480",
X"d22e81fe",
X"387480d2",
X"24893874",
X"bf2e8e38",
X"86a93974",
X"80d32e80",
X"e938869f",
X"3980ddf8",
X"518f863f",
X"02b30533",
X"70882b81",
X"fe800602",
X"8805b205",
X"33710551",
X"565688b0",
X"3f80c151",
X"87e43ff5",
X"943f860b",
X"83e0a834",
X"815283e0",
X"a851899f",
X"3f8151fd",
X"c43f748d",
X"38860b83",
X"e2c00c80",
X"dcc8518b",
X"39a80b83",
X"e2c00c80",
X"dcd0518e",
X"b43f83e2",
X"c0085280",
X"dcbc518e",
X"a83f80de",
X"80518ea1",
X"3f87e13f",
X"80c15187",
X"953ff4c5",
X"3f980b83",
X"e2b43383",
X"e2b53371",
X"882b0757",
X"59567481",
X"802e0981",
X"069a3883",
X"e2b23383",
X"e2b33371",
X"882b0756",
X"57ad8075",
X"27883881",
X"98568339",
X"b8567583",
X"e0a834ff",
X"0b83e0a9",
X"34e00b83",
X"e0aa3480",
X"0b83e0ab",
X"34845283",
X"e0a85188",
X"8a3f8451",
X"fcaf3f83",
X"e0a83352",
X"80dcbc51",
X"8daf3f80",
X"de885184",
X"b43902b3",
X"05337088",
X"2b81fe80",
X"06028805",
X"b2053358",
X"77055959",
X"80705d59",
X"86ce3f80",
X"c1518682",
X"3f80de90",
X"518cfe3f",
X"775280dc",
X"bc518cf5",
X"3f80ded4",
X"518cee3f",
X"83e2bc08",
X"792e8381",
X"3883e2d8",
X"0880fc05",
X"5580fd52",
X"7451b895",
X"3f83e080",
X"0880dd80",
X"525b8cc9",
X"3f778224",
X"b93880de",
X"98518cbd",
X"3fff1870",
X"872b83ff",
X"ff800680",
X"e1d80583",
X"e0a85957",
X"55818055",
X"75708105",
X"57337770",
X"81055934",
X"ff157081",
X"ff065155",
X"74ea3882",
X"9b397782",
X"e82e0981",
X"068b3880",
X"dea0518b",
X"fc3f81aa",
X"397782e9",
X"2e098106",
X"81b13880",
X"deb0518b",
X"e83f7858",
X"77873270",
X"30707207",
X"80257a8a",
X"32703070",
X"72078025",
X"73075354",
X"5a515755",
X"75802e97",
X"38787826",
X"9238a00b",
X"83e0a81a",
X"34811970",
X"81ff065a",
X"55eb3981",
X"187081ff",
X"0659558a",
X"7827ffbc",
X"388f5883",
X"e0a31833",
X"83e0a819",
X"34ff1870",
X"81ff0659",
X"55778426",
X"ea389058",
X"800b83e0",
X"a8193481",
X"187081ff",
X"0670982b",
X"52595574",
X"8025e938",
X"80c6557a",
X"858f2484",
X"3880c255",
X"7483e0a8",
X"3480f10b",
X"83e0ab34",
X"810b83e0",
X"ac347a83",
X"e0a9347a",
X"882c5574",
X"83e0aa34",
X"80ce3982",
X"f0782580",
X"c73880de",
X"b8518ab1",
X"3f7780fd",
X"29fd97d3",
X"05527951",
X"8d823f8f",
X"3df40554",
X"80fd5383",
X"e0a85279",
X"518c9e3f",
X"7b811959",
X"567580fc",
X"24833878",
X"5877882c",
X"557483e1",
X"a5347783",
X"e1a63475",
X"83e1a734",
X"80dec051",
X"89eb3f81",
X"805980d8",
X"3983e2d4",
X"08578378",
X"259b3883",
X"e2b43383",
X"e2b53371",
X"882b07fc",
X"1a712979",
X"05838005",
X"5951598d",
X"39778180",
X"2917ff80",
X"05578180",
X"59765280",
X"dcbc5189",
X"ac3f80dc",
X"9c5189a5",
X"3f765279",
X"518bfd3f",
X"8f3df405",
X"54785383",
X"e0a85279",
X"518b9a3f",
X"7851f7fd",
X"3f80decc",
X"5189823f",
X"805280dc",
X"bc5188f9",
X"3f80dc9c",
X"5188f23f",
X"82f73f80",
X"fb3f8b39",
X"83e2a808",
X"810583e2",
X"a80c8f3d",
X"0d04f8b1",
X"3fed8b3f",
X"f939fe3d",
X"0d80e0f4",
X"08703370",
X"81ff0670",
X"842a8132",
X"81065551",
X"52537180",
X"2e8c38a8",
X"733480e0",
X"f40851b8",
X"71347183",
X"e0800c84",
X"3d0d04fe",
X"3d0d80e0",
X"f4087033",
X"7081ff06",
X"70852a81",
X"32810655",
X"51525371",
X"802e8c38",
X"98733480",
X"e0f40851",
X"b8713471",
X"83e0800c",
X"843d0d04",
X"803d0d80",
X"e0f00851",
X"93713480",
X"e0fc0851",
X"ff713482",
X"3d0d04fe",
X"3d0d0293",
X"053380e0",
X"f0085353",
X"8072348a",
X"51ea913f",
X"d33f80e1",
X"80085280",
X"f8723480",
X"e1980852",
X"807234fa",
X"1380e1a0",
X"08535372",
X"723480e1",
X"88085280",
X"723480e1",
X"90085272",
X"723480e0",
X"f4085280",
X"723480e0",
X"f40852b8",
X"7234843d",
X"0d04ff3d",
X"0d028f05",
X"3380e0f8",
X"08525271",
X"7134fe9e",
X"3f83e080",
X"08802ef6",
X"38833d0d",
X"04803d0d",
X"8439eb92",
X"3ffeb83f",
X"83e08008",
X"802ef338",
X"80e0f808",
X"70337081",
X"ff0683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"e0f00851",
X"a3713480",
X"e0fc0851",
X"ff713480",
X"e0f40851",
X"a8713480",
X"e0f40851",
X"b8713482",
X"3d0d0480",
X"3d0d80e0",
X"f0087033",
X"7081c006",
X"70307080",
X"2583e080",
X"0c515151",
X"51823d0d",
X"04ff3d0d",
X"80e0f408",
X"70337081",
X"ff067083",
X"2a813270",
X"81065151",
X"51525270",
X"802ee538",
X"b0723480",
X"e0f40851",
X"b8713483",
X"3d0d0480",
X"3d0d80e1",
X"a8087008",
X"810683e0",
X"800c5182",
X"3d0d04fd",
X"3d0d7577",
X"54548073",
X"25943873",
X"70810555",
X"335280de",
X"d851859d",
X"3fff1353",
X"e939853d",
X"0d04f63d",
X"0d7c7e60",
X"625a5d5b",
X"56805981",
X"55853974",
X"7a295574",
X"527551b0",
X"b83f83e0",
X"80087a27",
X"ee387480",
X"2e80dd38",
X"74527551",
X"b0a33f83",
X"e0800875",
X"53765254",
X"b0ca3f83",
X"e080087a",
X"53755256",
X"b08b3f83",
X"e0800879",
X"30707b07",
X"9f2a7077",
X"80240751",
X"51545572",
X"873883e0",
X"8008c538",
X"768118b0",
X"16555858",
X"8974258b",
X"38b71453",
X"7a853880",
X"d7145372",
X"78348119",
X"59ff9f39",
X"8077348c",
X"3d0d04f7",
X"3d0d7b7d",
X"7f620290",
X"05bb0533",
X"5759565a",
X"5ab05872",
X"8338a058",
X"75707081",
X"05523371",
X"59545590",
X"39807425",
X"8e38ff14",
X"77708105",
X"59335454",
X"72ef3873",
X"ff155553",
X"80732589",
X"38775279",
X"51782def",
X"39753375",
X"57537280",
X"2e903872",
X"52795178",
X"2d757081",
X"05573353",
X"ed398b3d",
X"0d04ee3d",
X"0d646669",
X"69707081",
X"0552335b",
X"4a5c5e5e",
X"76802e82",
X"f93876a5",
X"2e098106",
X"82e03880",
X"70416770",
X"70810552",
X"33714a59",
X"575f76b0",
X"2e098106",
X"8c387570",
X"81055733",
X"76485781",
X"5fd01756",
X"75892680",
X"da387667",
X"5c59805c",
X"9339778a",
X"2480c338",
X"7b8a2918",
X"7b708105",
X"5d335a5c",
X"d0197081",
X"ff065858",
X"897727a4",
X"38ff9f19",
X"7081ff06",
X"ffa91b5a",
X"51568576",
X"279238ff",
X"bf197081",
X"ff065156",
X"7585268a",
X"38c91958",
X"778025ff",
X"b9387a47",
X"7b407881",
X"ff065776",
X"80e42e80",
X"e5387680",
X"e424a738",
X"7680d82e",
X"81863876",
X"80d82490",
X"3876802e",
X"81cc3876",
X"a52e81b6",
X"3881b939",
X"7680e32e",
X"818c3881",
X"af397680",
X"f52e9b38",
X"7680f524",
X"8b387680",
X"f32e8181",
X"38819939",
X"7680f82e",
X"80ca3881",
X"8f39913d",
X"70555780",
X"538a5279",
X"841b7108",
X"535b56fc",
X"813f7655",
X"ab397984",
X"1b710894",
X"3d705b5b",
X"525b5675",
X"80258c38",
X"753056ad",
X"78340280",
X"c1055776",
X"5480538a",
X"527551fb",
X"d53f7755",
X"7e54b839",
X"913d7055",
X"7780d832",
X"70307080",
X"25565158",
X"56905279",
X"841b7108",
X"535b57fb",
X"b13f7555",
X"db397984",
X"1b831233",
X"545b5698",
X"3979841b",
X"7108575b",
X"5680547f",
X"537c527d",
X"51fc9c3f",
X"87397652",
X"7d517c2d",
X"66703358",
X"810547fd",
X"8339943d",
X"0d047283",
X"e0900c71",
X"83e0940c",
X"04fb3d0d",
X"883d7070",
X"84055208",
X"57547553",
X"83e09008",
X"5283e094",
X"0851fcc6",
X"3f873d0d",
X"04ff3d0d",
X"73700853",
X"51029305",
X"33723470",
X"08810571",
X"0c833d0d",
X"04fc3d0d",
X"873d8811",
X"557854a8",
X"f55351fc",
X"993f8052",
X"873d51d1",
X"3f863d0d",
X"04803d0d",
X"72517080",
X"2e833881",
X"517083e0",
X"800c823d",
X"0d04ff3d",
X"0d028f05",
X"33703070",
X"9f2a83e0",
X"800c5252",
X"833d0d04",
X"fd3d0d75",
X"705254a2",
X"913f83e0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee38ff",
X"13537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83e0",
X"8008732e",
X"9e3883e0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb3980",
X"7434853d",
X"0d04803d",
X"0d7251ff",
X"933f823d",
X"0d04ff3d",
X"0d735283",
X"e2dc0872",
X"2e8b3871",
X"5193e23f",
X"7183e2dc",
X"0c833d0d",
X"04fc3d0d",
X"7651df3f",
X"863dfc05",
X"5302a205",
X"22527751",
X"95813f79",
X"863d2271",
X"0c5483e0",
X"800851fe",
X"a43f863d",
X"0d04fc3d",
X"0d7651ff",
X"b53f863d",
X"fc055302",
X"a2052252",
X"775196df",
X"3f79863d",
X"22710c54",
X"83e08008",
X"51fdfa3f",
X"863d0d04",
X"ff3d0d73",
X"51ff8b3f",
X"745199b6",
X"3f7151fd",
X"e43f833d",
X"0d04803d",
X"0d72bc11",
X"0883e080",
X"0c51823d",
X"0d0480c0",
X"0b83e080",
X"0c04fd3d",
X"0d757771",
X"54705354",
X"549fe33f",
X"80c01408",
X"bc140c72",
X"5192be3f",
X"7283e2dc",
X"0c83e080",
X"0851fda1",
X"3f853d0d",
X"04ff3d0d",
X"80dee051",
X"fcbf3f73",
X"83e2e00c",
X"7483e2fc",
X"0c80deec",
X"51fcae3f",
X"a0a73f83",
X"e0800881",
X"ff0680de",
X"fc5252fc",
X"9c3f7180",
X"2e883871",
X"51fcfb3f",
X"a03980df",
X"8c51fc89",
X"3f83e394",
X"518de33f",
X"83e08008",
X"80df9852",
X"52fbf63f",
X"7151fcc5",
X"3f833d0d",
X"04f83d0d",
X"7a598057",
X"80cc5283",
X"e2fc0851",
X"a79b3f83",
X"e0800880",
X"dfa85258",
X"fbcf3f78",
X"5283e380",
X"5199dd3f",
X"83e08008",
X"772e8d38",
X"80dfb451",
X"fbb73f76",
X"5581e639",
X"80dfbc51",
X"fbab3f81",
X"b03983e2",
X"ec337082",
X"2a708106",
X"51565674",
X"819f3875",
X"812a7081",
X"06515574",
X"81933876",
X"883883e2",
X"e008579d",
X"3977802e",
X"819d3880",
X"c8170853",
X"765280df",
X"c051faed",
X"3f80c817",
X"08ff1959",
X"57775376",
X"5280dfcc",
X"51fada3f",
X"83e2ec33",
X"70842a81",
X"0680c419",
X"0c83e2ed",
X"5380e08c",
X"5256fac1",
X"3f785276",
X"519db73f",
X"76519dce",
X"3f83e080",
X"081755af",
X"75708105",
X"573474bc",
X"180c83e2",
X"ed527451",
X"9d983f83",
X"e2e40880",
X"c0180c80",
X"cc177080",
X"c8190c54",
X"80c01708",
X"5383e2e4",
X"085280df",
X"d851f9f9",
X"3f83e2e4",
X"5283e380",
X"5199933f",
X"83e08008",
X"8a3883e2",
X"ed335574",
X"feb83880",
X"dfe451f9",
X"d83f800b",
X"80c8180c",
X"83e2e008",
X"557483e0",
X"800c8a3d",
X"0d04f03d",
X"0d627052",
X"54fab93f",
X"83e08008",
X"7453873d",
X"70535555",
X"fad93f73",
X"53745280",
X"dff851f9",
X"a03f7351",
X"fdaf3f83",
X"e0800854",
X"83e08008",
X"802eb138",
X"bc140852",
X"80e08c51",
X"f9833fbc",
X"14085274",
X"519bb73f",
X"83e08008",
X"8f386352",
X"7351fbfa",
X"3f83e080",
X"08548b39",
X"80c81408",
X"5473d138",
X"81547383",
X"e0800c92",
X"3d0d0471",
X"83e0800c",
X"04803d0d",
X"72bc1108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"7280c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7280c8",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7280",
X"c4110883",
X"e0800c51",
X"823d0d04",
X"f63d0d7c",
X"83e09808",
X"59598179",
X"2782a938",
X"78881908",
X"2782a138",
X"77335675",
X"822e819b",
X"38758224",
X"89387581",
X"2e8d3882",
X"8b397583",
X"2e81b738",
X"82823978",
X"83ffff06",
X"70812a11",
X"7083ffff",
X"067083ff",
X"0671892a",
X"903d5f52",
X"5a515155",
X"7683ff2e",
X"8e388254",
X"76538c18",
X"08155279",
X"51a93975",
X"5476538c",
X"18081552",
X"79519bc5",
X"3f83e080",
X"0881bd38",
X"755483e0",
X"8008538c",
X"18081581",
X"05528c3d",
X"fd05519b",
X"a83f83e0",
X"800881a0",
X"3802a905",
X"338c3d33",
X"71882b07",
X"7a810671",
X"842a5357",
X"58567486",
X"38769fff",
X"06567555",
X"81803975",
X"54781083",
X"fe065378",
X"882a8c19",
X"0805528c",
X"3dfc0551",
X"9ae73f83",
X"e0800880",
X"df3802a9",
X"05338c3d",
X"3371882b",
X"07565780",
X"d1398454",
X"78822b83",
X"fc065378",
X"872a8c19",
X"0805528c",
X"3dfc0551",
X"9ab73f83",
X"e08008b0",
X"3802ab05",
X"33028405",
X"aa053371",
X"982b7190",
X"2b07028c",
X"05a90533",
X"70882b72",
X"07903d33",
X"7180ffff",
X"fe800607",
X"51525357",
X"58568339",
X"81557483",
X"e0800c8c",
X"3d0d04fb",
X"3d0d83e0",
X"9808fe19",
X"881208fe",
X"05555654",
X"80567473",
X"278d3882",
X"14337571",
X"29941608",
X"05575375",
X"83e0800c",
X"873d0d04",
X"fc3d0d76",
X"83e09808",
X"55558075",
X"23881508",
X"5372812e",
X"88388814",
X"08732685",
X"388152b2",
X"39729038",
X"73335271",
X"832e0981",
X"06853890",
X"14085372",
X"8c160c72",
X"802e8d38",
X"7251ff93",
X"3f83e080",
X"08528539",
X"90140852",
X"7190160c",
X"80527183",
X"e0800c86",
X"3d0d04fa",
X"3d0d7883",
X"e0980871",
X"22810570",
X"83ffff06",
X"57545755",
X"73802e88",
X"38901508",
X"53728638",
X"835280e7",
X"39738f06",
X"527180da",
X"38811390",
X"160c8c15",
X"08537290",
X"38830b84",
X"17225752",
X"73762780",
X"c638bf39",
X"821633ff",
X"0574842a",
X"065271b2",
X"387251fb",
X"db3f8152",
X"7183e080",
X"0827a838",
X"835283e0",
X"80088817",
X"08279c38",
X"83e08008",
X"8c160c83",
X"e0800851",
X"fdf93f83",
X"e0800890",
X"160c7375",
X"23805271",
X"83e0800c",
X"883d0d04",
X"f23d0d60",
X"6264585d",
X"5b753355",
X"74a02e09",
X"81068838",
X"81167044",
X"56ef3962",
X"70335656",
X"74af2e09",
X"81068438",
X"81164380",
X"0b881c0c",
X"62703351",
X"5574a026",
X"91387a51",
X"fdd23f83",
X"e0800856",
X"807c3483",
X"a839933d",
X"841c0870",
X"585a5f8a",
X"55a07670",
X"81055834",
X"ff155574",
X"ff2e0981",
X"06ef3880",
X"70595d88",
X"7f085f5a",
X"7c811e70",
X"81ff0660",
X"13703370",
X"af327030",
X"a0732771",
X"80250751",
X"51525b53",
X"5f575574",
X"80d83876",
X"ae2e0981",
X"06833881",
X"55777a27",
X"75075574",
X"802e9f38",
X"79883270",
X"3078ae32",
X"70307073",
X"079f2a53",
X"51575156",
X"75ac3888",
X"588b5aff",
X"ab39ff9f",
X"17557499",
X"268938e0",
X"177081ff",
X"06585577",
X"81197081",
X"ff06721c",
X"535a5755",
X"767534ff",
X"87397c1e",
X"7f0c8055",
X"76a02683",
X"38815574",
X"8b1a347a",
X"51fc913f",
X"83e08008",
X"80f538a0",
X"547a2270",
X"852b83e0",
X"06545590",
X"1b08527b",
X"5195be3f",
X"83e08008",
X"5783e080",
X"08818238",
X"7b335574",
X"802e80f5",
X"388b1c33",
X"70832a70",
X"81065156",
X"5674b438",
X"8b7c841d",
X"0883e080",
X"08595b5b",
X"58ff1858",
X"77ff2e9a",
X"38797081",
X"055b3379",
X"7081055b",
X"33717131",
X"52565675",
X"802ee238",
X"86397580",
X"2ebc387a",
X"51fbf43f",
X"ff863983",
X"e0800856",
X"83e08008",
X"802ea938",
X"83e08008",
X"832e0981",
X"0680de38",
X"841b088b",
X"11335155",
X"7480d238",
X"845680cd",
X"398356ec",
X"39815680",
X"c4397656",
X"841b088b",
X"11335155",
X"74b7388b",
X"1c337084",
X"2a708106",
X"51565774",
X"802ed538",
X"951c3394",
X"1d337198",
X"2b71902b",
X"079b1f33",
X"7f9a0533",
X"71882b07",
X"72077f88",
X"050c5a58",
X"5658fcda",
X"397583e0",
X"800c903d",
X"0d04f83d",
X"0d7a7c59",
X"57825483",
X"fe537752",
X"765193cd",
X"3f835683",
X"e0800880",
X"ec388117",
X"33773371",
X"882b0756",
X"56825674",
X"82d4d52e",
X"09810680",
X"d4387554",
X"b6537752",
X"765193a1",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"ac388254",
X"80d25377",
X"52765192",
X"f83f83e0",
X"80089838",
X"81173377",
X"3371882b",
X"0783e080",
X"08525656",
X"748182c6",
X"2e833881",
X"567583e0",
X"800c8a3d",
X"0d04ec3d",
X"0d665980",
X"0b83e098",
X"0c785678",
X"802e83e8",
X"3892863f",
X"83e08008",
X"81065582",
X"567483d8",
X"38747553",
X"8e3d7053",
X"5858fec2",
X"3f83e080",
X"0881ff06",
X"5675812e",
X"09810680",
X"d4389054",
X"83be5374",
X"52765192",
X"843f83e0",
X"800880c9",
X"388e3d33",
X"5574802e",
X"80c93802",
X"bb053302",
X"8405ba05",
X"3371982b",
X"71902b07",
X"028c05b9",
X"05337088",
X"2b720794",
X"3d337107",
X"70587c57",
X"54525d57",
X"5956fde6",
X"3f83e080",
X"0881ff06",
X"5675832e",
X"09810686",
X"38815682",
X"db397580",
X"2e863887",
X"5682d139",
X"a4548d53",
X"77527651",
X"919b3f81",
X"5683e080",
X"0882bd38",
X"02ba0533",
X"028405b9",
X"05337188",
X"2b07585c",
X"76ab3802",
X"80ca0533",
X"02840580",
X"c9053371",
X"982b7190",
X"2b07963d",
X"3370882b",
X"72070294",
X"0580c705",
X"33710754",
X"525d5758",
X"5602b305",
X"33777129",
X"028805b2",
X"0533028c",
X"05b10533",
X"71882b07",
X"701c708c",
X"1f0c5e59",
X"57585c8d",
X"3d33821a",
X"3402b505",
X"338f3d33",
X"71882b07",
X"595b7784",
X"1a2302b7",
X"05330284",
X"05b60533",
X"71882b07",
X"565b74ab",
X"380280c6",
X"05330284",
X"0580c505",
X"3371982b",
X"71902b07",
X"953d3370",
X"882b7207",
X"02940580",
X"c3053371",
X"07515253",
X"575d5b74",
X"76317731",
X"78842a8f",
X"3d335471",
X"71315356",
X"5696da3f",
X"83e08008",
X"82057088",
X"1b0c709f",
X"f6268105",
X"575583ff",
X"f6752783",
X"38835675",
X"79347583",
X"2e098106",
X"af380280",
X"d2053302",
X"840580d1",
X"05337198",
X"2b71902b",
X"07983d33",
X"70882b72",
X"07029405",
X"80cf0533",
X"7107901f",
X"0c525d57",
X"59568639",
X"761a901a",
X"0c841922",
X"8c1a0818",
X"71842a05",
X"941b0c5c",
X"800b811a",
X"347883e0",
X"980c8056",
X"7583e080",
X"0c963d0d",
X"04e93d0d",
X"83e09808",
X"56865475",
X"802e81a6",
X"38800b81",
X"1734993d",
X"e011466a",
X"54c01153",
X"ec0551f6",
X"cf3f83e0",
X"80085483",
X"e0800881",
X"8538893d",
X"33547380",
X"2e933802",
X"ab053370",
X"842a7081",
X"06515555",
X"73802e86",
X"38835480",
X"e53902b5",
X"05338f3d",
X"3371982b",
X"71902b07",
X"028c05bb",
X"05330290",
X"05ba0533",
X"71882b07",
X"7207a01b",
X"0c029005",
X"bf053302",
X"9405be05",
X"3371982b",
X"71902b07",
X"029c05bd",
X"05337088",
X"2b720799",
X"3d337107",
X"7f9c050c",
X"5283e080",
X"08981f0c",
X"565a5252",
X"53575957",
X"810b8117",
X"3483e080",
X"08547383",
X"e0800c99",
X"3d0d04f5",
X"3d0d7d60",
X"028805ba",
X"05227283",
X"e098085b",
X"5d5a5c5c",
X"807b2386",
X"5676802e",
X"81e03881",
X"17338106",
X"55855674",
X"802e81d2",
X"389c1708",
X"98180831",
X"55747827",
X"87387483",
X"ffff0658",
X"77802e81",
X"ae389817",
X"087083ff",
X"06565674",
X"80ca3882",
X"1733ff05",
X"76892a06",
X"7081ff06",
X"5a5578a0",
X"38758738",
X"a0170855",
X"8d39a417",
X"0851efe0",
X"3f83e080",
X"08558175",
X"2780f838",
X"74a4180c",
X"a4170851",
X"f28d3f83",
X"e0800880",
X"2e80e438",
X"83e08008",
X"19a8180c",
X"98170883",
X"ff068480",
X"71317083",
X"ffff0658",
X"51557776",
X"27833877",
X"56755498",
X"170883ff",
X"0653a817",
X"08527955",
X"7b83387b",
X"5574518b",
X"c03f83e0",
X"8008a438",
X"98170816",
X"98180c75",
X"1a787731",
X"7083ffff",
X"067d2279",
X"05525a56",
X"5a747b23",
X"fece3980",
X"56883980",
X"0b811834",
X"81567583",
X"e0800c8d",
X"3d0d04f7",
X"3d0d7d02",
X"8405b205",
X"227d83e0",
X"9808595a",
X"58598079",
X"23865475",
X"802e82d1",
X"38811633",
X"70810654",
X"55855472",
X"802e82c1",
X"3874862a",
X"5376a838",
X"72810653",
X"72802e8f",
X"38765276",
X"518b883f",
X"83e08008",
X"829c3881",
X"163381bf",
X"06537281",
X"17347654",
X"82933972",
X"81065372",
X"8a389816",
X"08fc8006",
X"98170c9c",
X"16089817",
X"08315372",
X"77278738",
X"7283ffff",
X"06577680",
X"2e81df38",
X"98160870",
X"83ff0654",
X"547280e3",
X"38821633",
X"ff057489",
X"2a067081",
X"ff065653",
X"74a03873",
X"8738a016",
X"08548d39",
X"a4160851",
X"ed9a3f83",
X"e0800854",
X"81742781",
X"a93873a4",
X"170ca416",
X"0851efc7",
X"3f83e080",
X"08802e81",
X"953883e0",
X"80081570",
X"a8180c52",
X"805189eb",
X"3f83e080",
X"0880ff38",
X"81163380",
X"c0075372",
X"8117349a",
X"162283ff",
X"06848071",
X"317083ff",
X"ff065751",
X"53767527",
X"83387655",
X"74527751",
X"89b93f83",
X"e0800880",
X"cd389816",
X"08157098",
X"180c7519",
X"78773170",
X"83ffff06",
X"7c227905",
X"525a5659",
X"53737923",
X"7283ff06",
X"5372febe",
X"3883e080",
X"085283e0",
X"80085188",
X"fe3f83e0",
X"80089338",
X"81163381",
X"bf065372",
X"811734fe",
X"9d398054",
X"8839800b",
X"81173481",
X"547383e0",
X"800c8b3d",
X"0d04fa3d",
X"0d7883e0",
X"98085556",
X"86557380",
X"2e81dc38",
X"81143381",
X"06538555",
X"72802e81",
X"ce389c14",
X"08537276",
X"27833872",
X"56981408",
X"57800b98",
X"150c7580",
X"2e81a938",
X"82143370",
X"892b5653",
X"76802eb5",
X"387452ff",
X"16518ed1",
X"3f83e080",
X"08ff1876",
X"54705358",
X"538ec23f",
X"83e08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b4387251",
X"eaca3f83",
X"e0800853",
X"810b83e0",
X"80082780",
X"cb3883e0",
X"80088815",
X"082780c0",
X"3883e080",
X"08a4150c",
X"98140815",
X"98150c75",
X"753156c9",
X"39981408",
X"16709816",
X"0c735256",
X"ecd13f83",
X"e0800880",
X"2e963882",
X"1433ff05",
X"76892a06",
X"83e08008",
X"05a8150c",
X"80558839",
X"800b8115",
X"34815574",
X"83e0800c",
X"883d0d04",
X"ee3d0d64",
X"56865583",
X"e0980880",
X"2e80f638",
X"943df411",
X"84180c66",
X"54d40552",
X"7551eea0",
X"3f83e080",
X"085583e0",
X"800880cf",
X"38893d33",
X"5473802e",
X"bc3802ab",
X"05337084",
X"2a708106",
X"51555584",
X"5573802e",
X"bc3802b5",
X"05338f3d",
X"3371982b",
X"71902b07",
X"028c05bb",
X"05330290",
X"05ba0533",
X"71882b07",
X"7207881b",
X"0c535759",
X"577551eb",
X"db3f83e0",
X"80085574",
X"832e0981",
X"06833884",
X"557483e0",
X"800c943d",
X"0d04eb3d",
X"0d67695b",
X"59865583",
X"e0980880",
X"2e82fe38",
X"973df405",
X"841a0c79",
X"98387851",
X"eba23f83",
X"e0800855",
X"82e73981",
X"5580f739",
X"835580f2",
X"398c3d58",
X"83559019",
X"08802e80",
X"e538a054",
X"78227085",
X"2b83e006",
X"54569019",
X"08527751",
X"84b73f83",
X"e08008cf",
X"38773356",
X"75802ecc",
X"388b1833",
X"bf067681",
X"e5327030",
X"709f2a51",
X"51565775",
X"ae2e9338",
X"74802e8e",
X"3876832a",
X"70810651",
X"5574802e",
X"ad387851",
X"eb8d3f83",
X"e0800855",
X"83e08008",
X"89389019",
X"08ff9f38",
X"8639800b",
X"901a0c74",
X"832e0981",
X"068d3880",
X"0b901a0c",
X"8a3983e0",
X"80085574",
X"81cf3889",
X"1a579019",
X"08802e81",
X"a5388056",
X"75187033",
X"515574a0",
X"2ea03874",
X"852e0981",
X"06843881",
X"e5557477",
X"70810559",
X"34811670",
X"81ff0657",
X"55877627",
X"d7388818",
X"335574a0",
X"2ea938ae",
X"77708105",
X"59348856",
X"75187033",
X"515574a0",
X"2e953874",
X"77708105",
X"59348116",
X"7081ff06",
X"57558a76",
X"27e2388b",
X"1833881b",
X"349f1833",
X"9e193371",
X"982b7190",
X"2b079d1b",
X"3370882b",
X"72079c1d",
X"3371077f",
X"0c52991c",
X"33981d33",
X"71882b07",
X"53515357",
X"5c567484",
X"1b239718",
X"33961933",
X"71882b07",
X"56567486",
X"1b238077",
X"347851e9",
X"a63f83e0",
X"80085583",
X"e0800883",
X"2e098106",
X"8838800b",
X"901a0c80",
X"557483e0",
X"800c973d",
X"0d04fd3d",
X"0d757753",
X"54733351",
X"70893871",
X"33517080",
X"2ea13873",
X"33723352",
X"53727127",
X"8538ff51",
X"94397073",
X"27853881",
X"518b3981",
X"14811353",
X"54d33980",
X"517083e0",
X"800c853d",
X"0d04fe3d",
X"0d747653",
X"53717081",
X"05533351",
X"70737081",
X"05553470",
X"f038843d",
X"0d04fe3d",
X"0d745280",
X"72335253",
X"70732e8d",
X"38811281",
X"14713353",
X"545270f5",
X"387283e0",
X"800c843d",
X"0d04fc3d",
X"0d765574",
X"83e3c008",
X"2eaf3880",
X"53745184",
X"e03f83e0",
X"800881ff",
X"06ff1470",
X"81ff0672",
X"30709f2a",
X"51525553",
X"5472802e",
X"843871dd",
X"3873fe38",
X"7483e3c0",
X"0c863d0d",
X"04ff3d0d",
X"80e09051",
X"dbfb3fff",
X"0b83e3c0",
X"0c829a3f",
X"85943f83",
X"e0800881",
X"ff065271",
X"f03880e0",
X"9c51dbdd",
X"3f81863f",
X"7183e080",
X"0c833d0d",
X"04fc3d0d",
X"76028405",
X"a2052202",
X"8805a605",
X"227a5455",
X"5555fef6",
X"3f72802e",
X"a03883e3",
X"d0143375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552dd",
X"39800b83",
X"e0800c86",
X"3d0d0480",
X"3d0d7083",
X"e0800c82",
X"3d0d04ff",
X"3d0d83e3",
X"cc081083",
X"e3c40807",
X"80e1ac08",
X"52710c83",
X"3d0d0480",
X"0b83e3cc",
X"0ce13f04",
X"810b83e3",
X"cc0cd83f",
X"04ed3f04",
X"7183e3c8",
X"0c04803d",
X"0d8051f4",
X"3f810b83",
X"e3cc0c81",
X"0b83e3c4",
X"0cffb83f",
X"823d0d04",
X"803d0d72",
X"30707407",
X"802583e3",
X"c40c51ff",
X"a23f823d",
X"0d04fe3d",
X"0d029305",
X"3380e1b0",
X"0854730c",
X"80e1ac08",
X"52710870",
X"81065151",
X"70f73872",
X"087081ff",
X"0683e080",
X"0c51843d",
X"0d04803d",
X"0d81ff51",
X"cd3f83e0",
X"800881ff",
X"0683e080",
X"0c823d0d",
X"04803d0d",
X"ff883f80",
X"51ff9d3f",
X"823d0d04",
X"ff3d0d83",
X"e3d05281",
X"8051cf3f",
X"83e08008",
X"72708105",
X"5434ff11",
X"7083ffff",
X"06515170",
X"e9388180",
X"51ffb33f",
X"83e08008",
X"72708105",
X"5434ff11",
X"7083ffff",
X"06515170",
X"e8388180",
X"51ff973f",
X"83e08008",
X"72708105",
X"5434ff11",
X"7083ffff",
X"06515170",
X"e8388180",
X"51fefb3f",
X"83e08008",
X"72708105",
X"5434ff11",
X"7083ffff",
X"06515170",
X"e838833d",
X"0d04fd3d",
X"0d760284",
X"05970533",
X"535381ff",
X"54fecf3f",
X"fecc3ffe",
X"c93ffec6",
X"3f7180c0",
X"0751fe92",
X"3f72982a",
X"51fe8b3f",
X"72902a70",
X"81ff0652",
X"52fdff3f",
X"72882a70",
X"81ff0652",
X"52fdf33f",
X"7281ff06",
X"51fdeb3f",
X"819551fd",
X"e53ffe8e",
X"3f83e080",
X"0881ff06",
X"ff157081",
X"ff067030",
X"709f2a51",
X"52565353",
X"7281ff2e",
X"09810684",
X"3871db38",
X"7283e080",
X"0c853d0d",
X"04fd3d0d",
X"8151fd98",
X"3f75892b",
X"529151fe",
X"f13f83e0",
X"800881ff",
X"06705553",
X"72a538fd",
X"c13f83e0",
X"800881ff",
X"06537281",
X"fe2e0981",
X"06ed38fd",
X"d33ffdaa",
X"3ffda73f",
X"8051fce0",
X"3f805473",
X"83e0800c",
X"853d0d04",
X"fe3d0d02",
X"93053353",
X"8151fcc8",
X"3f755272",
X"51fea33f",
X"83e08008",
X"81ff0653",
X"8051fcb4",
X"3f7283e0",
X"800c843d",
X"0d04fd3d",
X"0d81ff53",
X"fce43fff",
X"137081ff",
X"06515372",
X"f3387252",
X"7251ffbc",
X"3f83e080",
X"0881ff06",
X"5381ff54",
X"72812e09",
X"810680e2",
X"3883ffff",
X"548052b7",
X"51ff9d3f",
X"83e08008",
X"81ff0653",
X"72812e09",
X"8106a138",
X"8052a951",
X"ff863f83",
X"e0800881",
X"ff065372",
X"802e8d38",
X"ff147083",
X"ffff0655",
X"5373ca38",
X"80528151",
X"fee63f83",
X"e0800881",
X"ff065381",
X"ff547292",
X"387252bb",
X"51fed13f",
X"84805290",
X"51fec93f",
X"72547383",
X"e0800c85",
X"3d0d04fb",
X"3d0d83e3",
X"d0568151",
X"fb863f77",
X"892b5298",
X"51fcdf3f",
X"83e08008",
X"81ff0670",
X"56547380",
X"d738fbae",
X"3f81fe51",
X"fafc3f84",
X"80537570",
X"81055733",
X"51faef3f",
X"ff137083",
X"ffff0651",
X"5372eb38",
X"fb8c3ffb",
X"893ffb86",
X"3f83e080",
X"0881ff06",
X"709f0654",
X"5572852e",
X"09810698",
X"38faef3f",
X"83e08008",
X"81ff0653",
X"72802ef1",
X"388051fa",
X"9b3f8055",
X"7483e080",
X"0c873d0d",
X"0483e08c",
X"080283e0",
X"8c0cfd3d",
X"0d805383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"05085183",
X"d43f83e0",
X"80087083",
X"e0800c54",
X"853d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cfd3d0d",
X"815383e0",
X"8c088c05",
X"085283e0",
X"8c088805",
X"085183a1",
X"3f83e080",
X"087083e0",
X"800c5485",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"f93d0d80",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"88050880",
X"25b93883",
X"e08c0888",
X"05083083",
X"e08c0888",
X"050c800b",
X"83e08c08",
X"f4050c83",
X"e08c08fc",
X"05088a38",
X"810b83e0",
X"8c08f405",
X"0c83e08c",
X"08f40508",
X"83e08c08",
X"fc050c83",
X"e08c088c",
X"05088025",
X"b93883e0",
X"8c088c05",
X"083083e0",
X"8c088c05",
X"0c800b83",
X"e08c08f0",
X"050c83e0",
X"8c08fc05",
X"088a3881",
X"0b83e08c",
X"08f0050c",
X"83e08c08",
X"f0050883",
X"e08c08fc",
X"050c8053",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"81df3f83",
X"e0800870",
X"83e08c08",
X"f8050c54",
X"83e08c08",
X"fc050880",
X"2e903883",
X"e08c08f8",
X"05083083",
X"e08c08f8",
X"050c83e0",
X"8c08f805",
X"087083e0",
X"800c5489",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"fb3d0d80",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"88050880",
X"25993883",
X"e08c0888",
X"05083083",
X"e08c0888",
X"050c810b",
X"83e08c08",
X"fc050c83",
X"e08c088c",
X"05088025",
X"903883e0",
X"8c088c05",
X"083083e0",
X"8c088c05",
X"0c815383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"050851bd",
X"3f83e080",
X"087083e0",
X"8c08f805",
X"0c5483e0",
X"8c08fc05",
X"08802e90",
X"3883e08c",
X"08f80508",
X"3083e08c",
X"08f8050c",
X"83e08c08",
X"f8050870",
X"83e0800c",
X"54873d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cfd3d",
X"0d810b83",
X"e08c08fc",
X"050c800b",
X"83e08c08",
X"f8050c83",
X"e08c088c",
X"050883e0",
X"8c088805",
X"0827b938",
X"83e08c08",
X"fc050880",
X"2eae3880",
X"0b83e08c",
X"088c0508",
X"24a23883",
X"e08c088c",
X"05081083",
X"e08c088c",
X"050c83e0",
X"8c08fc05",
X"081083e0",
X"8c08fc05",
X"0cffb839",
X"83e08c08",
X"fc050880",
X"2e80e138",
X"83e08c08",
X"8c050883",
X"e08c0888",
X"050826ad",
X"3883e08c",
X"08880508",
X"83e08c08",
X"8c050831",
X"83e08c08",
X"88050c83",
X"e08c08f8",
X"050883e0",
X"8c08fc05",
X"080783e0",
X"8c08f805",
X"0c83e08c",
X"08fc0508",
X"812a83e0",
X"8c08fc05",
X"0c83e08c",
X"088c0508",
X"812a83e0",
X"8c088c05",
X"0cff9539",
X"83e08c08",
X"90050880",
X"2e933883",
X"e08c0888",
X"05087083",
X"e08c08f4",
X"050c5191",
X"3983e08c",
X"08f80508",
X"7083e08c",
X"08f4050c",
X"5183e08c",
X"08f40508",
X"83e0800c",
X"853d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cff3d0d",
X"800b83e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"8106ff11",
X"70097083",
X"e08c088c",
X"05080683",
X"e08c08fc",
X"05081183",
X"e08c08fc",
X"050c83e0",
X"8c088805",
X"08812a83",
X"e08c0888",
X"050c83e0",
X"8c088c05",
X"081083e0",
X"8c088c05",
X"0c515151",
X"5183e08c",
X"08880508",
X"802e8438",
X"ffab3983",
X"e08c08fc",
X"05087083",
X"e0800c51",
X"833d0d83",
X"e08c0c04",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"48656c6c",
X"6f20576f",
X"726c640a",
X"20492061",
X"6d20616e",
X"20417461",
X"7269210a",
X"00000000",
X"44495220",
X"696e6974",
X"206f6b0a",
X"00000000",
X"4f70656e",
X"696e6720",
X"66696c65",
X"0a000000",
X"47554e50",
X"4f574452",
X"2e415452",
X"00000000",
X"46494c45",
X"206f7065",
X"6e206f6b",
X"0a000000",
X"46494c45",
X"206f7065",
X"6e206661",
X"696c6564",
X"0a000000",
X"44495220",
X"696e6974",
X"20666169",
X"6c65640a",
X"00000000",
X"636d643a",
X"00000000",
X"25640000",
X"45525220",
X"00000000",
X"53504446",
X"00000000",
X"53504453",
X"00000000",
X"436f756c",
X"64206e6f",
X"74207265",
X"61642068",
X"65616465",
X"720a0000",
X"58464400",
X"78666400",
X"58464420",
X"00000000",
X"58455820",
X"00000000",
X"41545220",
X"00000000",
X"556e6b6e",
X"6f776e20",
X"66696c65",
X"20747970",
X"65000000",
X"4d442000",
X"53442000",
X"44442000",
X"58442000",
X"42414420",
X"73656374",
X"6f722073",
X"697a6500",
X"300a0000",
X"2873656e",
X"643a0000",
X"3a63686b",
X"3a000000",
X"29000000",
X"44726976",
X"653a0000",
X"44726976",
X"65206e6f",
X"74207072",
X"6573656e",
X"74000000",
X"53706565",
X"643a0000",
X"53746174",
X"3a000000",
X"3a646f6e",
X"650a0000",
X"53656374",
X"6f723a00",
X"626f6f74",
X"20000000",
X"6e756d74",
X"6f627566",
X"66657220",
X"00000000",
X"6e616d65",
X"20000000",
X"64617461",
X"20000000",
X"2073656e",
X"64696e67",
X"0a000000",
X"20726563",
X"65697665",
X"3a000000",
X"25303278",
X"00000000",
X"6469725f",
X"696e6974",
X"0a000000",
X"6469736b",
X"5f696e69",
X"7420676f",
X"0a000000",
X"6469736b",
X"5f696e69",
X"7420646f",
X"6e650a00",
X"70665f6d",
X"6f756e74",
X"0a000000",
X"70665f6d",
X"6f756e74",
X"20646f6e",
X"650a0000",
X"6f70656e",
X"64697220",
X"00000000",
X"4641494c",
X"20000000",
X"4f4b2000",
X"696e6320",
X"25782025",
X"78200000",
X"6e657874",
X"20257820",
X"25642000",
X"6e202564",
X"20256420",
X"25782000",
X"6469725f",
X"656e7472",
X"69657320",
X"646f6e65",
X"20000000",
X"66696c65",
X"6e616d65",
X"3a257320",
X"6469726e",
X"616d653a",
X"25732000",
X"20696e20",
X"696e6974",
X"20000000",
X"20736574",
X"74696e67",
X"20667265",
X"71200000",
X"00000000",
X"00000000",
X"0001d20f",
X"0001d400",
X"0001d401",
X"0001d409",
X"0001d010",
X"0001d301",
X"0001d300",
X"0001d20a",
X"0001d01b",
X"0001d018",
X"0001d017",
X"0001d01a",
X"0001d403",
X"0001d402",
X"0001d40e",
X"0004007c",
X"00040078",
X"00040074",
X"00040068",
X"00040060",
X"0004005c",
X"00040058",
X"00040054",
X"00040050",
X"0004004c",
X"00040048",
X"00040044",
X"00040040",
X"00040030",
X"0004002c",
X"00040028",
X"00040024",
X"00040020",
X"0004001c",
X"00040018",
X"00040014",
X"00040010",
X"0004000c",
X"00040008",
X"00040004",
X"00040000",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
