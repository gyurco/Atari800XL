
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80dc",
X"e0738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80df",
X"fc0c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580d7",
X"902d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580d5a4",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80cef804",
X"fc3d0d76",
X"705255b3",
X"f33f83e0",
X"800815ff",
X"05547375",
X"2e8e3873",
X"335372ae",
X"2e8638ff",
X"1454ef39",
X"77528114",
X"51b38b3f",
X"83e08008",
X"307083e0",
X"80080780",
X"2583e080",
X"0c53863d",
X"0d04fc3d",
X"0d767052",
X"559aac3f",
X"83e08008",
X"54815383",
X"e0800880",
X"c7387451",
X"99ef3f83",
X"e080080b",
X"0b80dec0",
X"5383e080",
X"085253ff",
X"8f3f83e0",
X"8008a538",
X"0b0b80de",
X"c4527251",
X"fefe3f83",
X"e0800894",
X"380b0b80",
X"dec85272",
X"51feed3f",
X"83e08008",
X"802e8338",
X"81547353",
X"7283e080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"99c53f81",
X"5383e080",
X"08993873",
X"51998e3f",
X"0b0b80de",
X"cc5283e0",
X"800851fe",
X"b33f83e0",
X"80085372",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"70525499",
X"923f8153",
X"83e08008",
X"99387351",
X"98db3f0b",
X"0b80ded0",
X"5283e080",
X"0851fe80",
X"3f83e080",
X"08537283",
X"e0800c85",
X"3d0d04e0",
X"3d0da33d",
X"0870525e",
X"8f863f83",
X"e0800833",
X"943d5654",
X"73943880",
X"e1c85274",
X"5184c639",
X"7d527851",
X"92833f84",
X"d0397d51",
X"8eee3f83",
X"e0800852",
X"74518e9e",
X"3f83e09c",
X"0852933d",
X"70525d94",
X"f33f83e0",
X"80085980",
X"0b83e080",
X"08555b83",
X"e080087b",
X"2e943881",
X"1b74525b",
X"97f43f83",
X"e0800854",
X"83e08008",
X"ee38805a",
X"ff7a437a",
X"427a415f",
X"7909709f",
X"2c7b065b",
X"547a7a24",
X"8438ff1b",
X"5af61a70",
X"09709f2c",
X"72067bff",
X"125a5a52",
X"55558075",
X"25953876",
X"5197b33f",
X"83e08008",
X"76ff1858",
X"55577380",
X"24ed3874",
X"7f2e8638",
X"b8de3f74",
X"5f78ff1b",
X"70585d58",
X"807a2595",
X"38775197",
X"893f83e0",
X"800876ff",
X"18585558",
X"738024ed",
X"38800b83",
X"e3980c80",
X"0b83e3b8",
X"0c0b0b80",
X"ded4518b",
X"e23f8180",
X"0b83e3b8",
X"0c0b0b80",
X"dedc518b",
X"d23fa80b",
X"83e3980c",
X"76802e80",
X"e83883e3",
X"98087779",
X"32703070",
X"72078025",
X"70872b83",
X"e3b80c51",
X"56785356",
X"5696bc3f",
X"83e08008",
X"802e8a38",
X"0b0b80de",
X"e4518b97",
X"3f765195",
X"fc3f83e0",
X"8008520b",
X"0b80df98",
X"518b843f",
X"76519682",
X"3f83e080",
X"0883e398",
X"08555775",
X"74258638",
X"a81656f7",
X"397583e3",
X"980c86f0",
X"7624ff94",
X"3887980b",
X"83e3980c",
X"77802eb7",
X"38775195",
X"b83f83e0",
X"80087852",
X"5595d83f",
X"0b0b80de",
X"ec5483e0",
X"80088f38",
X"87398076",
X"34fd9639",
X"0b0b80de",
X"e8547453",
X"73520b0b",
X"80deb051",
X"8a9d3f80",
X"540b0b80",
X"deb8518a",
X"923f8114",
X"5473a82e",
X"098106ed",
X"38868da0",
X"51b4de3f",
X"8052903d",
X"70525480",
X"c2bc3f83",
X"52735180",
X"c2b43f61",
X"802e80ff",
X"387b5473",
X"ff2e9638",
X"78802e81",
X"80387851",
X"94d83f83",
X"e08008ff",
X"155559e7",
X"3978802e",
X"80eb3878",
X"5194d43f",
X"83e08008",
X"802efc84",
X"38785194",
X"9c3f83e0",
X"8008520b",
X"0b80debc",
X"51abfa3f",
X"83e08008",
X"a4387c51",
X"adb23f83",
X"e0800855",
X"74ff1656",
X"54807425",
X"fbef3874",
X"1d703355",
X"5673af2e",
X"fec838e8",
X"39785193",
X"da3f83e0",
X"8008527c",
X"51ace93f",
X"fbcf397f",
X"88296010",
X"057a0561",
X"055afc80",
X"39a23d0d",
X"04fe3d0d",
X"80e0d008",
X"70337081",
X"ff067084",
X"2a813281",
X"06555152",
X"5371802e",
X"8c38a873",
X"3480e0d0",
X"0851b871",
X"347183e0",
X"800c843d",
X"0d04fe3d",
X"0d80e0d0",
X"08703370",
X"81ff0670",
X"852a8132",
X"81065551",
X"52537180",
X"2e8c3898",
X"733480e0",
X"d00851b8",
X"71347183",
X"e0800c84",
X"3d0d0480",
X"3d0d80e0",
X"cc085193",
X"713480e0",
X"d80851ff",
X"7134823d",
X"0d04fe3d",
X"0d029305",
X"3380e0cc",
X"08535380",
X"72348a51",
X"b2a73fd3",
X"3f80e0dc",
X"085280f8",
X"723480e0",
X"f4085280",
X"7234fa13",
X"80e0fc08",
X"53537272",
X"3480e0e4",
X"08528072",
X"3480e0ec",
X"08527272",
X"3480e0d0",
X"08528072",
X"3480e0d0",
X"0852b872",
X"34843d0d",
X"04ff3d0d",
X"028f0533",
X"80e0d408",
X"52527171",
X"34fe9e3f",
X"83e08008",
X"802ef638",
X"833d0d04",
X"803d0d84",
X"39baf53f",
X"feb83f83",
X"e0800880",
X"2ef33880",
X"e0d40870",
X"337081ff",
X"0683e080",
X"0c515182",
X"3d0d0480",
X"3d0d80e0",
X"cc0851a3",
X"713480e0",
X"d80851ff",
X"713480e0",
X"d00851a8",
X"713480e0",
X"d00851b8",
X"7134823d",
X"0d04803d",
X"0d80e0cc",
X"08703370",
X"81c00670",
X"30708025",
X"83e0800c",
X"51515151",
X"823d0d04",
X"ff3d0d80",
X"e0d00870",
X"337081ff",
X"0670832a",
X"81327081",
X"06515151",
X"52527080",
X"2ee538b0",
X"723480e0",
X"d00851b8",
X"7134833d",
X"0d04803d",
X"0d80e188",
X"08700881",
X"0683e080",
X"0c51823d",
X"0d04fd3d",
X"0d757754",
X"54807325",
X"94387370",
X"81055533",
X"5280def0",
X"5185a03f",
X"ff1353e9",
X"39853d0d",
X"04f63d0d",
X"7c7e6062",
X"5a5d5b56",
X"80598155",
X"8539747a",
X"29557452",
X"755180c0",
X"a13f83e0",
X"80087a27",
X"ed387480",
X"2e80df38",
X"74527551",
X"80c08b3f",
X"83e08008",
X"75537652",
X"5480c0b1",
X"3f83e080",
X"087a5375",
X"5256bff2",
X"3f83e080",
X"08793070",
X"7b079f2a",
X"70778024",
X"07515154",
X"55728738",
X"83e08008",
X"c3387681",
X"18b01655",
X"58588974",
X"258b38b7",
X"14537a85",
X"3880d714",
X"53727834",
X"811959ff",
X"9d398077",
X"348c3d0d",
X"04f73d0d",
X"7b7d7f62",
X"029005bb",
X"05335759",
X"565a5ab0",
X"58728338",
X"a0587570",
X"70810552",
X"33715954",
X"55903980",
X"74258e38",
X"ff147770",
X"81055933",
X"545472ef",
X"3873ff15",
X"55538073",
X"25893877",
X"52795178",
X"2def3975",
X"33755753",
X"72802e90",
X"38725279",
X"51782d75",
X"70810557",
X"3353ed39",
X"8b3d0d04",
X"ee3d0d64",
X"66696970",
X"70810552",
X"335b4a5c",
X"5e5e7680",
X"2e82f938",
X"76a52e09",
X"810682e0",
X"38807041",
X"67707081",
X"05523371",
X"4a59575f",
X"76b02e09",
X"81068c38",
X"75708105",
X"57337648",
X"57815fd0",
X"17567589",
X"2680da38",
X"76675c59",
X"805c9339",
X"778a2480",
X"c3387b8a",
X"29187b70",
X"81055d33",
X"5a5cd019",
X"7081ff06",
X"58588977",
X"27a438ff",
X"9f197081",
X"ff06ffa9",
X"1b5a5156",
X"85762792",
X"38ffbf19",
X"7081ff06",
X"51567585",
X"268a38c9",
X"19587780",
X"25ffb938",
X"7a477b40",
X"7881ff06",
X"577680e4",
X"2e80e538",
X"7680e424",
X"a7387680",
X"d82e8186",
X"387680d8",
X"24903876",
X"802e81cc",
X"3876a52e",
X"81b63881",
X"b9397680",
X"e32e818c",
X"3881af39",
X"7680f52e",
X"9b387680",
X"f5248b38",
X"7680f32e",
X"81813881",
X"99397680",
X"f82e80ca",
X"38818f39",
X"913d7055",
X"5780538a",
X"5279841b",
X"7108535b",
X"56fbfe3f",
X"7655ab39",
X"79841b71",
X"08943d70",
X"5b5b525b",
X"56758025",
X"8c387530",
X"56ad7834",
X"0280c105",
X"57765480",
X"538a5275",
X"51fbd23f",
X"77557e54",
X"b839913d",
X"70557780",
X"d8327030",
X"70802556",
X"51585690",
X"5279841b",
X"7108535b",
X"57fbae3f",
X"7555db39",
X"79841b83",
X"1233545b",
X"56983979",
X"841b7108",
X"575b5680",
X"547f537c",
X"527d51fc",
X"9c3f8739",
X"76527d51",
X"7c2d6670",
X"33588105",
X"47fd8339",
X"943d0d04",
X"7283e090",
X"0c7183e0",
X"940c04fb",
X"3d0d883d",
X"70708405",
X"52085754",
X"755383e0",
X"90085283",
X"e0940851",
X"fcc63f87",
X"3d0d04ff",
X"3d0d7370",
X"08535102",
X"93053372",
X"34700881",
X"05710c83",
X"3d0d04fc",
X"3d0d873d",
X"88115578",
X"5499b753",
X"51fc993f",
X"8052873d",
X"51d13f86",
X"3d0d04fd",
X"3d0d7570",
X"5254a3bc",
X"3f83e080",
X"08145372",
X"742e9238",
X"ff137033",
X"535371af",
X"2e098106",
X"ee388113",
X"537283e0",
X"800c853d",
X"0d04fd3d",
X"0d757770",
X"535454c7",
X"3f83e080",
X"08732ea1",
X"3883e080",
X"08733152",
X"ff125271",
X"ff2e8f38",
X"72708105",
X"54337470",
X"81055634",
X"eb39ff14",
X"54807434",
X"853d0d04",
X"803d0d72",
X"51ff903f",
X"823d0d04",
X"7183e080",
X"0c04803d",
X"0d725180",
X"7134810b",
X"bc120c80",
X"0b80c012",
X"0c823d0d",
X"04800b83",
X"e2c40824",
X"8a38b98b",
X"3fff0b83",
X"e2c40c80",
X"0b83e080",
X"0c04ff3d",
X"0d735283",
X"e0a00872",
X"2e8d38d9",
X"3f715196",
X"913f7183",
X"e0a00c83",
X"3d0d04f4",
X"3d0d7e60",
X"625c5a55",
X"8154bc15",
X"08819138",
X"7451cf3f",
X"7958807a",
X"2580f738",
X"83e2f408",
X"70892a57",
X"83ff0678",
X"84807231",
X"56565773",
X"78258338",
X"73557583",
X"e2c4082e",
X"8438ff89",
X"3f83e2c4",
X"088025a6",
X"3875892b",
X"5198d43f",
X"83e2f408",
X"8f3dfc11",
X"555c5481",
X"52f81b51",
X"96be3f76",
X"1483e2f4",
X"0c7583e2",
X"c40c7453",
X"76527851",
X"b79e3f83",
X"e0800883",
X"e2f40816",
X"83e2f40c",
X"78763176",
X"1b5b5956",
X"778024ff",
X"8b38617a",
X"710c5475",
X"5475802e",
X"83388154",
X"7383e080",
X"0c8e3d0d",
X"04fc3d0d",
X"fe9b3f76",
X"51feaf3f",
X"863dfc05",
X"53785277",
X"5195e13f",
X"7975710c",
X"5483e080",
X"085483e0",
X"8008802e",
X"83388154",
X"7383e080",
X"0c863d0d",
X"04fd3d0d",
X"7683e2c4",
X"08535380",
X"72248938",
X"71732e84",
X"38fdd63f",
X"7551fdea",
X"3f725197",
X"a63f7352",
X"73802e83",
X"38815271",
X"83e0800c",
X"853d0d04",
X"803d0d72",
X"80c01108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"72bc1108",
X"83e0800c",
X"51823d0d",
X"0480c40b",
X"83e0800c",
X"04fd3d0d",
X"75777154",
X"70535553",
X"9f9a3f82",
X"c81308bc",
X"150c82c0",
X"130880c0",
X"150cfcf1",
X"3f735193",
X"a93f7383",
X"e0a00c83",
X"e0800853",
X"83e08008",
X"802e8338",
X"81537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"5553fcc5",
X"3f72802e",
X"a538bc13",
X"08527351",
X"9ea43f83",
X"e080088f",
X"38775272",
X"51ff9a3f",
X"83e08008",
X"538a3982",
X"cc130853",
X"d8398153",
X"7283e080",
X"0c853d0d",
X"04fe3d0d",
X"ff0b83e2",
X"c40c7483",
X"e0a40c75",
X"83e2c00c",
X"b3e83f83",
X"e0800881",
X"ff065281",
X"53719938",
X"83e2dc51",
X"8e933f83",
X"e0800852",
X"83e08008",
X"802e8338",
X"72527153",
X"7283e080",
X"0c843d0d",
X"04fa3d0d",
X"787a82c4",
X"120882c4",
X"12087072",
X"24595656",
X"57577373",
X"2e098106",
X"913880c0",
X"165280c0",
X"17519c95",
X"3f83e080",
X"08557483",
X"e0800c88",
X"3d0d04f6",
X"3d0d7c5b",
X"807b715c",
X"54577a77",
X"2e8c3881",
X"1a82cc14",
X"08545a72",
X"f6388059",
X"80d9397a",
X"54815780",
X"707b7b31",
X"5a5755ff",
X"18537473",
X"2580c138",
X"82cc1408",
X"527351ff",
X"8c3f800b",
X"83e08008",
X"25a13882",
X"cc140882",
X"cc110882",
X"cc160c74",
X"82cc120c",
X"5375802e",
X"86387282",
X"cc170c72",
X"54805773",
X"82cc1508",
X"81175755",
X"56ffb839",
X"81195980",
X"0bff1b54",
X"54787325",
X"83388154",
X"76813270",
X"75065153",
X"72ff9038",
X"8c3d0d04",
X"f73d0d7b",
X"7d5a5a82",
X"d05283e2",
X"c00851b3",
X"b13f83e0",
X"800857f9",
X"e83f7952",
X"83e2c851",
X"95b43f83",
X"e0800854",
X"805383e0",
X"8008732e",
X"09810682",
X"833883e0",
X"a4080b0b",
X"80debc53",
X"7052569b",
X"d33f0b0b",
X"80debc52",
X"80c01651",
X"9bc63f75",
X"bc170c73",
X"82c0170c",
X"810b82c4",
X"170c810b",
X"82c8170c",
X"7382cc17",
X"0cff1782",
X"d0175557",
X"81913983",
X"e0b03370",
X"822a7081",
X"06515455",
X"72818038",
X"74812a81",
X"06587780",
X"f6387484",
X"2a810682",
X"c4150c83",
X"e0b03381",
X"0682c815",
X"0c795273",
X"519aed3f",
X"73519b84",
X"3f83e080",
X"081453af",
X"73708105",
X"553472bc",
X"150c83e0",
X"b1527251",
X"9ace3f83",
X"e0a80882",
X"c0150c83",
X"e0be5280",
X"c014519a",
X"bb3f7880",
X"2e8d3873",
X"51782d83",
X"e0800880",
X"2e993877",
X"82cc150c",
X"75802e86",
X"387382cc",
X"170c7382",
X"d015ff19",
X"59555676",
X"802e9b38",
X"83e0a852",
X"83e2c851",
X"94aa3f83",
X"e080088a",
X"3883e0b1",
X"335372fe",
X"d2387880",
X"2e893883",
X"e0a40851",
X"fcb93f83",
X"e0a40853",
X"7283e080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb63f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f697",
X"3f83e080",
X"08745387",
X"3d705355",
X"55f6b73f",
X"f7973f73",
X"51d33f63",
X"53745283",
X"e0800851",
X"fab93f92",
X"3d0d0471",
X"83e0800c",
X"0480c012",
X"83e0800c",
X"04803d0d",
X"7282c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"e0800c51",
X"823d0d04",
X"f93d0d79",
X"83e09808",
X"57578177",
X"27819638",
X"76881708",
X"27818e38",
X"75335574",
X"822e8938",
X"74832eb3",
X"3880fe39",
X"74547610",
X"83fe0653",
X"76882a8c",
X"17080552",
X"893dfc05",
X"51ae843f",
X"83e08008",
X"80df3802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d13984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"51add43f",
X"83e08008",
X"b038029f",
X"05330284",
X"059e0533",
X"71982b71",
X"902b0702",
X"8c059d05",
X"3370882b",
X"72078d3d",
X"337180ff",
X"fffe8006",
X"07515253",
X"57585683",
X"39815574",
X"83e0800c",
X"893d0d04",
X"fb3d0d83",
X"e09808fe",
X"19881208",
X"fe055556",
X"54805674",
X"73278d38",
X"82143375",
X"71299416",
X"08055753",
X"7583e080",
X"0c873d0d",
X"04fc3d0d",
X"7652800b",
X"83e09808",
X"70335152",
X"5370832e",
X"09810691",
X"38951233",
X"94133371",
X"982b7190",
X"2b075555",
X"519b1233",
X"9a133371",
X"882b0774",
X"0783e080",
X"0c55863d",
X"0d04fc3d",
X"0d7683e0",
X"98085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"fed63f83",
X"e0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183e080",
X"0c863d0d",
X"04fa3d0d",
X"7883e098",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fcb13f",
X"81527183",
X"e0800827",
X"a8388352",
X"83e08008",
X"88170827",
X"9c3883e0",
X"80088c16",
X"0c83e080",
X"0851fdbc",
X"3f83e080",
X"0890160c",
X"73752380",
X"527183e0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585e5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"9f269138",
X"7a51fdd2",
X"3f83e080",
X"0856807d",
X"34838139",
X"933d841c",
X"08705859",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"3880705a",
X"5c887f08",
X"5f5a7b81",
X"1d7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535e57",
X"557480e7",
X"3876ae2e",
X"09810683",
X"38815578",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675bb",
X"3888598b",
X"5affab39",
X"76982b55",
X"74802587",
X"3880dbf0",
X"173357ff",
X"9f175574",
X"99268938",
X"e0177081",
X"ff065855",
X"78811a70",
X"81ff0672",
X"1b535b57",
X"55767534",
X"fef8397b",
X"1e7f0c80",
X"5576a026",
X"83388155",
X"748b1934",
X"7a51fc82",
X"3f83e080",
X"0880f538",
X"a0547a22",
X"70852b83",
X"e0065455",
X"901b0852",
X"7c51a88f",
X"3f83e080",
X"085783e0",
X"80088181",
X"387c3355",
X"74802e80",
X"f4388b1d",
X"3370832a",
X"70810651",
X"565674b4",
X"388b7d84",
X"1d0883e0",
X"8008595b",
X"5b58ff18",
X"5877ff2e",
X"9a387970",
X"81055b33",
X"79708105",
X"5b337171",
X"31525656",
X"75802ee2",
X"38863975",
X"802e9638",
X"7a51fbe5",
X"3fff8639",
X"83e08008",
X"5683e080",
X"08b63883",
X"39765684",
X"1b088b11",
X"33515574",
X"a7388b1d",
X"3370842a",
X"70810651",
X"56567489",
X"38835694",
X"39815690",
X"397c51fa",
X"943f83e0",
X"8008881c",
X"0cfd8139",
X"7583e080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"51a6d43f",
X"835683e0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"51a6a83f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"7651a5ff",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583e080",
X"0c8a3d0d",
X"04eb3d0d",
X"675a800b",
X"83e0980c",
X"a5b43f83",
X"e0800881",
X"06558256",
X"7483ee38",
X"7475538f",
X"3d705357",
X"59feca3f",
X"83e08008",
X"81ff0657",
X"76812e09",
X"810680d4",
X"38905483",
X"be537452",
X"7551a593",
X"3f83e080",
X"0880c938",
X"8f3d3355",
X"74802e80",
X"c93802bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"33710770",
X"587b575e",
X"525e5759",
X"57fdee3f",
X"83e08008",
X"81ff0657",
X"76832e09",
X"81068638",
X"815682f1",
X"3976802e",
X"86388656",
X"82e739a4",
X"548d5378",
X"527551a4",
X"aa3f8156",
X"83e08008",
X"82d33802",
X"be053302",
X"8405bd05",
X"3371882b",
X"07595d77",
X"ab380280",
X"ce053302",
X"840580cd",
X"05337198",
X"2b71902b",
X"07973d33",
X"70882b72",
X"07029405",
X"80cb0533",
X"71075452",
X"5e575956",
X"02b70533",
X"78712902",
X"8805b605",
X"33028c05",
X"b5053371",
X"882b0770",
X"1d707f8c",
X"050c5f59",
X"57595d8e",
X"3d33821b",
X"3402b905",
X"33903d33",
X"71882b07",
X"5a5c7884",
X"1b2302bb",
X"05330284",
X"05ba0533",
X"71882b07",
X"565c74ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"07515253",
X"575e5c74",
X"76317831",
X"79842a90",
X"3d335471",
X"71315356",
X"56a4973f",
X"83e08008",
X"82057088",
X"1c0c83e0",
X"8008e08a",
X"05565674",
X"83dffe26",
X"83388257",
X"83fff676",
X"27853883",
X"57893986",
X"5676802e",
X"80db3876",
X"7a347683",
X"2e098106",
X"b0380280",
X"d6053302",
X"840580d5",
X"05337198",
X"2b71902b",
X"07993d33",
X"70882b72",
X"07029405",
X"80d30533",
X"71077f90",
X"050c525e",
X"57585686",
X"39771b90",
X"1b0c841a",
X"228c1b08",
X"1971842a",
X"05941c0c",
X"5d800b81",
X"1b347983",
X"e0980c80",
X"567583e0",
X"800c973d",
X"0d04e93d",
X"0d83e098",
X"08568554",
X"75802e81",
X"8238800b",
X"81173499",
X"3de01146",
X"6a548a3d",
X"705458ec",
X"0551f6e6",
X"3f83e080",
X"085483e0",
X"800880df",
X"38893d33",
X"5473802e",
X"913802ab",
X"05337084",
X"2a810651",
X"5574802e",
X"86388354",
X"80c13976",
X"51f48a3f",
X"83e08008",
X"a0170c02",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"9c1c0c52",
X"78981b0c",
X"53565957",
X"810b8117",
X"34745473",
X"83e0800c",
X"993d0d04",
X"f53d0d7d",
X"7f617283",
X"e098085a",
X"5d5d595c",
X"807b0c85",
X"5775802e",
X"81e03881",
X"16338106",
X"55845774",
X"802e81d2",
X"38913974",
X"81173486",
X"39800b81",
X"17348157",
X"81c0399c",
X"16089817",
X"08315574",
X"78278338",
X"74587780",
X"2e81a938",
X"98160870",
X"83ff0656",
X"577480cf",
X"38821633",
X"ff057789",
X"2a067081",
X"ff065a55",
X"78a03876",
X"8738a016",
X"08558d39",
X"a4160851",
X"f0ea3f83",
X"e0800855",
X"817527ff",
X"a83874a4",
X"170ca416",
X"0851f284",
X"3f83e080",
X"085583e0",
X"8008802e",
X"ff893883",
X"e0800819",
X"a8170c98",
X"160883ff",
X"06848071",
X"31515577",
X"75278338",
X"77557483",
X"ffff0654",
X"98160883",
X"ff0653a8",
X"16085279",
X"577b8338",
X"7b577651",
X"9ed13f83",
X"e08008fe",
X"d0389816",
X"08159817",
X"0c741a78",
X"76317c08",
X"177d0c59",
X"5afed339",
X"80577683",
X"e0800c8d",
X"3d0d04fa",
X"3d0d7883",
X"e0980855",
X"56855573",
X"802e81e1",
X"38811433",
X"81065384",
X"5572802e",
X"81d3389c",
X"14085372",
X"76278338",
X"72569814",
X"0857800b",
X"98150c75",
X"802e81b7",
X"38821433",
X"70892b56",
X"5376802e",
X"b5387452",
X"ff16519f",
X"993f83e0",
X"8008ff18",
X"76547053",
X"58539f8a",
X"3f83e080",
X"08732696",
X"38743070",
X"78067098",
X"170c7771",
X"31a41708",
X"52585153",
X"8939a014",
X"0870a416",
X"0c537476",
X"27b93872",
X"51eed93f",
X"83e08008",
X"53810b83",
X"e0800827",
X"8b388814",
X"0883e080",
X"08268838",
X"800b8115",
X"34b03983",
X"e08008a4",
X"150c9814",
X"08159815",
X"0c757531",
X"56c43998",
X"14081670",
X"98160c73",
X"5256efc8",
X"3f83e080",
X"088c3883",
X"e0800881",
X"15348155",
X"94398214",
X"33ff0576",
X"892a0683",
X"e0800805",
X"a8150c80",
X"557483e0",
X"800c883d",
X"0d04ef3d",
X"0d635685",
X"5583e098",
X"08802e80",
X"d238933d",
X"f4058417",
X"0c645388",
X"3d705376",
X"5257f1d2",
X"3f83e080",
X"085583e0",
X"8008b438",
X"883d3354",
X"73802ea1",
X"3802a705",
X"3370842a",
X"70810651",
X"55558355",
X"73802e97",
X"387651ee",
X"f83f83e0",
X"80088817",
X"0c7551ef",
X"a93f83e0",
X"80085574",
X"83e0800c",
X"933d0d04",
X"e43d0d6e",
X"a13d0840",
X"5e855683",
X"e0980880",
X"2e848538",
X"9e3df405",
X"841f0c7e",
X"98387d51",
X"eef83f83",
X"e0800856",
X"83ee3981",
X"4181f639",
X"834181f1",
X"39933d7f",
X"96054159",
X"807f8295",
X"055e5675",
X"6081ff05",
X"34834190",
X"1e08762e",
X"81d338a0",
X"547d2270",
X"852b83e0",
X"06545890",
X"1e085278",
X"519adc3f",
X"83e08008",
X"4183e080",
X"08ffb838",
X"78335c7b",
X"802effb4",
X"388b1933",
X"70bf0671",
X"81065243",
X"5574802e",
X"80de387b",
X"81bf0655",
X"748f2480",
X"d3389a19",
X"33557480",
X"cb38f31d",
X"70585d81",
X"56758b2e",
X"09810685",
X"388e568b",
X"39759a2e",
X"09810683",
X"389c5675",
X"19707081",
X"05523371",
X"33811a82",
X"1a5f5b52",
X"5b557486",
X"38797734",
X"853980df",
X"7734777b",
X"57577aa0",
X"2e098106",
X"c0388156",
X"7b81e532",
X"7030709f",
X"2a515155",
X"7bae2e93",
X"3874802e",
X"8e386183",
X"2a708106",
X"51557480",
X"2e97387d",
X"51ede23f",
X"83e08008",
X"4183e080",
X"08873890",
X"1e08feaf",
X"38806034",
X"75802e88",
X"387c527f",
X"5183a53f",
X"60802e86",
X"38800b90",
X"1f0c6056",
X"60832e85",
X"386081d0",
X"38891f57",
X"901e0880",
X"2e81a838",
X"80567519",
X"70335155",
X"74a02ea0",
X"3874852e",
X"09810684",
X"3881e555",
X"74777081",
X"05593481",
X"167081ff",
X"06575587",
X"7627d738",
X"88193355",
X"74a02ea9",
X"38ae7770",
X"81055934",
X"88567519",
X"70335155",
X"74a02e95",
X"38747770",
X"81055934",
X"81167081",
X"ff065755",
X"8a7627e2",
X"388b1933",
X"7f880534",
X"9f19339e",
X"1a337198",
X"2b71902b",
X"079d1c33",
X"70882b72",
X"079c1e33",
X"7107640c",
X"52991d33",
X"981e3371",
X"882b0753",
X"51535759",
X"56747f84",
X"05239719",
X"33961a33",
X"71882b07",
X"5656747f",
X"86052380",
X"77347d51",
X"ebf33f83",
X"e0800883",
X"32703070",
X"72079f2c",
X"83e08008",
X"06525656",
X"961f3355",
X"748a3889",
X"1f52961f",
X"5181b13f",
X"7583e080",
X"0c9e3d0d",
X"04fd3d0d",
X"75775354",
X"73335170",
X"89387133",
X"5170802e",
X"a1387333",
X"72335253",
X"72712785",
X"38ff5194",
X"39707327",
X"85388151",
X"8b398114",
X"81135354",
X"d3398051",
X"7083e080",
X"0c853d0d",
X"04fd3d0d",
X"75775454",
X"72337081",
X"ff065252",
X"70802ea3",
X"387181ff",
X"068114ff",
X"bf125354",
X"52709926",
X"8938a012",
X"7081ff06",
X"53517174",
X"70810556",
X"34d23980",
X"7434853d",
X"0d04ffbd",
X"3d0d80c6",
X"3d0852a5",
X"3d705254",
X"ffb33f80",
X"c73d0852",
X"853d7052",
X"53ffa63f",
X"72527351",
X"fedf3f80",
X"c53d0d04",
X"fe3d0d74",
X"76535371",
X"70810553",
X"33517073",
X"70810555",
X"3470f038",
X"843d0d04",
X"fe3d0d74",
X"52807233",
X"52537073",
X"2e8d3881",
X"12811471",
X"33535452",
X"70f53872",
X"83e0800c",
X"843d0d04",
X"7183e38c",
X"0c888080",
X"0b83e388",
X"0c848080",
X"0b83e390",
X"0c04f03d",
X"0d838080",
X"5683e38c",
X"081683e3",
X"88081756",
X"54743374",
X"3483e390",
X"08165480",
X"74348116",
X"56758380",
X"a02e0981",
X"06db3883",
X"d0805683",
X"e38c0816",
X"83e38808",
X"17565474",
X"33743483",
X"e3900816",
X"54807434",
X"81165675",
X"83d0a02e",
X"098106db",
X"3883a880",
X"5683e38c",
X"081683e3",
X"88081756",
X"54743374",
X"3483e390",
X"08165480",
X"74348116",
X"567583a8",
X"902e0981",
X"06db3880",
X"5683e38c",
X"081683e3",
X"90081755",
X"55733375",
X"34811656",
X"75818080",
X"2e098106",
X"e43886d0",
X"3f893d58",
X"a25380dd",
X"f0527751",
X"9cab3f80",
X"578c8056",
X"83e39008",
X"16771955",
X"55733375",
X"34811681",
X"18585676",
X"a22e0981",
X"06e63880",
X"e0940854",
X"86743480",
X"e0980854",
X"80743480",
X"e0c80854",
X"80743480",
X"e0b80854",
X"af743480",
X"e0c40854",
X"bf743480",
X"e0c00854",
X"80743480",
X"e0bc0854",
X"9f743480",
X"e0b40854",
X"80743480",
X"e0a40854",
X"f8743480",
X"e09c0854",
X"76743480",
X"e08c0854",
X"82743480",
X"e0a00854",
X"82743492",
X"3d0d04fe",
X"3d0d8053",
X"83e39008",
X"1383e38c",
X"08145252",
X"70337234",
X"81135372",
X"8180802e",
X"098106e4",
X"38838080",
X"5383e390",
X"081383e3",
X"8c081452",
X"52703372",
X"34811353",
X"728380a0",
X"2e098106",
X"e43883d0",
X"805383e3",
X"90081383",
X"e38c0814",
X"52527033",
X"72348113",
X"537283d0",
X"a02e0981",
X"06e43883",
X"a8805383",
X"e3900813",
X"83e38c08",
X"14525270",
X"33723481",
X"13537283",
X"a8902e09",
X"8106e438",
X"843d0d04",
X"803d0d80",
X"e1a40870",
X"08810683",
X"e0800c51",
X"823d0d04",
X"ff3d0d80",
X"e1a40870",
X"0870fe06",
X"7607720c",
X"5252833d",
X"0d04803d",
X"0d80e1a4",
X"08700870",
X"812c8106",
X"83e0800c",
X"5151823d",
X"0d04ff3d",
X"0d80e1a4",
X"08700870",
X"fd067610",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80e1a408",
X"70087082",
X"2cbf0683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80e1a408",
X"700870fe",
X"83067682",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d80e1a4",
X"08700870",
X"882c8706",
X"83e0800c",
X"5151823d",
X"0d04ff3d",
X"0d80e1a4",
X"08700870",
X"f1ff0676",
X"882b0772",
X"0c525283",
X"3d0d0480",
X"3d0d80e1",
X"a4087008",
X"708b2cbf",
X"0683e080",
X"0c515182",
X"3d0d04ff",
X"3d0d80e1",
X"a4087008",
X"70f88fff",
X"06768b2b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80e1b408",
X"70087088",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04803d0d",
X"80e1b408",
X"70087089",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04803d0d",
X"80e1b408",
X"7008708a",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04803d0d",
X"80e1b408",
X"7008708b",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04fd3d0d",
X"7581e629",
X"872a80e1",
X"94085473",
X"0c853d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727081",
X"055434ff",
X"1151f039",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708405",
X"540cff11",
X"51f03984",
X"3d0d04fe",
X"3d0d8180",
X"80538052",
X"88800a51",
X"ffb33fa0",
X"80538052",
X"82800a51",
X"c73f843d",
X"0d04803d",
X"0d8151fc",
X"cf3f7280",
X"2e8338d3",
X"3f8151fc",
X"f13f8051",
X"fcec3f80",
X"51fcb93f",
X"823d0d04",
X"fd3d0d75",
X"52805480",
X"ff722588",
X"38810bff",
X"80135354",
X"ffbf1251",
X"70992686",
X"38e01252",
X"9e39ff9f",
X"12519971",
X"279538d0",
X"12e01370",
X"54545189",
X"71278838",
X"8f732783",
X"38805273",
X"802e8538",
X"81801252",
X"7181ff06",
X"83e0800c",
X"853d0d04",
X"803d0d84",
X"d8c05180",
X"71708105",
X"53347084",
X"e0c02e09",
X"8106f038",
X"823d0d04",
X"fe3d0d02",
X"97053351",
X"ff863f83",
X"e0800881",
X"ff0683e3",
X"98085452",
X"8073249b",
X"3883e3b4",
X"08137283",
X"e3b80807",
X"53537173",
X"3483e398",
X"08810583",
X"e3980c84",
X"3d0d04fa",
X"3d0d8280",
X"0a1b5580",
X"57883dfc",
X"05547953",
X"74527851",
X"d6933f88",
X"3d0d04fe",
X"3d0d83e3",
X"ac085274",
X"51dcf03f",
X"83e08008",
X"8c387653",
X"755283e3",
X"ac0851c7",
X"3f843d0d",
X"04fe3d0d",
X"83e3ac08",
X"53755274",
X"51d7b03f",
X"83e08008",
X"8d387753",
X"765283e3",
X"ac0851ff",
X"a23f843d",
X"0d04fd3d",
X"0d83e3b0",
X"0851d6a4",
X"3f83e080",
X"0890802e",
X"098106ad",
X"38805483",
X"c1808053",
X"83e08008",
X"5283e3b0",
X"0851fef3",
X"3f87c180",
X"80143387",
X"c1908015",
X"34811454",
X"7390802e",
X"098106e9",
X"38853d0d",
X"0480def8",
X"0b83e080",
X"0c04f73d",
X"0d805a80",
X"59805880",
X"705757fd",
X"e73f800b",
X"83e3980c",
X"800b83e3",
X"b80c80de",
X"fc51d18f",
X"3f81800b",
X"83e3b80c",
X"80df8051",
X"d1813f80",
X"d00b83e3",
X"980c7530",
X"70770780",
X"2570872b",
X"83e3b80c",
X"5154f9d1",
X"3f83e080",
X"085280df",
X"8851d0db",
X"3f80f80b",
X"83e3980c",
X"75813270",
X"30707207",
X"80257087",
X"2b83e3b8",
X"0c515555",
X"ff833f83",
X"e0800852",
X"80df9451",
X"d0b13f81",
X"a00b83e3",
X"980c7582",
X"32703070",
X"72078025",
X"70872b83",
X"e3b80c51",
X"5583e3b0",
X"085255d1",
X"cb3f83e0",
X"80085280",
X"df9c51d0",
X"823f81c8",
X"0b83e398",
X"0c758332",
X"70307072",
X"07802570",
X"872b83e3",
X"b80c5155",
X"80dfa452",
X"55cfe03f",
X"81f00b83",
X"e3980c75",
X"84327030",
X"70720780",
X"2570872b",
X"83e3b80c",
X"515580df",
X"b45255cf",
X"be3f8298",
X"0b83e398",
X"0c758532",
X"70307072",
X"07802570",
X"872b83e3",
X"b80c5155",
X"80dfcc52",
X"55cf9c3f",
X"82c00b83",
X"e3980c75",
X"86327030",
X"70720780",
X"2570872b",
X"83e3b80c",
X"515580df",
X"e45255ce",
X"fa3f868d",
X"a051f9d1",
X"3f805288",
X"3d705254",
X"87b03f83",
X"52735187",
X"a93f7816",
X"56758025",
X"85388056",
X"90398676",
X"25853886",
X"56873975",
X"862682cb",
X"38758429",
X"80de9405",
X"54730804",
X"f7a33f83",
X"e0800878",
X"56547481",
X"2e098106",
X"893883e0",
X"80081054",
X"903974ff",
X"2e098106",
X"883883e0",
X"8008812c",
X"54907425",
X"85389054",
X"88397380",
X"24833881",
X"547351f7",
X"803f81ff",
X"39f7933f",
X"83e08008",
X"18547380",
X"25853880",
X"54883987",
X"74258338",
X"87547351",
X"f7903f81",
X"de397787",
X"3879802e",
X"81d5388a",
X"dd0b83e0",
X"9c0c83e3",
X"b00851ff",
X"bfed3ffb",
X"bd3f81bf",
X"3979802e",
X"81b9388b",
X"900b83e0",
X"9c0c83e3",
X"ac0851ff",
X"bfd13f75",
X"832e0981",
X"06943881",
X"80805382",
X"80805283",
X"e3ac0851",
X"faa93f81",
X"87397584",
X"2e098106",
X"af388280",
X"80538180",
X"805283e3",
X"ac0851fa",
X"8e3f8054",
X"84828080",
X"14338481",
X"80801534",
X"81145473",
X"8180802e",
X"098106e8",
X"3880d139",
X"75852e09",
X"810680c8",
X"38805481",
X"80805380",
X"c0805283",
X"e3ac0851",
X"f9d53f82",
X"80805380",
X"c0805283",
X"e3ac0851",
X"f9c53f84",
X"81808014",
X"338481c0",
X"80153484",
X"82808014",
X"338482c0",
X"80153481",
X"14547380",
X"c0802e09",
X"8106dc38",
X"81548c39",
X"79873876",
X"802efad3",
X"38805473",
X"83e0800c",
X"8b3d0d04",
X"ff3d0df5",
X"e43f83e0",
X"8008802e",
X"86388051",
X"80dd39f5",
X"ec3f83e0",
X"800880d1",
X"38f6923f",
X"83e08008",
X"802eaa38",
X"8151f3e4",
X"3ff08f3f",
X"800b83e3",
X"980cfa82",
X"3f83e080",
X"0852ff0b",
X"83e3980c",
X"f2ad3f71",
X"a4387151",
X"f3c23fa2",
X"39f5c63f",
X"83e08008",
X"802e9738",
X"8151f3b0",
X"3fefdb3f",
X"ff0b83e3",
X"980cf287",
X"3f8151f6",
X"c93f833d",
X"0d04fc3d",
X"0d908080",
X"52868480",
X"8051d0bd",
X"3f83e080",
X"08b83880",
X"e1b851d5",
X"803f83e0",
X"800883e3",
X"b0085480",
X"dff05383",
X"e0800852",
X"55cfdc3f",
X"83e08008",
X"8438f8ba",
X"3f818080",
X"54828080",
X"5380dfec",
X"527451f8",
X"843f8151",
X"f5f43ffe",
X"b73ffc39",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"0283e08c",
X"08fc050c",
X"800b83e3",
X"9c0b83e0",
X"8c08f805",
X"0c83e08c",
X"08f4050c",
X"cec33f83",
X"e0800886",
X"05fc0683",
X"e08c08f0",
X"050c0283",
X"e08c08f0",
X"0508310d",
X"833d7083",
X"e08c08f8",
X"05087084",
X"0583e08c",
X"08f8050c",
X"0c51cb92",
X"3f83e08c",
X"08f40508",
X"810583e0",
X"8c08f405",
X"0c83e08c",
X"08f40508",
X"862e0981",
X"06ffad38",
X"86948080",
X"51edd93f",
X"ff0b83e3",
X"980c800b",
X"83e3b80c",
X"84d8c00b",
X"83e3b40c",
X"8151f1a8",
X"3f8151f1",
X"d13f8051",
X"f1cc3f81",
X"51f1f63f",
X"8151f2d3",
X"3f8251f2",
X"9d3f80c5",
X"f8528051",
X"c8d63ffd",
X"e93f83e0",
X"8c08fc05",
X"080d800b",
X"83e0800c",
X"873d0d83",
X"e08c0c04",
X"fd3d0d75",
X"5480740c",
X"800b8415",
X"0c800b88",
X"150c80e0",
X"88087033",
X"80e08c08",
X"70337082",
X"2a708106",
X"70307072",
X"07700970",
X"9f2c7806",
X"9e065451",
X"51545151",
X"55525451",
X"80729806",
X"52537088",
X"2e098106",
X"83388153",
X"70983270",
X"30708025",
X"75713184",
X"180c5151",
X"51807286",
X"06525370",
X"822e0981",
X"06833881",
X"53708632",
X"70307080",
X"25757131",
X"770c5151",
X"51719432",
X"70307080",
X"2588170c",
X"5151853d",
X"0d04fe3d",
X"0d747654",
X"527151fe",
X"e73f7281",
X"2ea23881",
X"73268d38",
X"72822eab",
X"3872832e",
X"9f38e639",
X"7108e238",
X"841208dd",
X"38881208",
X"d838a039",
X"88120881",
X"2e098106",
X"cc389439",
X"88120881",
X"2e8d3871",
X"08893884",
X"1208802e",
X"ffb73884",
X"3d0d04fd",
X"3d0d7554",
X"7383e3c0",
X"082ea738",
X"80e19808",
X"74a00a07",
X"710c80e1",
X"a8085353",
X"71085170",
X"802ef938",
X"80730c71",
X"085170fb",
X"387383e3",
X"c00c853d",
X"0d04ff0b",
X"83e3c00c",
X"8180800b",
X"83e3bc0c",
X"800b83e0",
X"800c04fc",
X"3d0d7602",
X"8405a205",
X"22028805",
X"a605227a",
X"54555555",
X"ff9d3f72",
X"802ea338",
X"83e3bc08",
X"14527133",
X"75708105",
X"57348114",
X"7083ffff",
X"06ff1570",
X"83ffff06",
X"56525552",
X"da39800b",
X"83e0800c",
X"863d0d04",
X"f73d0d7b",
X"7d7f1158",
X"55598055",
X"73762eb1",
X"3883e3bc",
X"088b3d59",
X"57741970",
X"3375fc06",
X"1970085d",
X"7683067b",
X"07535454",
X"51727134",
X"79720c81",
X"14811656",
X"5473762e",
X"098106d9",
X"38800b83",
X"e0800c8b",
X"3d0d04fe",
X"3d0d80e1",
X"980883e3",
X"c008900a",
X"07710c80",
X"e1a80853",
X"53710851",
X"70802ef9",
X"3880730c",
X"71085170",
X"fb38843d",
X"0d0483e0",
X"8c080283",
X"e08c0cfd",
X"3d0d8053",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"83d43f83",
X"e0800870",
X"83e0800c",
X"54853d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cfd3d",
X"0d815383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"05085183",
X"a13f83e0",
X"80087083",
X"e0800c54",
X"853d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cf93d0d",
X"800b83e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"8025b938",
X"83e08c08",
X"88050830",
X"83e08c08",
X"88050c80",
X"0b83e08c",
X"08f4050c",
X"83e08c08",
X"fc05088a",
X"38810b83",
X"e08c08f4",
X"050c83e0",
X"8c08f405",
X"0883e08c",
X"08fc050c",
X"83e08c08",
X"8c050880",
X"25b93883",
X"e08c088c",
X"05083083",
X"e08c088c",
X"050c800b",
X"83e08c08",
X"f0050c83",
X"e08c08fc",
X"05088a38",
X"810b83e0",
X"8c08f005",
X"0c83e08c",
X"08f00508",
X"83e08c08",
X"fc050c80",
X"5383e08c",
X"088c0508",
X"5283e08c",
X"08880508",
X"5181df3f",
X"83e08008",
X"7083e08c",
X"08f8050c",
X"5483e08c",
X"08fc0508",
X"802e9038",
X"83e08c08",
X"f8050830",
X"83e08c08",
X"f8050c83",
X"e08c08f8",
X"05087083",
X"e0800c54",
X"893d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"800b83e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"80259938",
X"83e08c08",
X"88050830",
X"83e08c08",
X"88050c81",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"8c050880",
X"25903883",
X"e08c088c",
X"05083083",
X"e08c088c",
X"050c8153",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"bd3f83e0",
X"80087083",
X"e08c08f8",
X"050c5483",
X"e08c08fc",
X"0508802e",
X"903883e0",
X"8c08f805",
X"083083e0",
X"8c08f805",
X"0c83e08c",
X"08f80508",
X"7083e080",
X"0c54873d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cfd",
X"3d0d810b",
X"83e08c08",
X"fc050c80",
X"0b83e08c",
X"08f8050c",
X"83e08c08",
X"8c050883",
X"e08c0888",
X"050827b9",
X"3883e08c",
X"08fc0508",
X"802eae38",
X"800b83e0",
X"8c088c05",
X"0824a238",
X"83e08c08",
X"8c050810",
X"83e08c08",
X"8c050c83",
X"e08c08fc",
X"05081083",
X"e08c08fc",
X"050cffb8",
X"3983e08c",
X"08fc0508",
X"802e80e1",
X"3883e08c",
X"088c0508",
X"83e08c08",
X"88050826",
X"ad3883e0",
X"8c088805",
X"0883e08c",
X"088c0508",
X"3183e08c",
X"0888050c",
X"83e08c08",
X"f8050883",
X"e08c08fc",
X"05080783",
X"e08c08f8",
X"050c83e0",
X"8c08fc05",
X"08812a83",
X"e08c08fc",
X"050c83e0",
X"8c088c05",
X"08812a83",
X"e08c088c",
X"050cff95",
X"3983e08c",
X"08900508",
X"802e9338",
X"83e08c08",
X"88050870",
X"83e08c08",
X"f4050c51",
X"913983e0",
X"8c08f805",
X"087083e0",
X"8c08f405",
X"0c5183e0",
X"8c08f405",
X"0883e080",
X"0c853d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cff3d",
X"0d800b83",
X"e08c08fc",
X"050c83e0",
X"8c088805",
X"088106ff",
X"11700970",
X"83e08c08",
X"8c050806",
X"83e08c08",
X"fc050811",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"0508812a",
X"83e08c08",
X"88050c83",
X"e08c088c",
X"05081083",
X"e08c088c",
X"050c5151",
X"515183e0",
X"8c088805",
X"08802e84",
X"38ffab39",
X"83e08c08",
X"fc050870",
X"83e0800c",
X"51833d0d",
X"83e08c0c",
X"04fc3d0d",
X"7670797b",
X"55555555",
X"8f72278c",
X"38727507",
X"83065170",
X"802ea938",
X"ff125271",
X"ff2e9838",
X"72708105",
X"54337470",
X"81055634",
X"ff125271",
X"ff2e0981",
X"06ea3874",
X"83e0800c",
X"863d0d04",
X"74517270",
X"84055408",
X"71708405",
X"530c7270",
X"84055408",
X"71708405",
X"530c7270",
X"84055408",
X"71708405",
X"530c7270",
X"84055408",
X"71708405",
X"530cf012",
X"52718f26",
X"c9388372",
X"27953872",
X"70840554",
X"08717084",
X"05530cfc",
X"12527183",
X"26ed3870",
X"54ff8139",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"0000255c",
X"0000259d",
X"000025be",
X"000025dd",
X"000025dd",
X"000025dd",
X"00002698",
X"25732025",
X"73000000",
X"20000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"524f4d00",
X"42494e00",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"31364b00",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"43617274",
X"72696467",
X"65203332",
X"6b000000",
X"43617274",
X"72696467",
X"65203136",
X"6b206f6e",
X"65206368",
X"69700000",
X"43617274",
X"72696467",
X"65203136",
X"6b207477",
X"6f206368",
X"69700000",
X"45786974",
X"00000000",
X"61636964",
X"35323030",
X"2e726f6d",
X"00000000",
X"00000000",
X"00000000",
X"0001e80a",
X"0001e809",
X"0001e80f",
X"0001d40e",
X"0001d403",
X"0001d402",
X"0001d400",
X"0001d401",
X"0001d409",
X"0001d301",
X"0001d300",
X"0001c010",
X"0001c01b",
X"0001c016",
X"0001c019",
X"0001c018",
X"0001c017",
X"0001c01a",
X"0004007c",
X"00040078",
X"00040074",
X"00040068",
X"00040060",
X"0004005c",
X"00040058",
X"00040054",
X"00040050",
X"0004004c",
X"00040048",
X"00040044",
X"00040040",
X"00040034",
X"00040030",
X"0004002c",
X"00040028",
X"00040024",
X"00040020",
X"0004001c",
X"00040018",
X"00040014",
X"00040010",
X"0004000c",
X"00040008",
X"00040004",
X"00040000",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
