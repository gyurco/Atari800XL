
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81d3",
X"a8738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81da",
X"bc0c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757580f1",
X"922d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7580f0d1",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80dbdd04",
X"fd3d0d75",
X"705254ae",
X"a63f83c0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"c0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83c0",
X"8008732e",
X"a13883c0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183c0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83c2d008",
X"248a38b4",
X"f73fff0b",
X"83c2d00c",
X"800b83c0",
X"800c04ff",
X"3d0d7352",
X"83c0ac08",
X"722e8d38",
X"d93f7151",
X"96993f71",
X"83c0ac0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"558154bc",
X"15088191",
X"387451cf",
X"3f795880",
X"7a2580f7",
X"3883c380",
X"0870892a",
X"5783ff06",
X"78848072",
X"31565657",
X"73782583",
X"38735575",
X"83c2d008",
X"2e8438ff",
X"893f83c2",
X"d0088025",
X"a6387589",
X"2b5198dc",
X"3f83c380",
X"088f3dfc",
X"11555c54",
X"8152f81b",
X"5196c63f",
X"761483c3",
X"800c7583",
X"c2d00c74",
X"53765278",
X"51b3a83f",
X"83c08008",
X"83c38008",
X"1683c380",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8b3861",
X"7a710c54",
X"75547580",
X"2e833881",
X"547383c0",
X"800c8e3d",
X"0d04fc3d",
X"0dfe9b3f",
X"7651feaf",
X"3f863dfc",
X"05537852",
X"775195e9",
X"3f797571",
X"0c5483c0",
X"80085483",
X"c0800880",
X"2e833881",
X"547383c0",
X"800c863d",
X"0d04fe3d",
X"0d7583c2",
X"d0085353",
X"80722489",
X"3871732e",
X"8438fdd6",
X"3f7451fd",
X"ea3f7251",
X"97ae3f83",
X"c0800852",
X"83c08008",
X"802e8338",
X"81527183",
X"c0800c84",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"c0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"c0800c51",
X"823d0d04",
X"80c40b83",
X"c0800c04",
X"fd3d0d75",
X"77715470",
X"535553a9",
X"fe3f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfceb3f",
X"735193ab",
X"3f7383c0",
X"ac0c83c0",
X"80085383",
X"c0800880",
X"2e833881",
X"537283c0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcbf3f",
X"72802ea5",
X"38bc1308",
X"527351a9",
X"883f83c0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"c0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83c0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83c2d0",
X"0c7483c0",
X"b00c7583",
X"c2cc0caf",
X"dc3f83c0",
X"800881ff",
X"06528153",
X"71993883",
X"c2e8518e",
X"943f83c0",
X"80085283",
X"c0800880",
X"2e833872",
X"52715372",
X"83c0800c",
X"843d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"51a6f93f",
X"83c08008",
X"557483c0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"c0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283c2cc",
X"085180df",
X"d43f83c0",
X"800857f9",
X"e13f7952",
X"83c2d451",
X"95b73f83",
X"c0800854",
X"805383c0",
X"8008732e",
X"09810682",
X"833883c0",
X"b0080b0b",
X"81d8b053",
X"705256a6",
X"b63f0b0b",
X"81d8b052",
X"80c01651",
X"a6a93f75",
X"bc170c73",
X"82c0170c",
X"810b82c4",
X"170c810b",
X"82c8170c",
X"7382cc17",
X"0cff1782",
X"d0175557",
X"81913983",
X"c0bc3370",
X"822a7081",
X"06515455",
X"72818038",
X"74812a81",
X"06587780",
X"f6387484",
X"2a810682",
X"c4150c83",
X"c0bc3381",
X"0682c815",
X"0c795273",
X"51a5d03f",
X"7351a5e7",
X"3f83c080",
X"081453af",
X"73708105",
X"553472bc",
X"150c83c0",
X"bd527251",
X"a5b13f83",
X"c0b40882",
X"c0150c83",
X"c0ca5280",
X"c01451a5",
X"9e3f7880",
X"2e8d3873",
X"51782d83",
X"c0800880",
X"2e993877",
X"82cc150c",
X"75802e86",
X"387382cc",
X"170c7382",
X"d015ff19",
X"59555676",
X"802e9b38",
X"83c0b452",
X"83c2d451",
X"94ad3f83",
X"c080088a",
X"3883c0bd",
X"335372fe",
X"d2387880",
X"2e893883",
X"c0b00851",
X"fcb83f83",
X"c0b00853",
X"7283c080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb53f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f690",
X"3f83c080",
X"08745387",
X"3d705355",
X"55f6b03f",
X"f7903f73",
X"51d33f63",
X"53745283",
X"c0800851",
X"fab83f92",
X"3d0d0471",
X"83c0800c",
X"0480c012",
X"83c0800c",
X"04803d0d",
X"7282c011",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"c0800c51",
X"823d0d04",
X"f93d0d79",
X"83c09008",
X"57578177",
X"27819638",
X"76881708",
X"27818e38",
X"75335574",
X"822e8938",
X"74832eb3",
X"3880fe39",
X"74547610",
X"83fe0653",
X"76882a8c",
X"17080552",
X"893dfc05",
X"51aa8a3f",
X"83c08008",
X"80df3802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d13984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"51a9da3f",
X"83c08008",
X"b038029f",
X"05330284",
X"059e0533",
X"71982b71",
X"902b0702",
X"8c059d05",
X"3370882b",
X"72078d3d",
X"337180ff",
X"fffe8006",
X"07515253",
X"57585683",
X"39815574",
X"83c0800c",
X"893d0d04",
X"fb3d0d83",
X"c09008fe",
X"19881208",
X"fe055556",
X"54805674",
X"73278d38",
X"82143375",
X"71299416",
X"08055753",
X"7583c080",
X"0c873d0d",
X"04fc3d0d",
X"7652800b",
X"83c09008",
X"70335152",
X"5370832e",
X"09810691",
X"38951233",
X"94133371",
X"982b7190",
X"2b075555",
X"519b1233",
X"9a133371",
X"882b0774",
X"0783c080",
X"0c55863d",
X"0d04fc3d",
X"0d7683c0",
X"90085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"fed63f83",
X"c0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183c080",
X"0c863d0d",
X"04fa3d0d",
X"7883c090",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fcb13f",
X"81527183",
X"c0800827",
X"a8388352",
X"83c08008",
X"88170827",
X"9c3883c0",
X"80088c16",
X"0c83c080",
X"0851fdbc",
X"3f83c080",
X"0890160c",
X"73752380",
X"527183c0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585e5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"9f269138",
X"7a51fdd2",
X"3f83c080",
X"0856807d",
X"34838139",
X"933d841c",
X"08705859",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"3880705a",
X"5c887f08",
X"5f5a7b81",
X"1d7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535e57",
X"557480e7",
X"3876ae2e",
X"09810683",
X"38815578",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675bb",
X"3888598b",
X"5affab39",
X"76982b55",
X"74802587",
X"3881d2b8",
X"173357ff",
X"9f175574",
X"99268938",
X"e0177081",
X"ff065855",
X"78811a70",
X"81ff0672",
X"1b535b57",
X"55767534",
X"fef8397b",
X"1e7f0c80",
X"5576a026",
X"83388155",
X"748b1934",
X"7a51fc82",
X"3f83c080",
X"0880f538",
X"a0547a22",
X"70852b83",
X"e0065455",
X"901b0852",
X"7c51a495",
X"3f83c080",
X"085783c0",
X"80088181",
X"387c3355",
X"74802e80",
X"f4388b1d",
X"3370832a",
X"70810651",
X"565674b4",
X"388b7d84",
X"1d0883c0",
X"8008595b",
X"5b58ff18",
X"5877ff2e",
X"9a387970",
X"81055b33",
X"79708105",
X"5b337171",
X"31525656",
X"75802ee2",
X"38863975",
X"802e9638",
X"7a51fbe5",
X"3fff8639",
X"83c08008",
X"5683c080",
X"08b63883",
X"39765684",
X"1b088b11",
X"33515574",
X"a7388b1d",
X"3370842a",
X"70810651",
X"56567489",
X"38835694",
X"39815690",
X"397c51fa",
X"943f83c0",
X"8008881c",
X"0cfd8139",
X"7583c080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"51a2da3f",
X"835683c0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"51a2ae3f",
X"83c08008",
X"98388117",
X"33773371",
X"882b0783",
X"c0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"7651a285",
X"3f83c080",
X"08983881",
X"17337733",
X"71882b07",
X"83c08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583c080",
X"0c8a3d0d",
X"04eb3d0d",
X"675a800b",
X"83c0900c",
X"a1a73f83",
X"c0800881",
X"06558256",
X"7483ef38",
X"7475538f",
X"3d705357",
X"59feca3f",
X"83c08008",
X"81ff0657",
X"76812e09",
X"810680d4",
X"38905483",
X"be537452",
X"7551a199",
X"3f83c080",
X"0880c938",
X"8f3d3355",
X"74802e80",
X"c93802bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"33710770",
X"587b575e",
X"525e5759",
X"57fdee3f",
X"83c08008",
X"81ff0657",
X"76832e09",
X"81068638",
X"815682f2",
X"3976802e",
X"86388656",
X"82e839a4",
X"548d5378",
X"527551a0",
X"b03f8156",
X"83c08008",
X"82d43802",
X"be053302",
X"8405bd05",
X"3371882b",
X"07595d77",
X"ab380280",
X"ce053302",
X"840580cd",
X"05337198",
X"2b71902b",
X"07973d33",
X"70882b72",
X"07029405",
X"80cb0533",
X"71075452",
X"5e575956",
X"02b70533",
X"78712902",
X"8805b605",
X"33028c05",
X"b5053371",
X"882b0770",
X"1d707f8c",
X"050c5f59",
X"57595d8e",
X"3d33821b",
X"3402b905",
X"33903d33",
X"71882b07",
X"5a5c7884",
X"1b2302bb",
X"05330284",
X"05ba0533",
X"71882b07",
X"565c74ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"07515253",
X"575e5c74",
X"76317831",
X"79842a90",
X"3d335471",
X"71315356",
X"5680d0b9",
X"3f83c080",
X"08820570",
X"881c0c83",
X"c08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83c0900c",
X"80567583",
X"c0800c97",
X"3d0d04e9",
X"3d0d83c0",
X"90085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e53f83c0",
X"80085483",
X"c0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f489",
X"3f83c080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383c080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83c09008",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0e93f",
X"83c08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"833f83c0",
X"80085583",
X"c0800880",
X"2eff8938",
X"83c08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"519ad63f",
X"83c08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83c0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83c09008",
X"55568555",
X"73802e81",
X"e3388114",
X"33810653",
X"84557280",
X"2e81d538",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b9388214",
X"3370892b",
X"56537680",
X"2eb73874",
X"52ff1651",
X"80cbba3f",
X"83c08008",
X"ff187654",
X"70535853",
X"80cbaa3f",
X"83c08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed63f83",
X"c0800853",
X"810b83c0",
X"8008278b",
X"38881408",
X"83c08008",
X"26883880",
X"0b811534",
X"b03983c0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc53f",
X"83c08008",
X"8c3883c0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683c0",
X"800805a8",
X"150c8055",
X"7483c080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83c09008",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1cf3f",
X"83c08008",
X"5583c080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef5",
X"3f83c080",
X"0888170c",
X"7551efa6",
X"3f83c080",
X"08557483",
X"c0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683c0",
X"9008802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f53f83c0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"96df3f83",
X"c0800841",
X"83c08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"eddf3f83",
X"c0800841",
X"83c08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"8e853f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f03f83c0",
X"80088332",
X"70307072",
X"079f2c83",
X"c0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"8c913f75",
X"83c0800c",
X"9e3d0d04",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"7751e0d2",
X"3f83c080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3381dac4",
X"0b81dac4",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"527751e0",
X"813f83c0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583c0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"558b983f",
X"83c08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"8114518a",
X"b03f83c0",
X"80083070",
X"83c08008",
X"07802583",
X"c0800c53",
X"863d0d04",
X"fc3d0d76",
X"705255e6",
X"ee3f83c0",
X"80085481",
X"5383c080",
X"0880c138",
X"7451e6b1",
X"3f83c080",
X"0881d8c0",
X"5383c080",
X"085253ff",
X"913f83c0",
X"8008a138",
X"81d8c452",
X"7251ff82",
X"3f83c080",
X"08923881",
X"d8c85272",
X"51fef33f",
X"83c08008",
X"802e8338",
X"81547353",
X"7283c080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"e68d3f81",
X"5383c080",
X"08983873",
X"51e5d63f",
X"83c39808",
X"5283c080",
X"0851feba",
X"3f83c080",
X"08537283",
X"c0800c85",
X"3d0d04df",
X"3d0da43d",
X"0870525e",
X"dbfb3f83",
X"c0800833",
X"953d5654",
X"73963881",
X"ddd45274",
X"5189903f",
X"9a397d52",
X"7851defc",
X"3f84cf39",
X"7d51dbe1",
X"3f83c080",
X"08527451",
X"db913f80",
X"43804280",
X"41804083",
X"c3a00852",
X"943d7052",
X"5de1e43f",
X"83c08008",
X"59800b83",
X"c0800855",
X"5b83c080",
X"087b2e94",
X"38811b74",
X"525be4e6",
X"3f83c080",
X"085483c0",
X"8008ee38",
X"805aff5f",
X"7909709f",
X"2c7b065b",
X"547a7a24",
X"8438ff1b",
X"5af61a70",
X"09709f2c",
X"72067bff",
X"125a5a52",
X"55558075",
X"25953876",
X"51e4ab3f",
X"83c08008",
X"76ff1858",
X"55577380",
X"24ed3874",
X"7f2e8638",
X"a0d83f74",
X"5f78ff1b",
X"70585d58",
X"807a2595",
X"387751e4",
X"813f83c0",
X"800876ff",
X"18585558",
X"738024ed",
X"38800b83",
X"c7d00c80",
X"0b83c884",
X"0c81d8cc",
X"518d8f3f",
X"81800b83",
X"c8840c81",
X"d8d4518d",
X"813fa80b",
X"83c7d00c",
X"76802e80",
X"e43883c7",
X"d0087779",
X"32703070",
X"72078025",
X"70872b83",
X"c8840c51",
X"56785356",
X"56e3b83f",
X"83c08008",
X"802e8838",
X"81d8dc51",
X"8cc83f76",
X"51e2fa3f",
X"83c08008",
X"5281d9e8",
X"518cb73f",
X"7651e382",
X"3f83c080",
X"0883c7d0",
X"08555775",
X"74258638",
X"a81656f7",
X"397583c7",
X"d00c86f0",
X"7624ff98",
X"3887980b",
X"83c7d00c",
X"77802eb1",
X"387751e2",
X"b83f83c0",
X"80087852",
X"55e2d83f",
X"81d8e454",
X"83c08008",
X"8d388739",
X"80763481",
X"d03981d8",
X"e0547453",
X"735281d8",
X"b4518bd6",
X"3f805481",
X"d8bc518b",
X"cd3f8114",
X"5473a82e",
X"098106ef",
X"38868da0",
X"519cdd3f",
X"8052903d",
X"70525780",
X"c1943f83",
X"52765180",
X"c18c3f62",
X"818f3861",
X"802e80fb",
X"387b5473",
X"ff2e9638",
X"78802e81",
X"89387851",
X"e1dc3f83",
X"c08008ff",
X"155559e7",
X"3978802e",
X"80f43878",
X"51e1d83f",
X"83c08008",
X"802efc8e",
X"387851e1",
X"a03f83c0",
X"80085281",
X"d8b05183",
X"e33f83c0",
X"8008a338",
X"7c51859b",
X"3f83c080",
X"085574ff",
X"16565480",
X"7425ae38",
X"741d7033",
X"555673af",
X"2efecd38",
X"e9397851",
X"e0e13f83",
X"c0800852",
X"7c5184d3",
X"3f8f397f",
X"88296010",
X"057a0561",
X"055afc90",
X"3962802e",
X"fbd13880",
X"527651bf",
X"ed3fa33d",
X"0d04803d",
X"0d9088b8",
X"337081ff",
X"0670842a",
X"81327081",
X"06515151",
X"5170802e",
X"8d38a80b",
X"9088b834",
X"b80b9088",
X"b8347083",
X"c0800c82",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067085",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d3898",
X"0b9088b8",
X"34b80b90",
X"88b83470",
X"83c0800c",
X"823d0d04",
X"930b9088",
X"bc34ff0b",
X"9088a834",
X"04ff3d0d",
X"028f0533",
X"52800b90",
X"88bc348a",
X"519aa53f",
X"df3f80f8",
X"0b9088a0",
X"34800b90",
X"888834fa",
X"12527190",
X"88803480",
X"0b908898",
X"34719088",
X"90349088",
X"b8528072",
X"34b87234",
X"833d0d04",
X"803d0d02",
X"8b053351",
X"709088b4",
X"34febf3f",
X"83c08008",
X"802ef638",
X"823d0d04",
X"803d0d84",
X"39a3fe3f",
X"fed93f83",
X"c0800880",
X"2ef33890",
X"88b43370",
X"81ff0683",
X"c0800c51",
X"823d0d04",
X"803d0da3",
X"0b9088bc",
X"34ff0b90",
X"88a83490",
X"88b851a8",
X"7134b871",
X"34823d0d",
X"04803d0d",
X"9088bc33",
X"7081c006",
X"70307080",
X"2583c080",
X"0c515151",
X"823d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"832a8132",
X"70810651",
X"51515170",
X"802ee838",
X"b00b9088",
X"b834b80b",
X"9088b834",
X"823d0d04",
X"803d0d90",
X"80ac0881",
X"0683c080",
X"0c823d0d",
X"04fd3d0d",
X"75775454",
X"80732594",
X"38737081",
X"05553352",
X"81d8e851",
X"87843fff",
X"1353e939",
X"853d0d04",
X"fd3d0d75",
X"77535473",
X"33517089",
X"38713351",
X"70802ea1",
X"38733372",
X"33525372",
X"71278538",
X"ff519439",
X"70732785",
X"3881518b",
X"39811481",
X"135354d3",
X"39805170",
X"83c0800c",
X"853d0d04",
X"fd3d0d75",
X"77545472",
X"337081ff",
X"06525270",
X"802ea338",
X"7181ff06",
X"8114ffbf",
X"12535452",
X"70992689",
X"38a01270",
X"81ff0653",
X"51717470",
X"81055634",
X"d2398074",
X"34853d0d",
X"04ffbd3d",
X"0d80c63d",
X"0852a53d",
X"705254ff",
X"b33f80c7",
X"3d085285",
X"3d705253",
X"ffa63f72",
X"527351fe",
X"df3f80c5",
X"3d0d04fe",
X"3d0d7476",
X"53537170",
X"81055333",
X"51707370",
X"81055534",
X"70f03884",
X"3d0d04fe",
X"3d0d7452",
X"80723352",
X"5370732e",
X"8d388112",
X"81147133",
X"53545270",
X"f5387283",
X"c0800c84",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"b88f3f83",
X"c080087a",
X"27ee3874",
X"802e80dd",
X"38745275",
X"51b7fa3f",
X"83c08008",
X"75537652",
X"54b7fe3f",
X"83c08008",
X"7a537552",
X"56b7e23f",
X"83c08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"c08008c5",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9f",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fc813f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd53f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbb13f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83c0940c",
X"7183c098",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383c094",
X"085283c0",
X"980851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"bdba5351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fc3d",
X"0d765574",
X"83c3a808",
X"2eaf3880",
X"53745187",
X"c13f83c0",
X"800881ff",
X"06ff1470",
X"81ff0672",
X"30709f2a",
X"51525553",
X"5472802e",
X"843871dd",
X"3873fe38",
X"7483c3a8",
X"0c863d0d",
X"04ff3d0d",
X"ff0b83c3",
X"a80c84a5",
X"3f815187",
X"853f83c0",
X"800881ff",
X"065271ee",
X"3881d33f",
X"7183c080",
X"0c833d0d",
X"04fc3d0d",
X"76028405",
X"a2052202",
X"8805a605",
X"227a5455",
X"5555ff82",
X"3f72802e",
X"a03883c3",
X"bc143375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552dd",
X"39800b83",
X"c0800c86",
X"3d0d04fc",
X"3d0d7678",
X"7a115653",
X"55805371",
X"742e9338",
X"72155170",
X"3383c3bc",
X"13348112",
X"81145452",
X"ea39800b",
X"83c0800c",
X"863d0d04",
X"fd3d0d90",
X"5483c3a8",
X"085186f4",
X"3f83c080",
X"0881ff06",
X"ff157130",
X"71307073",
X"079f2a72",
X"9f2a0652",
X"55525553",
X"72db3885",
X"3d0d0480",
X"3d0d83c3",
X"b4081083",
X"c3ac0807",
X"9080a80c",
X"823d0d04",
X"800b83c3",
X"b40ce43f",
X"04810b83",
X"c3b40cdb",
X"3f04ed3f",
X"047183c3",
X"b00c0480",
X"3d0d8051",
X"f43f810b",
X"83c3b40c",
X"810b83c3",
X"ac0cffbb",
X"3f823d0d",
X"04803d0d",
X"72307074",
X"07802583",
X"c3ac0c51",
X"ffa53f82",
X"3d0d0480",
X"3d0d028b",
X"05339080",
X"a40c9080",
X"a8087081",
X"06515170",
X"f5389080",
X"a4087081",
X"ff0683c0",
X"800c5182",
X"3d0d0480",
X"3d0d81ff",
X"51d13f83",
X"c0800881",
X"ff0683c0",
X"800c823d",
X"0d04803d",
X"0d73902b",
X"73079080",
X"b40c823d",
X"0d0404fb",
X"3d0d7802",
X"84059f05",
X"3370982b",
X"55575572",
X"80259b38",
X"7580ff06",
X"56805280",
X"f751e03f",
X"83c08008",
X"81ff0654",
X"73812680",
X"ff388051",
X"fee73fff",
X"a23f8151",
X"fedf3fff",
X"9a3f7551",
X"feed3f74",
X"982a51fe",
X"e63f7490",
X"2a7081ff",
X"065253fe",
X"da3f7488",
X"2a7081ff",
X"065253fe",
X"ce3f7481",
X"ff0651fe",
X"c63f8155",
X"7580c02e",
X"09810686",
X"38819555",
X"8d397580",
X"c82e0981",
X"06843881",
X"87557451",
X"fea53f8a",
X"55fec83f",
X"83c08008",
X"81ff0670",
X"982b5454",
X"7280258c",
X"38ff1570",
X"81ff0656",
X"5374e238",
X"7383c080",
X"0c873d0d",
X"04fa3d0d",
X"fdc53f80",
X"51fdda3f",
X"8a54fe93",
X"3fff1470",
X"81ff0655",
X"5373f338",
X"73745355",
X"80c051fe",
X"a63f83c0",
X"800881ff",
X"06547381",
X"2e098106",
X"829f3883",
X"aa5280c8",
X"51fe8c3f",
X"83c08008",
X"81ff0653",
X"72812e09",
X"810681a8",
X"38745487",
X"3d741154",
X"56fdc83f",
X"83c08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e53802",
X"9a053353",
X"72812e09",
X"810681d9",
X"38029b05",
X"335380ce",
X"90547281",
X"aa2e8d38",
X"81c73980",
X"e4518acc",
X"3fff1454",
X"73802e81",
X"b838820a",
X"5281e951",
X"fda53f83",
X"c0800881",
X"ff065372",
X"de387252",
X"80fa51fd",
X"923f83c0",
X"800881ff",
X"06537281",
X"90387254",
X"731653fc",
X"d63f83c0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e8",
X"38873d33",
X"70862a70",
X"81065154",
X"548c5572",
X"80e33884",
X"5580de39",
X"745281e9",
X"51fccc3f",
X"83c08008",
X"81ff0653",
X"825581e9",
X"56817327",
X"86387355",
X"80c15680",
X"ce90548a",
X"3980e451",
X"89be3fff",
X"14547380",
X"2ea93880",
X"527551fc",
X"9a3f83c0",
X"800881ff",
X"065372e1",
X"38848052",
X"80d051fc",
X"863f83c0",
X"800881ff",
X"06537280",
X"2e833880",
X"557483c3",
X"b8348051",
X"fb873ffb",
X"c23f883d",
X"0d04fb3d",
X"0d775480",
X"0b83c3b8",
X"3370832a",
X"70810651",
X"55575572",
X"752e0981",
X"06853873",
X"892b5473",
X"5280d151",
X"fbbd3f83",
X"c0800881",
X"ff065372",
X"bd3882b8",
X"c054fb83",
X"3f83c080",
X"0881ff06",
X"537281ff",
X"2e098106",
X"8938ff14",
X"5473e738",
X"9f397281",
X"fe2e0981",
X"06963883",
X"c7bc5283",
X"c3bc51fa",
X"ed3ffad3",
X"3ffad03f",
X"83398155",
X"8051fa89",
X"3ffac43f",
X"7481ff06",
X"83c0800c",
X"873d0d04",
X"fb3d0d77",
X"83c3bc56",
X"548151f9",
X"ec3f83c3",
X"b8337083",
X"2a708106",
X"51545672",
X"85387389",
X"2b547352",
X"80d851fa",
X"b63f83c0",
X"800881ff",
X"06537280",
X"e43881ff",
X"51f9d43f",
X"81fe51f9",
X"ce3f8480",
X"53747081",
X"05563351",
X"f9c13fff",
X"137083ff",
X"ff065153",
X"72eb3872",
X"51f9b03f",
X"7251f9ab",
X"3ff9d03f",
X"83c08008",
X"9f0653a7",
X"88547285",
X"2e8c3899",
X"3980e451",
X"86f63fff",
X"1454f9b3",
X"3f83c080",
X"0881ff2e",
X"843873e9",
X"388051f8",
X"e43ff99f",
X"3f800b83",
X"c0800c87",
X"3d0d0471",
X"83c7c00c",
X"8880800b",
X"83c7bc0c",
X"8480800b",
X"83c7c40c",
X"04fd3d0d",
X"77701755",
X"7705ff1a",
X"535371ff",
X"2e943873",
X"70810555",
X"33517073",
X"70810555",
X"34ff1252",
X"e939853d",
X"0d04fc3d",
X"0d87a681",
X"55743383",
X"c7c834a0",
X"5483a080",
X"5383c7c0",
X"085283c7",
X"bc0851ff",
X"b83fa054",
X"83a48053",
X"83c7c008",
X"5283c7bc",
X"0851ffa5",
X"3f905483",
X"a8805383",
X"c7c00852",
X"83c7bc08",
X"51ff923f",
X"a0538052",
X"83c7c408",
X"83a08005",
X"5185ce3f",
X"a0538052",
X"83c7c408",
X"83a48005",
X"5185be3f",
X"90538052",
X"83c7c408",
X"83a88005",
X"5185ae3f",
X"ff753483",
X"a0805480",
X"5383c7c0",
X"085283c7",
X"c40851fe",
X"cc3f80d0",
X"805483b0",
X"805383c7",
X"c0085283",
X"c7c40851",
X"feb73f86",
X"e13fa254",
X"805383c7",
X"c4088c80",
X"055281db",
X"b851fea1",
X"3f860b87",
X"a8833480",
X"0b87a882",
X"34800b87",
X"a09a34af",
X"0b87a096",
X"34bf0b87",
X"a0973480",
X"0b87a098",
X"349f0b87",
X"a0993480",
X"0b87a09b",
X"34e00b87",
X"a88934a2",
X"0b87a880",
X"34830b87",
X"a48f3482",
X"0b87a881",
X"34863d0d",
X"04fd3d0d",
X"83a08054",
X"805383c7",
X"c4085283",
X"c7c00851",
X"fdbf3f80",
X"d0805483",
X"b0805383",
X"c7c40852",
X"83c7c008",
X"51fdaa3f",
X"a05483a0",
X"805383c7",
X"c4085283",
X"c7c00851",
X"fd973fa0",
X"5483a480",
X"5383c7c4",
X"085283c7",
X"c00851fd",
X"843f9054",
X"83a88053",
X"83c7c408",
X"5283c7c0",
X"0851fcf1",
X"3f83c7c8",
X"3387a681",
X"34853d0d",
X"04803d0d",
X"90809008",
X"810683c0",
X"800c823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087081",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fd0676",
X"1007720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870822c",
X"bf0683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe830676",
X"822b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087088",
X"2c870683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f1ff06",
X"76882b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"8b2cbf06",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f88f",
X"ff06768b",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870912c",
X"bf0683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fc87ffff",
X"0676912b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70992c81",
X"0683c080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870ff",
X"bf0a0676",
X"992b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"80087088",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"892c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708a2c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708b2c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708c",
X"2cbf0683",
X"c0800c51",
X"823d0d04",
X"fe3d0d74",
X"81e62987",
X"2a9080a0",
X"0c843d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727081",
X"055434ff",
X"1151f039",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708405",
X"540cff11",
X"51f03984",
X"3d0d04fe",
X"3d0d8480",
X"80538052",
X"88800a51",
X"ffb33f81",
X"80805380",
X"5282800a",
X"51c63f84",
X"3d0d0480",
X"3d0d8151",
X"fbfc3f72",
X"802e9038",
X"8051fdfe",
X"3fcd3f83",
X"c7cc3351",
X"fdf43f81",
X"51fc8d3f",
X"8051fc88",
X"3f8051fb",
X"d93f823d",
X"0d04fd3d",
X"0d755280",
X"5480ff72",
X"25883881",
X"0bff8013",
X"5354ffbf",
X"12517099",
X"268638e0",
X"12529e39",
X"ff9f1251",
X"99712795",
X"38d012e0",
X"13705454",
X"51897127",
X"88388f73",
X"27833880",
X"5273802e",
X"85388180",
X"12527181",
X"ff0683c0",
X"800c853d",
X"0d04803d",
X"0d84d8c0",
X"51807170",
X"81055334",
X"7084e0c0",
X"2e098106",
X"f038823d",
X"0d04fe3d",
X"0d029705",
X"3351ff86",
X"3f83c080",
X"0881ff06",
X"83c7d008",
X"54528073",
X"249b3883",
X"c8800813",
X"7283c884",
X"08075353",
X"71733483",
X"c7d00881",
X"0583c7d0",
X"0c843d0d",
X"04fa3d0d",
X"82800a1b",
X"55805788",
X"3dfc0554",
X"79537452",
X"7851ffbb",
X"893f883d",
X"0d04fe3d",
X"0d83c7e8",
X"08527451",
X"c1ed3f83",
X"c080088c",
X"38765375",
X"5283c7e8",
X"0851c63f",
X"843d0d04",
X"fe3d0d83",
X"c7e80853",
X"75527451",
X"ffbcab3f",
X"83c08008",
X"8d387753",
X"765283c7",
X"e80851ff",
X"a03f843d",
X"0d04fe3d",
X"0d83c7e8",
X"0851ffbb",
X"9e3f83c0",
X"80088180",
X"802e0981",
X"06883883",
X"c1808053",
X"9c3983c7",
X"e80851ff",
X"bb813f83",
X"c0800880",
X"d0802e09",
X"81069338",
X"83c1b080",
X"5383c080",
X"085283c7",
X"e80851fe",
X"d43f843d",
X"0d04803d",
X"0df9e03f",
X"83c08008",
X"842981db",
X"dc057008",
X"83c0800c",
X"51823d0d",
X"04ed3d0d",
X"80448043",
X"80428041",
X"80705a5b",
X"fdcc3f80",
X"0b83c7d0",
X"0c800b83",
X"c8840c81",
X"d9b451ea",
X"a53f8180",
X"0b83c884",
X"0c81d9b8",
X"51ea973f",
X"80d00b83",
X"c7d00c78",
X"30707a07",
X"80257087",
X"2b83c884",
X"0c5155f8",
X"d13f83c0",
X"80085281",
X"d9c051e9",
X"f13f80f8",
X"0b83c7d0",
X"0c788132",
X"70307072",
X"07802570",
X"872b83c8",
X"840c5156",
X"56feef3f",
X"83c08008",
X"5281d9cc",
X"51e9c73f",
X"81a00b83",
X"c7d00c78",
X"82327030",
X"70720780",
X"2570872b",
X"83c8840c",
X"515683c7",
X"e8085256",
X"ffb6a63f",
X"83c08008",
X"5281d9d4",
X"51e9973f",
X"81f00b83",
X"c7d00c81",
X"0b83c7d4",
X"5b5883c7",
X"d0088219",
X"7a327030",
X"70720780",
X"2570872b",
X"83c8840c",
X"51578e3d",
X"7055ff1b",
X"54575757",
X"9a8d3f79",
X"7084055b",
X"0851ffb5",
X"dc3f7454",
X"83c08008",
X"53775281",
X"d9dc51e8",
X"c93fa817",
X"83c7d00c",
X"81185877",
X"852e0981",
X"06ffaf38",
X"83900b83",
X"c7d00c78",
X"87327030",
X"70720780",
X"2570872b",
X"83c8840c",
X"515656f7",
X"f53f81d9",
X"ec5583c0",
X"8008802e",
X"8f3883c7",
X"e40851ff",
X"b5873f83",
X"c0800855",
X"745281d9",
X"f451e7f6",
X"3f83e00b",
X"83c7d00c",
X"78883270",
X"30707207",
X"80257087",
X"2b83c884",
X"0c515781",
X"da805255",
X"e7d43f86",
X"8da051f8",
X"ef3f8052",
X"913d7052",
X"559da73f",
X"83527451",
X"9da03f63",
X"557482fa",
X"38611959",
X"78802585",
X"38745990",
X"39887925",
X"85388859",
X"87397888",
X"2682d938",
X"78822b55",
X"81d4b815",
X"0804f5e2",
X"3f83c080",
X"08615755",
X"75812e09",
X"81068938",
X"83c08008",
X"10559039",
X"75ff2e09",
X"81068838",
X"83c08008",
X"812c5590",
X"75258538",
X"90558839",
X"74802483",
X"38815574",
X"51f5bc3f",
X"828e39f5",
X"ce3f83c0",
X"80086105",
X"55748025",
X"85388055",
X"88398675",
X"25833886",
X"557451f5",
X"c73f81ec",
X"39608738",
X"62802e81",
X"e33883c3",
X"9c0883c3",
X"980cade5",
X"0b83c3a0",
X"0c83c7e8",
X"0851d78b",
X"3ffadb3f",
X"81c63960",
X"56807625",
X"9838ad84",
X"0b83c3a0",
X"0c83c7c8",
X"15700852",
X"55d6ec3f",
X"74085292",
X"39758025",
X"923883c7",
X"c8150851",
X"ffb2f03f",
X"8052fd19",
X"51b83962",
X"802e818c",
X"3883c7c8",
X"15700883",
X"c7d40872",
X"0c83c7d4",
X"0cfd1a70",
X"5351558c",
X"883f83c0",
X"80085680",
X"518bfe3f",
X"83c08008",
X"52745188",
X"953f7552",
X"8051888e",
X"3f80d539",
X"60558075",
X"25b63883",
X"c3a40883",
X"c3980cad",
X"e50b83c3",
X"a00c83c7",
X"e40851d5",
X"f63f83c7",
X"e40851d3",
X"973f83c0",
X"800881ff",
X"06705255",
X"f4d53f74",
X"802e9d38",
X"8155a139",
X"74802594",
X"3883c7e4",
X"0851ffb1",
X"e23f8051",
X"f4b93f84",
X"39628738",
X"7a802efa",
X"83388055",
X"7483c080",
X"0c953d0d",
X"04fe3d0d",
X"83c7f051",
X"80f3c63f",
X"f4dd3f83",
X"c0800880",
X"2e863880",
X"51818a39",
X"f4e23f83",
X"c0800880",
X"fe38f582",
X"3f83c080",
X"08802eb9",
X"388151f2",
X"913f8051",
X"f4983fef",
X"853f800b",
X"83c7d00c",
X"f9a33f83",
X"c0800853",
X"ff0b83c7",
X"d00cf0f1",
X"3f7280cb",
X"3883c7cc",
X"3351f3f2",
X"3f7251f1",
X"e13f80c0",
X"39f4aa3f",
X"83c08008",
X"802eb538",
X"8151f1ce",
X"3f8051f3",
X"d53feec2",
X"3fad840b",
X"83c3a00c",
X"83c7d408",
X"51d4a03f",
X"ff0b83c7",
X"d00cf0ad",
X"3f83c7d4",
X"08528051",
X"86843f81",
X"51f59c3f",
X"843d0d04",
X"fb3d0d80",
X"5283c7f0",
X"5180e2d5",
X"3f800b83",
X"c7cc3490",
X"80805286",
X"84808051",
X"ffb4893f",
X"83c08008",
X"81973889",
X"c53f81dd",
X"bc51ffb8",
X"c83f83c0",
X"8008559c",
X"800a5480",
X"c0805381",
X"da885283",
X"c0800851",
X"f6e63f83",
X"c7e80853",
X"81da9852",
X"7451ffb3",
X"913f83c0",
X"80088438",
X"f6f43f83",
X"c7ec0853",
X"81daa452",
X"7451ffb2",
X"f93f83c0",
X"8008b638",
X"873dfc05",
X"54848080",
X"5386a880",
X"805283c7",
X"ec0851ff",
X"b1843f83",
X"c0800893",
X"38758480",
X"802e0981",
X"06893881",
X"0b83c7cc",
X"34873980",
X"0b83c7cc",
X"3483c7cc",
X"3351f1f2",
X"3f8151f3",
X"de3f92ee",
X"3f8151f3",
X"d63f8151",
X"fd8f3ffa",
X"3983c08c",
X"080283c0",
X"8c0cfb3d",
X"0d0281da",
X"b00b83c3",
X"9c0c81da",
X"b40b83c3",
X"940c81da",
X"b80b83c3",
X"a40c83c0",
X"8c08fc05",
X"0c800b83",
X"c7d40b83",
X"c08c08f8",
X"050c83c0",
X"8c08f405",
X"0cffb194",
X"3f83c080",
X"088605fc",
X"0683c08c",
X"08f0050c",
X"0283c08c",
X"08f00508",
X"310d833d",
X"7083c08c",
X"08f80508",
X"70840583",
X"c08c08f8",
X"050c0c51",
X"ffaddc3f",
X"83c08c08",
X"f4050881",
X"0583c08c",
X"08f4050c",
X"83c08c08",
X"f4050887",
X"2e098106",
X"ffab3886",
X"94808051",
X"eaf13fff",
X"0b83c7d0",
X"0c800b83",
X"c8840c84",
X"d8c00b83",
X"c8800c81",
X"51ee9b3f",
X"8151eec0",
X"3f8051ee",
X"bb3f8151",
X"eee13f81",
X"51efb63f",
X"8251ef84",
X"3f8051ef",
X"da3f8051",
X"f0843f80",
X"d0ca5280",
X"51dfd03f",
X"fcd23f83",
X"c08c08fc",
X"05080d80",
X"0b83c080",
X"0c873d0d",
X"83c08c0c",
X"04803d0d",
X"81ff5180",
X"0b83c890",
X"1234ff11",
X"5170f438",
X"823d0d04",
X"ff3d0d73",
X"70335351",
X"81113371",
X"34718112",
X"34833d0d",
X"04fb3d0d",
X"77795656",
X"80707155",
X"55527175",
X"25ac3872",
X"16703370",
X"147081ff",
X"06555151",
X"51717427",
X"89388112",
X"7081ff06",
X"53517181",
X"147083ff",
X"ff065552",
X"54747324",
X"d6387183",
X"c0800c87",
X"3d0d04fb",
X"3d0d7756",
X"d79a3f83",
X"c0800880",
X"2ef63883",
X"caac0886",
X"057081ff",
X"065253d5",
X"9c3f810b",
X"9088d434",
X"9088d433",
X"7081ff06",
X"5153728b",
X"38f9ea3f",
X"8351efb8",
X"3fea3980",
X"55741675",
X"822b5454",
X"9088c013",
X"33743481",
X"15557485",
X"2e098106",
X"e838810b",
X"9088d434",
X"753383c8",
X"90348116",
X"3383c891",
X"34821633",
X"83c89234",
X"83163383",
X"c8933484",
X"5283c890",
X"51feba3f",
X"83c08008",
X"81ff0684",
X"17335753",
X"72762e09",
X"81068c38",
X"d5c33f83",
X"c0800880",
X"2e9a3883",
X"caac08a8",
X"2e098106",
X"8938860b",
X"83caac0c",
X"8739a80b",
X"83caac0c",
X"80e451ee",
X"b33f873d",
X"0d04f43d",
X"0d7e6059",
X"55805d80",
X"75822b71",
X"83cab012",
X"0c83cac4",
X"175b5b57",
X"76793477",
X"772e83b9",
X"38765277",
X"51ffaca2",
X"3f8e3dfc",
X"05549053",
X"83ca9852",
X"7751ffab",
X"dd3f7c56",
X"75902e09",
X"81068395",
X"3883ca98",
X"51fd953f",
X"83ca9a51",
X"fd8e3f83",
X"ca9c51fd",
X"873f7683",
X"caa80c77",
X"51ffa9a9",
X"3f0b0b81",
X"d8c45283",
X"c0800851",
X"cbc03f83",
X"c0800881",
X"2e098106",
X"80d43876",
X"83cac00c",
X"820b83ca",
X"9834ff96",
X"0b83ca99",
X"347751ff",
X"abed3f83",
X"c0800855",
X"83c08008",
X"77258838",
X"83c08008",
X"8f055574",
X"842c7083",
X"ffff0670",
X"882a5851",
X"557583ca",
X"9a347483",
X"ca9b3476",
X"83ca9c34",
X"ff800b83",
X"ca9d3481",
X"903983ca",
X"983383ca",
X"99337188",
X"2b07565b",
X"7483ffff",
X"2e098106",
X"80e838fe",
X"800b83ca",
X"c00c810b",
X"83caa80c",
X"ff0b83ca",
X"9834ff0b",
X"83ca9934",
X"7751ffaa",
X"fa3f83c0",
X"800883ca",
X"c80c83c0",
X"80085583",
X"c0800880",
X"25883883",
X"c080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583ca9a",
X"347483ca",
X"9b347683",
X"ca9c34ff",
X"800b83ca",
X"9d34810b",
X"83caa734",
X"a5397485",
X"962e0981",
X"0680fe38",
X"7583cac0",
X"0c7751ff",
X"aaae3f83",
X"caa73383",
X"c0800807",
X"557483ca",
X"a73483ca",
X"a7338106",
X"5574802e",
X"83388457",
X"83ca9c33",
X"83ca9d33",
X"71882b07",
X"565c7481",
X"802e0981",
X"06a13883",
X"ca9a3383",
X"ca9b3371",
X"882b0756",
X"5bad8075",
X"27873876",
X"8207579c",
X"39768107",
X"57963974",
X"82802e09",
X"81068738",
X"76830757",
X"87397481",
X"ff268a38",
X"7783cab0",
X"1b0c7679",
X"348e3d0d",
X"04803d0d",
X"72842983",
X"cab00570",
X"0883c080",
X"0c51823d",
X"0d04fe3d",
X"0d800b83",
X"ca940c80",
X"0b83ca90",
X"0cff0b83",
X"c88c0ca8",
X"0b83caac",
X"0cae51cf",
X"e43f800b",
X"83cab054",
X"52807370",
X"8405550c",
X"81125271",
X"842e0981",
X"06ef3884",
X"3d0d04fe",
X"3d0d7402",
X"84059605",
X"22535371",
X"802e9638",
X"72708105",
X"543351cf",
X"ef3fff12",
X"7083ffff",
X"065152e7",
X"39843d0d",
X"04fe3d0d",
X"02920522",
X"5382ac51",
X"e9c63f80",
X"c351cfcc",
X"3f819651",
X"e9ba3f72",
X"5283c890",
X"51ffb43f",
X"725283c8",
X"9051f8f1",
X"3f83c080",
X"0881ff06",
X"51cfa93f",
X"843d0d04",
X"ffb13d0d",
X"80d13df8",
X"0551f99b",
X"3f83ca94",
X"08810583",
X"ca940c80",
X"cf3d33cf",
X"117081ff",
X"06515656",
X"74832688",
X"e238758f",
X"06ff0556",
X"7583c88c",
X"082e9b38",
X"75832696",
X"387583c8",
X"8c0c7584",
X"2983cab0",
X"05700853",
X"557551fa",
X"993f8076",
X"2488be38",
X"75842983",
X"cab00555",
X"7408802e",
X"88af3883",
X"c88c0884",
X"2983cab0",
X"05700802",
X"880582b9",
X"0533525b",
X"557480d2",
X"2e84ac38",
X"7480d224",
X"903874bf",
X"2e9c3874",
X"80d02e81",
X"d13887ee",
X"397480d3",
X"2e80cf38",
X"7480d72e",
X"81c03887",
X"dd390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290556",
X"56cea53f",
X"80c151cd",
X"df3ff6ed",
X"3f860b83",
X"c8903481",
X"5283c890",
X"51cf823f",
X"8151fde9",
X"3f748938",
X"860b83ca",
X"ac0c8739",
X"a80b83ca",
X"ac0ccdf4",
X"3f80c151",
X"cdae3ff6",
X"bc3f900b",
X"83caa733",
X"81065656",
X"74802e83",
X"38985683",
X"ca9c3383",
X"ca9d3371",
X"882b0756",
X"59748180",
X"2e098106",
X"9c3883ca",
X"9a3383ca",
X"9b337188",
X"2b075657",
X"ad807527",
X"8c387581",
X"80075685",
X"3975a007",
X"567583c8",
X"9034ff0b",
X"83c89134",
X"e00b83c8",
X"9234800b",
X"83c89334",
X"845283c8",
X"9051cdf9",
X"3f845186",
X"9b390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290556",
X"59cce93f",
X"7951ffa4",
X"ff3f83c0",
X"8008802e",
X"8a3880ce",
X"51cc953f",
X"85f13980",
X"c151cc8c",
X"3fcd813f",
X"cbb63f83",
X"cac00858",
X"8375259b",
X"3883ca9c",
X"3383ca9d",
X"3371882b",
X"07fc1771",
X"297a0583",
X"80055a51",
X"578d3974",
X"81802918",
X"ff800558",
X"81805780",
X"5676762e",
X"9238cbe8",
X"3f83c080",
X"0883c890",
X"17348116",
X"56eb39cb",
X"d73f83c0",
X"800881ff",
X"06775383",
X"c8905256",
X"f4e73f83",
X"c0800881",
X"ff065575",
X"752e0981",
X"06819538",
X"9451e588",
X"3fcbd13f",
X"80c151cb",
X"8b3fcc80",
X"3f775279",
X"51ffa392",
X"3f805e80",
X"d13dfdf4",
X"05547653",
X"83c89052",
X"7951ffa1",
X"9f3f0282",
X"b9053355",
X"81597480",
X"d72e0981",
X"0680c538",
X"77527951",
X"ffa2e33f",
X"80d13dfd",
X"f0055476",
X"538f3d70",
X"537a5258",
X"ffa29b3f",
X"80567676",
X"2ea23875",
X"1883c890",
X"17337133",
X"70723270",
X"30708025",
X"70307f06",
X"811d5d5f",
X"51515152",
X"5b55db39",
X"82ac51e4",
X"833f7880",
X"2e863880",
X"c3518439",
X"80ce51c9",
X"ff3fcaf4",
X"3fc9a93f",
X"83d83902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"59558070",
X"5d5980e4",
X"51e3cd3f",
X"ca963f80",
X"c151c9d0",
X"3f83caa8",
X"08792e82",
X"d63883ca",
X"c80880fc",
X"055580fd",
X"52745185",
X"a03f83c0",
X"80085b77",
X"8224b238",
X"ff187087",
X"2b83ffff",
X"800681db",
X"fc0583c8",
X"90595755",
X"81805575",
X"70810557",
X"33777081",
X"055934ff",
X"157081ff",
X"06515574",
X"ea388285",
X"397782e8",
X"2e81a338",
X"7782e92e",
X"09810681",
X"aa387858",
X"77873270",
X"30707207",
X"80257a8a",
X"32703070",
X"72078025",
X"73075354",
X"5a515755",
X"75802e97",
X"38787826",
X"9238a00b",
X"83c8901a",
X"34811970",
X"81ff065a",
X"55eb3981",
X"187081ff",
X"0659558a",
X"7827ffbc",
X"388f5883",
X"c88b1833",
X"83c89019",
X"34ff1870",
X"81ff0659",
X"55778426",
X"ea389058",
X"800b83c8",
X"90193481",
X"187081ff",
X"0670982b",
X"52595574",
X"8025e938",
X"80c6557a",
X"858f2484",
X"3880c255",
X"7483c890",
X"3480f10b",
X"83c89334",
X"810b83c8",
X"94347a83",
X"c891347a",
X"882c5574",
X"83c89234",
X"80cb3982",
X"f0782580",
X"c4387780",
X"fd29fd97",
X"d3055279",
X"51ff9fbe",
X"3f80d13d",
X"fdec0554",
X"80fd5383",
X"c8905279",
X"51ff9ef6",
X"3f7b8119",
X"59567580",
X"fc248338",
X"78587788",
X"2c557483",
X"c98d3477",
X"83c98e34",
X"7583c98f",
X"34818059",
X"80cc3983",
X"cac00857",
X"8378259b",
X"3883ca9c",
X"3383ca9d",
X"3371882b",
X"07fc1a71",
X"29790583",
X"80055951",
X"598d3977",
X"81802917",
X"ff800557",
X"81805976",
X"527951ff",
X"9ecc3f80",
X"d13dfdec",
X"05547853",
X"83c89052",
X"7951ff9e",
X"853f7851",
X"f6c33fc7",
X"973fc5cc",
X"3f8b3983",
X"ca900881",
X"0583ca90",
X"0c80d13d",
X"0d04f6e4",
X"3ffc39fc",
X"3d0d7678",
X"71842983",
X"cab00570",
X"08515353",
X"53709e38",
X"80ce7234",
X"80cf0b81",
X"133480ce",
X"0b821334",
X"80c50b83",
X"13347084",
X"133480e7",
X"3983cac4",
X"13335480",
X"d2723473",
X"822a7081",
X"06515180",
X"cf537084",
X"3880d753",
X"72811334",
X"a00b8213",
X"34738306",
X"5170812e",
X"9e387081",
X"24883870",
X"802e8f38",
X"9f397082",
X"2e923870",
X"832e9238",
X"933980d8",
X"558e3980",
X"d3558939",
X"80cd5584",
X"3980c455",
X"74831334",
X"80c40b84",
X"1334800b",
X"85133486",
X"3d0d04fc",
X"3d0d7678",
X"53548153",
X"80558739",
X"71107310",
X"54527372",
X"26517280",
X"2ea73870",
X"802e8638",
X"718025e8",
X"3872802e",
X"98387174",
X"26893873",
X"72317574",
X"07565472",
X"812a7281",
X"2a5353e5",
X"39735178",
X"83387451",
X"7083c080",
X"0c863d0d",
X"04fe3d0d",
X"80537552",
X"7451ffa3",
X"3f843d0d",
X"04fe3d0d",
X"81537552",
X"7451ff93",
X"3f843d0d",
X"04fb3d0d",
X"77795555",
X"80567476",
X"25863874",
X"30558156",
X"73802588",
X"38733076",
X"81325754",
X"80537352",
X"7451fee7",
X"3f83c080",
X"08547580",
X"2e873883",
X"c0800830",
X"547383c0",
X"800c873d",
X"0d04fa3d",
X"0d787a57",
X"55805774",
X"77258638",
X"74305581",
X"57759f2c",
X"54815375",
X"74327431",
X"527451fe",
X"aa3f83c0",
X"80085476",
X"802e8738",
X"83c08008",
X"30547383",
X"c0800c88",
X"3d0d04fc",
X"3d0d7655",
X"80750c80",
X"0b84160c",
X"800b8816",
X"0c800b8c",
X"160c83c7",
X"f05180da",
X"cc3f87a6",
X"80337081",
X"ff065152",
X"dcad3f71",
X"812a8132",
X"72813271",
X"81067181",
X"06318418",
X"0c545471",
X"832a8132",
X"72822a81",
X"32718106",
X"71810631",
X"770c5353",
X"87a09033",
X"70098106",
X"88170c52",
X"83c08008",
X"802e80c2",
X"3883c080",
X"08812a70",
X"810683c0",
X"80088106",
X"3184170c",
X"5283c080",
X"08832a83",
X"c0800882",
X"2a718106",
X"71810631",
X"770c5353",
X"83c08008",
X"842a8106",
X"88160c83",
X"c0800885",
X"2a81068c",
X"160c863d",
X"0d04fe3d",
X"0d747654",
X"527151fe",
X"c63f7281",
X"2ea23881",
X"73268d38",
X"72822ea8",
X"3872832e",
X"9c38e639",
X"7108e238",
X"841208dd",
X"38881208",
X"d838a539",
X"88120881",
X"2e9e3891",
X"39881208",
X"812e9538",
X"71089138",
X"8412088c",
X"388c1208",
X"812e0981",
X"06ffb238",
X"843d0d04",
X"fb3d0d78",
X"0284059f",
X"05335556",
X"800b81d6",
X"c8565381",
X"732b7406",
X"5271802e",
X"83388152",
X"74708205",
X"56227073",
X"902b0790",
X"809c0c51",
X"81135372",
X"882e0981",
X"06d93880",
X"5383cad0",
X"13335170",
X"81ff2eb2",
X"38701081",
X"d4e80570",
X"22555180",
X"73177033",
X"701081d4",
X"e8057022",
X"51515152",
X"5273712e",
X"91388112",
X"5271862e",
X"098106f1",
X"38739080",
X"9c0c8113",
X"5372862e",
X"098106ff",
X"b8388053",
X"72167033",
X"51517081",
X"ff2e9438",
X"701081d4",
X"e8057022",
X"70848080",
X"0790809c",
X"0c515181",
X"13537286",
X"2e098106",
X"d7388053",
X"72165170",
X"3383cad0",
X"14348113",
X"5372862e",
X"098106ec",
X"38873d0d",
X"0404ff3d",
X"0d740284",
X"058f0533",
X"52527088",
X"38719080",
X"940c8e39",
X"70812e09",
X"81068638",
X"71908098",
X"0c833d0d",
X"04fb3d0d",
X"029f0533",
X"79982b70",
X"982c7c98",
X"2b70982c",
X"83caec15",
X"70337098",
X"2b70982c",
X"51585c5a",
X"51555154",
X"5470732e",
X"09810694",
X"3883cacc",
X"14337098",
X"2b70982c",
X"51525670",
X"722eb138",
X"72753471",
X"83cacc15",
X"3483cacd",
X"3383caed",
X"3371982b",
X"71902b07",
X"83cacc33",
X"70882b72",
X"0783caec",
X"33710790",
X"80b80c52",
X"59535452",
X"873d0d04",
X"fe3d0d74",
X"81113371",
X"3371882b",
X"0783c080",
X"0c535184",
X"3d0d0483",
X"cad83383",
X"c0800c04",
X"f53d0d02",
X"bb053302",
X"8405bf05",
X"33028805",
X"80c30533",
X"028c0580",
X"c6052266",
X"5c5a5e5c",
X"567a557b",
X"548953a1",
X"527d5180",
X"d0c03f83",
X"c0800881",
X"ff0683c0",
X"800c8d3d",
X"0d0483c0",
X"8c080283",
X"c08c0cf5",
X"3d0d83c0",
X"8c088805",
X"0883c08c",
X"088f0533",
X"83c08c08",
X"92052202",
X"8c057390",
X"0583c08c",
X"08e8050c",
X"83c08c08",
X"f8050c83",
X"c08c08f0",
X"050c83c0",
X"8c08ec05",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08f005",
X"0883c08c",
X"08e0050c",
X"83c08c08",
X"fc050c83",
X"c08c08f0",
X"05088927",
X"8a38890b",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"05088605",
X"87fffc06",
X"83c08c08",
X"e0050c02",
X"83c08c08",
X"e0050831",
X"0d853d70",
X"5583c08c",
X"08ec0508",
X"5483c08c",
X"08f00508",
X"5383c08c",
X"08f40508",
X"5283c08c",
X"08e4050c",
X"80d9f23f",
X"83c08008",
X"81ff0683",
X"c08c08e4",
X"050883c0",
X"8c08ec05",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"e0050880",
X"2e8c3883",
X"c08c08f8",
X"05080d89",
X"c83983c0",
X"8c08f005",
X"08802e89",
X"a63883c0",
X"8c08ec05",
X"08810533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508842e",
X"a938840b",
X"83c08c08",
X"e0050825",
X"88c73883",
X"c08c08e0",
X"0508852e",
X"859b3883",
X"c08c08e0",
X"0508a12e",
X"87ad3888",
X"ac39800b",
X"83c08c08",
X"ec050885",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08fc050c",
X"83c08c08",
X"e0050883",
X"2e098106",
X"88833883",
X"c08c08e8",
X"05088105",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e0050881",
X"2687e638",
X"810b83c0",
X"8c08e005",
X"0880d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08fc",
X"050c83c0",
X"8c08ec05",
X"08820533",
X"83c08c08",
X"e0050887",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088b",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"e005088c",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088d",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"e005088e",
X"052383c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088a",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"70940508",
X"fcffff06",
X"7194050c",
X"83c08c08",
X"e0050c83",
X"c08c08ec",
X"05088605",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"f4050c83",
X"c08c08e0",
X"050883c0",
X"8c08fc05",
X"082e0981",
X"06b63883",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c83",
X"c08c08fc",
X"050883c0",
X"8c08e005",
X"088b0534",
X"83c08c08",
X"ec050887",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"812e8f38",
X"83c08c08",
X"e0050882",
X"2eb73884",
X"8c3983c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c820b",
X"83c08c08",
X"e005088a",
X"053483d9",
X"3983c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08fc0508",
X"83c08c08",
X"e005088a",
X"053483a1",
X"3983c08c",
X"08fc0508",
X"802e8395",
X"3883c08c",
X"08ec0508",
X"83053383",
X"0683c08c",
X"08e0050c",
X"83c08c08",
X"e0050883",
X"2e098106",
X"82f33883",
X"c08c08ec",
X"05088205",
X"3370982b",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c83c0",
X"8c08e005",
X"08802582",
X"cc3883c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c83c0",
X"8c08ec05",
X"08860533",
X"83c08c08",
X"e0050880",
X"d6053483",
X"c08c08e0",
X"05088405",
X"83c08c08",
X"ec050882",
X"05338f06",
X"83c08c08",
X"e4050c83",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0883c08c",
X"08e00508",
X"3483c08c",
X"08ec0508",
X"84053383",
X"c08c08e0",
X"05088105",
X"34800b83",
X"c08c08e0",
X"05088205",
X"3483c08c",
X"08e00508",
X"08ff83ff",
X"06828007",
X"83c08c08",
X"e005080c",
X"83c08c08",
X"e8050881",
X"05338105",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"050883c0",
X"8c08e805",
X"08810534",
X"81833983",
X"c08c08fc",
X"0508802e",
X"80f73883",
X"c08c08ec",
X"05088605",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e00508a2",
X"2e098106",
X"80d73883",
X"c08c08ec",
X"05088805",
X"3383c08c",
X"08ec0508",
X"87053371",
X"82802905",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c5283c0",
X"8c08e405",
X"0c83c08c",
X"08f4050c",
X"83c08c08",
X"e4050883",
X"c08c08e0",
X"05088805",
X"2383c08c",
X"08ec0508",
X"3383c08c",
X"08f00508",
X"71317083",
X"ffff0683",
X"c08c08f0",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08ec0508",
X"0583c08c",
X"08ec050c",
X"f6d03983",
X"c08c08f8",
X"05080d83",
X"c08c08f0",
X"050883c0",
X"8c08e005",
X"0c83c08c",
X"08f80508",
X"0d83c08c",
X"08e00508",
X"83c0800c",
X"8d3d0d83",
X"c08c0c04",
X"83c08c08",
X"0283c08c",
X"0ce63d0d",
X"83c08c08",
X"88050802",
X"840583c0",
X"8c08e805",
X"0c83c08c",
X"08d4050c",
X"800b83ca",
X"f43483c0",
X"8c08d405",
X"08900583",
X"c08c08c0",
X"050c800b",
X"83c08c08",
X"c0050834",
X"800b83c0",
X"8c08c005",
X"08810534",
X"800b83c0",
X"8c08c405",
X"0c83c08c",
X"08c40508",
X"80d82983",
X"c08c08c0",
X"05080583",
X"c08c08ff",
X"b4050c80",
X"0b83c08c",
X"08ffb405",
X"0880d805",
X"0c83c08c",
X"08ffb405",
X"08840583",
X"c08c08ff",
X"b4050c83",
X"c08c08c4",
X"050883c0",
X"8c08ffb4",
X"05083488",
X"0b83c08c",
X"08ffb405",
X"08810534",
X"800b83c0",
X"8c08ffb4",
X"05088205",
X"3483c08c",
X"08ffb405",
X"0808ffa1",
X"ff06a080",
X"0783c08c",
X"08ffb405",
X"080c83c0",
X"8c08c405",
X"08810570",
X"81ff0683",
X"c08c08c4",
X"050c83c0",
X"8c08ffb4",
X"050c810b",
X"83c08c08",
X"c4050827",
X"fedb3883",
X"c08c08ec",
X"05705483",
X"c08c08c8",
X"050c9252",
X"83c08c08",
X"d4050851",
X"80cd993f",
X"83c08008",
X"81ff0670",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"8dea3883",
X"c08c08f4",
X"0551f18c",
X"3f83c080",
X"0883ffff",
X"0683c08c",
X"08f60552",
X"83c08c08",
X"e4050cf0",
X"f33f83c0",
X"800883ff",
X"ff0683c0",
X"8c08fd05",
X"3383c08c",
X"08ffb805",
X"0883c08c",
X"08c4050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"e0050c83",
X"c08c08c4",
X"050883c0",
X"8c08ffbc",
X"05082780",
X"fe3883c0",
X"8c08c805",
X"085483c0",
X"8c08c405",
X"08538952",
X"83c08c08",
X"d4050851",
X"80cc9e3f",
X"83c08008",
X"81ff0683",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b8050880",
X"f23883c0",
X"8c08ee05",
X"51eff13f",
X"83c08008",
X"83ffff06",
X"5383c08c",
X"08c40508",
X"5283c08c",
X"08d40508",
X"51f0b33f",
X"83c08c08",
X"c4050881",
X"057081ff",
X"0683c08c",
X"08c4050c",
X"83c08c08",
X"ffb4050c",
X"fef13983",
X"c08c08c0",
X"05088105",
X"3383c08c",
X"08ffb405",
X"0c81db0b",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb40508",
X"802e8be0",
X"38943983",
X"c08c08ff",
X"b8050883",
X"c08c08ff",
X"bc050c8b",
X"cb3983c0",
X"8c08f105",
X"335283c0",
X"8c08d405",
X"085180cb",
X"9c3f800b",
X"83c08c08",
X"c0050881",
X"053383c0",
X"8c08ffb4",
X"050c83c0",
X"8c08c405",
X"0c83c08c",
X"08c40508",
X"83c08c08",
X"ffb40508",
X"2789e638",
X"83c08c08",
X"c4050880",
X"d8297083",
X"c08c08c0",
X"05080570",
X"88057083",
X"053383c0",
X"8c08cc05",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"d8050c83",
X"c08c08cc",
X"050887a6",
X"3883c08c",
X"08c80508",
X"22028405",
X"71860587",
X"fffc0683",
X"c08c08ff",
X"b4050c83",
X"c08c08dc",
X"050c83c0",
X"8c08ffb8",
X"050c0283",
X"c08c08ff",
X"b4050831",
X"0d893d70",
X"5983c08c",
X"08ffb805",
X"085883c0",
X"8c08ffbc",
X"05088705",
X"335783c0",
X"8c08ffb4",
X"050ca255",
X"83c08c08",
X"cc050854",
X"86538181",
X"5283c08c",
X"08d40508",
X"51be933f",
X"83c08008",
X"81ff0683",
X"c08c08d0",
X"050c83c0",
X"8c08d005",
X"0881c138",
X"83c08c08",
X"ffbc0508",
X"96055383",
X"c08c08ff",
X"b8050852",
X"83c08c08",
X"ffb40508",
X"51a1c63f",
X"83c08008",
X"81ff0683",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b4050880",
X"2e818538",
X"83c08c08",
X"ffbc0508",
X"940583c0",
X"8c08ffbc",
X"05089605",
X"3370862a",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"cc050c83",
X"c08c08ff",
X"b4050883",
X"2e098106",
X"80c63883",
X"c08c08ff",
X"b4050883",
X"c08c08c8",
X"05088205",
X"3483cad8",
X"33708105",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb40508",
X"83cad834",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"cc050834",
X"83c08c08",
X"dc05080d",
X"83c08c08",
X"d0050881",
X"ff0683c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"0508fbff",
X"3883c08c",
X"08d80508",
X"83c08c08",
X"c0050805",
X"88057082",
X"05335183",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b4050883",
X"2e098106",
X"80e33883",
X"c08c08ff",
X"b8050883",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b4050881",
X"057081ff",
X"065183c0",
X"8c08ffb4",
X"050c810b",
X"83c08c08",
X"ffb40508",
X"27dd3880",
X"0b83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb405",
X"08810570",
X"81ff0651",
X"83c08c08",
X"ffb4050c",
X"970b83c0",
X"8c08ffb4",
X"050827dd",
X"3883c08c",
X"08e40508",
X"80f93270",
X"30708025",
X"515183c0",
X"8c08ffb4",
X"050c83c0",
X"8c08e005",
X"08912e09",
X"810680f9",
X"3883c08c",
X"08ffb405",
X"08802e80",
X"ec3883c0",
X"8c08c405",
X"0880e238",
X"850b83c0",
X"8c08c005",
X"08a60534",
X"a00b83c0",
X"8c08c005",
X"08a70534",
X"850b83c0",
X"8c08c005",
X"08a80534",
X"80c00b83",
X"c08c08c0",
X"0508a905",
X"34860b83",
X"c08c08c0",
X"0508aa05",
X"34900b83",
X"c08c08c0",
X"0508ab05",
X"34860b83",
X"c08c08c0",
X"0508ac05",
X"34a00b83",
X"c08c08c0",
X"0508ad05",
X"3483c08c",
X"08e40508",
X"89d83270",
X"30708025",
X"515183c0",
X"8c08ffb4",
X"050c83c0",
X"8c08e005",
X"0883edec",
X"2e098106",
X"80f63881",
X"7083c08c",
X"08ffb405",
X"080683c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb4",
X"0508802e",
X"80ce3883",
X"c08c08c4",
X"050880c4",
X"38840b83",
X"c08c08c0",
X"0508aa05",
X"3480c00b",
X"83c08c08",
X"c00508ab",
X"0534840b",
X"83c08c08",
X"c00508ac",
X"0534900b",
X"83c08c08",
X"c00508ad",
X"053483c0",
X"8c08ffb8",
X"050883c0",
X"8c08c005",
X"088c0534",
X"83c08c08",
X"e4050880",
X"f9327030",
X"70802551",
X"5183c08c",
X"08ffb405",
X"0c83c08c",
X"08e00508",
X"862e0981",
X"0680c338",
X"817083c0",
X"8c08ffb4",
X"05080683",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b4050880",
X"2e9c3883",
X"c08c08c4",
X"05089338",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"c005088d",
X"053483c0",
X"8c08c405",
X"0880d829",
X"83c08c08",
X"c0050805",
X"70840570",
X"83053383",
X"c08c08ff",
X"b4050c83",
X"c08c08c8",
X"050c83c0",
X"8c08ffbc",
X"050c8058",
X"805783c0",
X"8c08ffb4",
X"05085680",
X"5580548a",
X"53a15283",
X"c08c08d4",
X"050851b7",
X"8d3f83c0",
X"800881ff",
X"06703070",
X"9f2a5183",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b80508a0",
X"2e8c3883",
X"c08c08ff",
X"b40508f6",
X"c23883c0",
X"8c08ffbc",
X"05088b05",
X"3383c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb405",
X"08802eb3",
X"3883c08c",
X"08c80508",
X"83053383",
X"c08c08ff",
X"b4050c80",
X"58805783",
X"c08c08ff",
X"b4050856",
X"80558054",
X"8b53a152",
X"83c08c08",
X"d4050851",
X"b6883f83",
X"c08c08c4",
X"05088105",
X"7081ff06",
X"83c08c08",
X"c0050881",
X"05335283",
X"c08c08c4",
X"050c83c0",
X"8c08ffb4",
X"050cf689",
X"39800b83",
X"c08c08c4",
X"050c83c0",
X"8c08c405",
X"0880d829",
X"83c08c08",
X"d4050805",
X"709a0533",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb40508",
X"822e0981",
X"06a93883",
X"caf45681",
X"55805483",
X"c08c08ff",
X"b4050853",
X"83c08c08",
X"ffb80508",
X"97053352",
X"83c08c08",
X"d4050851",
X"e48a3f83",
X"c08c08c4",
X"05088105",
X"7081ff06",
X"83c08c08",
X"c4050c83",
X"c08c08ff",
X"b4050c81",
X"0b83c08c",
X"08c40508",
X"27fefb38",
X"810b83c0",
X"8c08c005",
X"0834800b",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"e805080d",
X"83c08c08",
X"ffbc0508",
X"83c0800c",
X"9c3d0d83",
X"c08c0c04",
X"f53d0d90",
X"1e57800b",
X"81183354",
X"59787327",
X"819d3878",
X"80d82917",
X"8a113354",
X"5472832e",
X"09810680",
X"f8389414",
X"335ba98c",
X"3f83c080",
X"085a8056",
X"7581c429",
X"1a871133",
X"54547280",
X"2e80c038",
X"730881d4",
X"dc2e0981",
X"06b53880",
X"74595574",
X"80d82918",
X"9a113354",
X"5472832e",
X"09810692",
X"38a41470",
X"3354547a",
X"73278738",
X"ff135372",
X"74348115",
X"7081ff06",
X"56538175",
X"27d13881",
X"167081ff",
X"0657538f",
X"7627ffa4",
X"3883cad8",
X"33ff0553",
X"7283cad8",
X"34811970",
X"81ff0681",
X"19335e5a",
X"537b7926",
X"fee53880",
X"0b83c080",
X"0c8d3d0d",
X"0483c08c",
X"080283c0",
X"8c0ce63d",
X"0d83c08c",
X"08880508",
X"02840571",
X"90057033",
X"7083c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"dc050c83",
X"c08c08e0",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"94b53880",
X"0b83c08c",
X"08c80508",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08d4",
X"050c83c0",
X"8c08d405",
X"0883c08c",
X"08ffa405",
X"082593fd",
X"3883c08c",
X"08d40508",
X"80d82983",
X"c08c08c8",
X"05080584",
X"05708605",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffa405",
X"08802e93",
X"8938a6b2",
X"3f83c08c",
X"08ffb805",
X"0880d405",
X"0883c080",
X"082692f2",
X"380283c0",
X"8c08ffb8",
X"05088105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08d8050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"fc052383",
X"c08c08ff",
X"a4050886",
X"0583fc06",
X"83c08c08",
X"ffa4050c",
X"0283c08c",
X"08ffa405",
X"08310d85",
X"3d705583",
X"c08c08fc",
X"055483c0",
X"8c08ffb8",
X"05085383",
X"c08c08e0",
X"05085283",
X"c08c08c0",
X"050cae8a",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"91bb3883",
X"c08c08ff",
X"b8050887",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"80d53883",
X"c08c08ff",
X"b8050886",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508822e",
X"098106b3",
X"3883c08c",
X"08fc0522",
X"83c08c08",
X"ffa4050c",
X"870b83c0",
X"8c08ffa4",
X"05082797",
X"3883c08c",
X"08c00508",
X"82055283",
X"c08c08c0",
X"05083351",
X"dba63f83",
X"c08c08ff",
X"b8050886",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508832e",
X"09810690",
X"a43883c0",
X"8c08ffb8",
X"05089205",
X"70820533",
X"83c08c08",
X"fc052283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08c4",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffa8",
X"0508268f",
X"e438800b",
X"83c08c08",
X"e4050c80",
X"0b83c08c",
X"08ffb005",
X"0c83c08c",
X"08ffb005",
X"081083c0",
X"8c0805f8",
X"0583c08c",
X"08ffb005",
X"08842983",
X"c08c08ff",
X"b0050810",
X"0583c08c",
X"08c40508",
X"05708405",
X"703383c0",
X"8c08c005",
X"08057033",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffbc0508",
X"2383c08c",
X"08ffa805",
X"08810533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"902e0981",
X"06be3883",
X"c08c08ff",
X"a8050833",
X"83c08c08",
X"c0050805",
X"81057033",
X"70828029",
X"83c08c08",
X"ffb40508",
X"05515183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"bc050823",
X"83c08c08",
X"ffac0508",
X"86052283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a80508a2",
X"3883c08c",
X"08ffac05",
X"08880522",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"81ff2e80",
X"e53883c0",
X"8c08ffbc",
X"05082270",
X"83c08c08",
X"ffa80508",
X"31708280",
X"29713183",
X"c08c08ff",
X"ac050888",
X"05227083",
X"c08c08ff",
X"a8050831",
X"70733553",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffbc05",
X"082383c0",
X"8c08ffb0",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa4050c",
X"810b83c0",
X"8c08ffb0",
X"050827fc",
X"e03883c0",
X"8c08f805",
X"2283c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08bf2691",
X"3883c08c",
X"08e40508",
X"820783c0",
X"8c08e405",
X"0c81c00b",
X"83c08c08",
X"ffa40508",
X"27913883",
X"c08c08e4",
X"05088107",
X"83c08c08",
X"e4050c83",
X"c08c08fa",
X"052283c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508bf26",
X"913883c0",
X"8c08e405",
X"08880783",
X"c08c08e4",
X"050c81c0",
X"0b83c08c",
X"08ffa405",
X"08279138",
X"83c08c08",
X"e4050884",
X"0783c08c",
X"08e4050c",
X"800b83c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffb0",
X"05081083",
X"c08c08c4",
X"05080570",
X"90057033",
X"83c08c08",
X"c0050805",
X"70337281",
X"05337072",
X"06515351",
X"83c08c08",
X"ffa8050c",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e9b",
X"38900b83",
X"c08c08ff",
X"b005082b",
X"83c08c08",
X"e4050807",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"b0050881",
X"057081ff",
X"0683c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa405",
X"0c970b83",
X"c08c08ff",
X"b0050827",
X"fef43883",
X"c08c08ff",
X"b8050890",
X"053383c0",
X"8c08e405",
X"0883c08c",
X"08ffb405",
X"0c83c08c",
X"08c4050c",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffb80508",
X"8c05082e",
X"83ff3883",
X"c08c08ff",
X"b4050883",
X"c08c08ff",
X"b805088c",
X"050c83c0",
X"8c08ffb8",
X"05088905",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e83",
X"b93883c0",
X"8c08e405",
X"83c08c08",
X"ffb40508",
X"8f0683c0",
X"8c08e405",
X"0c83c08c",
X"08cc050c",
X"800b83c0",
X"8c08f005",
X"0c800b83",
X"c08c08f4",
X"0523800b",
X"81d6d833",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffbc0508",
X"2e82d338",
X"83c08c08",
X"f00581d6",
X"d80b83c0",
X"8c08ffac",
X"050c83c0",
X"8c08d005",
X"0c83c08c",
X"08ffac05",
X"083383c0",
X"8c08ffac",
X"05088105",
X"3381722b",
X"81722b07",
X"7083c08c",
X"08ffb405",
X"08065283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"a805082e",
X"09810681",
X"be3883c0",
X"8c08ffbc",
X"05088526",
X"80f63883",
X"c08c08ff",
X"ac050882",
X"05337081",
X"ff0683c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"80ca3883",
X"c08c08ff",
X"bc050883",
X"c08c08ff",
X"bc050881",
X"057081ff",
X"0683c08c",
X"08d00508",
X"73055383",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b0050883",
X"c08c08ff",
X"a4050834",
X"83c08c08",
X"ffac0508",
X"83053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e9d3881",
X"0b83c08c",
X"08ffa405",
X"082b83c0",
X"8c08cc05",
X"08080783",
X"c08c08cc",
X"05080c83",
X"c08c08ff",
X"ac050884",
X"05703383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a40508fd",
X"c83883c0",
X"8c08f005",
X"528051d0",
X"c33f83c0",
X"8c08e405",
X"085283c0",
X"8c08c405",
X"0851d1fe",
X"3f83c08c",
X"08fb0533",
X"7081800a",
X"29810a05",
X"70982c55",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"f9053370",
X"81800a29",
X"810a0570",
X"982c5583",
X"c08c08ff",
X"a4050c83",
X"c08c08c4",
X"05085383",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a8050cd1",
X"d43f83c0",
X"8c08ffb8",
X"05088805",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e84",
X"e03883c0",
X"8c08ffb8",
X"05089005",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08812684",
X"c0388070",
X"81d78c0b",
X"81d78c0b",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"b405082e",
X"81ae3883",
X"c08c08ff",
X"ac050884",
X"2983c08c",
X"08ffa805",
X"08057033",
X"83c08c08",
X"c0050805",
X"70337281",
X"05337072",
X"06515351",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802eaa38",
X"810b83c0",
X"8c08ffac",
X"05082b83",
X"c08c08ff",
X"b4050807",
X"7083ffff",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffac05",
X"08810570",
X"81ff0681",
X"d78c7184",
X"29710570",
X"81053351",
X"5383c08c",
X"08ffa805",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08fed438",
X"83c08c08",
X"ffb80508",
X"8a052283",
X"c08c08c0",
X"050c83c0",
X"8c08ffb4",
X"050883c0",
X"8c08c005",
X"082e82ad",
X"38800b83",
X"c08c08e8",
X"050c800b",
X"83c08c08",
X"ec052380",
X"7083c08c",
X"08e80583",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"b0050c81",
X"af3983c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffac",
X"05082c70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e80e738",
X"83c08c08",
X"ffb00508",
X"83c08c08",
X"ffb00508",
X"81057081",
X"ff0683c0",
X"8c08ffbc",
X"05087305",
X"83c08c08",
X"ffb80508",
X"90053383",
X"c08c08ff",
X"ac050884",
X"29055353",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa80508",
X"81d78e05",
X"3383c08c",
X"08ffa405",
X"083483c0",
X"8c08ffac",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa4050c",
X"8f0b83c0",
X"8c08ffac",
X"05082783",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b0050885",
X"268c3883",
X"c08c08ff",
X"a40508fe",
X"a93883c0",
X"8c08e805",
X"528051ca",
X"f33f83c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffb8",
X"05088a05",
X"2383c08c",
X"08ffb805",
X"0880d205",
X"3383c08c",
X"08ffb805",
X"0880d405",
X"080583c0",
X"8c08ffb8",
X"050880d4",
X"050c83c0",
X"8c08d805",
X"080d83c0",
X"8c08d405",
X"0881800a",
X"2981800a",
X"0570982c",
X"83c08c08",
X"c8050881",
X"053383c0",
X"8c08ffa8",
X"050c5183",
X"c08c08d4",
X"050c83c0",
X"8c08ffa8",
X"050883c0",
X"8c08d405",
X"0824ec85",
X"38800b83",
X"c08c08ff",
X"a8050c83",
X"c08c08dc",
X"05080d83",
X"c08c08ff",
X"a8050883",
X"c0800c9c",
X"3d0d83c0",
X"8c0c04f3",
X"3d0d02bf",
X"05330284",
X"0580c305",
X"3383caf4",
X"335a5b59",
X"79802e8d",
X"38787806",
X"5776802e",
X"8e388189",
X"39787806",
X"5776802e",
X"80ff3883",
X"caf43370",
X"7a075858",
X"79883878",
X"09707906",
X"51577683",
X"caf43492",
X"973f83c0",
X"80085e80",
X"5c8f5d7d",
X"1c871133",
X"58587680",
X"2e80c138",
X"770881d4",
X"dc2e0981",
X"06b63880",
X"5b815a7d",
X"1c701c9a",
X"11335959",
X"5976822e",
X"09810694",
X"3883caf4",
X"56815580",
X"54765397",
X"18335278",
X"51cbc53f",
X"ff1a80d8",
X"1c5c5a79",
X"8025d038",
X"ff1d81c4",
X"1d5d5d7c",
X"8025ffa7",
X"388f3d0d",
X"04e93d0d",
X"696c0288",
X"0580ea05",
X"225c5a5b",
X"80707141",
X"5e58ff78",
X"797a7b7c",
X"7d464c4a",
X"45405d43",
X"62993d34",
X"62028405",
X"80dd0534",
X"77792280",
X"ffff0654",
X"45727923",
X"79782e88",
X"87387a70",
X"81055c33",
X"70842a71",
X"8c067082",
X"2a5a5656",
X"8306ff1b",
X"7083ffff",
X"065c5456",
X"80547574",
X"2e91387a",
X"7081055c",
X"33ff1b70",
X"83ffff06",
X"5c545481",
X"76279b38",
X"7381ff06",
X"7b708105",
X"5d335574",
X"82802905",
X"ff1b7083",
X"ffff065c",
X"54548276",
X"27aa3873",
X"83ffff06",
X"7b708105",
X"5d337090",
X"2b72077d",
X"7081055f",
X"3370982b",
X"7207fe1f",
X"7083ffff",
X"06405252",
X"52525454",
X"7e802e80",
X"c4387686",
X"f738748a",
X"2e098106",
X"9438811f",
X"7081ff06",
X"811e7081",
X"ff065f52",
X"405386dc",
X"39748c2e",
X"09810686",
X"d338ff1f",
X"7081ff06",
X"ff1e7081",
X"ff065f52",
X"40537b63",
X"2586bd38",
X"ff4386b8",
X"3976812e",
X"83bb3876",
X"81248938",
X"76802e8d",
X"3886a539",
X"76822e84",
X"a638869c",
X"39f81553",
X"72842684",
X"95387284",
X"2981d7cc",
X"05537208",
X"0464802e",
X"80cd3878",
X"22838080",
X"06537283",
X"80802e09",
X"8106bc38",
X"80567564",
X"27a43875",
X"1e7083ff",
X"ff067710",
X"1b901172",
X"832a5851",
X"57515373",
X"75347287",
X"0681712b",
X"51537281",
X"16348116",
X"7081ff06",
X"57539776",
X"27cc387f",
X"84074080",
X"0b993d43",
X"56611670",
X"3370982b",
X"70982c51",
X"51515380",
X"732480fb",
X"38607329",
X"1e7083ff",
X"ff067a22",
X"83808006",
X"52585372",
X"8380802e",
X"09810680",
X"de386088",
X"32703070",
X"72078025",
X"63903270",
X"30707207",
X"80257307",
X"53545851",
X"55537380",
X"2ebd3876",
X"87065372",
X"b6387584",
X"29761005",
X"79118411",
X"79832a57",
X"57515373",
X"75346081",
X"16346586",
X"14236688",
X"14237587",
X"387f8107",
X"408d3975",
X"812e0981",
X"0685387f",
X"82074081",
X"167081ff",
X"06575381",
X"7627fee5",
X"38636129",
X"1e7083ff",
X"ff065f53",
X"80704642",
X"ff028405",
X"80dd0534",
X"ff0b993d",
X"3483f539",
X"811c7081",
X"ff065d53",
X"80427381",
X"2e098106",
X"8e387781",
X"800a2981",
X"800a0558",
X"80d33973",
X"802e8938",
X"73822e09",
X"81068d38",
X"7c81800a",
X"2981800a",
X"055da439",
X"815f83b8",
X"39ff1c70",
X"81ff065d",
X"537b6325",
X"8338ff43",
X"7c802e92",
X"387c8180",
X"0a2981ff",
X"0a055d7c",
X"982c5d83",
X"93397780",
X"2e923877",
X"81800a29",
X"81ff0a05",
X"5877982c",
X"5882fd39",
X"7753839e",
X"39748926",
X"80f43874",
X"842981d7",
X"e0055372",
X"08047387",
X"2e82e138",
X"73852e82",
X"db387388",
X"2e82d538",
X"738c2e82",
X"cf387389",
X"2e098106",
X"86388145",
X"82c23973",
X"812e0981",
X"0682b938",
X"62802582",
X"b3387b98",
X"2b70982c",
X"514382a8",
X"397383ff",
X"ff064682",
X"9f397383",
X"ffff0647",
X"82963973",
X"81ff0641",
X"828e3973",
X"811a3482",
X"87397381",
X"ff064481",
X"ff397e53",
X"82a03974",
X"812e81e3",
X"38748124",
X"89387480",
X"2e8d3881",
X"e7397482",
X"2e81d838",
X"81de3974",
X"567b8338",
X"81567453",
X"73862e09",
X"81069738",
X"75810653",
X"72802e8e",
X"38782282",
X"ffff06fe",
X"80800753",
X"b6397b83",
X"38815373",
X"822e0981",
X"06973872",
X"81065372",
X"802e8e38",
X"782281ff",
X"ff068180",
X"80075393",
X"397b9638",
X"fc145372",
X"81268e38",
X"7822ff80",
X"80075372",
X"792380e5",
X"39805573",
X"812e0981",
X"06833873",
X"55775377",
X"802e8938",
X"74810653",
X"7280ca38",
X"72d01554",
X"55728126",
X"83388155",
X"77802eb9",
X"38748106",
X"5372802e",
X"b0387822",
X"83808006",
X"53728380",
X"802e0981",
X"069f3873",
X"b02e0981",
X"06873861",
X"993d3491",
X"3973b12e",
X"09810689",
X"38610284",
X"0580dd05",
X"34618105",
X"538c3961",
X"74318105",
X"53843961",
X"14537283",
X"ffff0642",
X"79f7fb38",
X"7d832a53",
X"72821a34",
X"78228380",
X"80065372",
X"8380802e",
X"09810688",
X"3881537f",
X"872e8338",
X"80537283",
X"c0800c99",
X"3d0d04fd",
X"3d0d7583",
X"11338212",
X"3371982b",
X"71902b07",
X"81143370",
X"882b7207",
X"75337107",
X"83c0800c",
X"52535456",
X"5452853d",
X"0d04f63d",
X"0d02b705",
X"33028405",
X"bb053302",
X"8805bf05",
X"335b5b5b",
X"80588057",
X"78882b7a",
X"07568055",
X"7a548153",
X"a3527c51",
X"92cc3f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f63d",
X"0d02b705",
X"33028405",
X"bb053302",
X"8805bf05",
X"335b5b5b",
X"80588057",
X"78882b7a",
X"07568055",
X"7a548353",
X"a3527c51",
X"92903f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f73d",
X"0d02b305",
X"33028405",
X"b6052260",
X"5a585680",
X"55805480",
X"5381a352",
X"7b5191e2",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8b3d0d04",
X"ee3d0d64",
X"90115c5c",
X"807b3480",
X"0b841c0c",
X"800b881c",
X"34810b89",
X"1c34880b",
X"8a1c3480",
X"0b8b1c34",
X"881b08c1",
X"06810788",
X"1c0c8f3d",
X"70545d88",
X"527b519b",
X"eb3f83c0",
X"800881ff",
X"06705b59",
X"7881a938",
X"903d335e",
X"81db5a7d",
X"892e0981",
X"06819938",
X"7c539252",
X"7b519bc4",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"8182387c",
X"58885778",
X"56a95578",
X"54865381",
X"a0527b51",
X"90d03f83",
X"c0800881",
X"ff06705b",
X"597880e0",
X"3802ba05",
X"337b347c",
X"5478537d",
X"527b519b",
X"ac3f83c0",
X"800881ff",
X"06705b59",
X"7880c138",
X"02bd0533",
X"527b519b",
X"c43f83c0",
X"800881ff",
X"06705b59",
X"78aa3881",
X"7b335a5a",
X"79792699",
X"38805479",
X"5388527b",
X"51fdbb3f",
X"811a7081",
X"ff067c33",
X"525b59e4",
X"39810b88",
X"1c34805a",
X"7983c080",
X"0c943d0d",
X"04800b83",
X"c0800c04",
X"f93d0d79",
X"028405ab",
X"05338e3d",
X"70545858",
X"58ffbeb0",
X"3f8a3d8a",
X"0551ffbe",
X"a73f7551",
X"fc8d3f83",
X"c0800884",
X"86812ebe",
X"3883c080",
X"08848681",
X"26993883",
X"c0800884",
X"82802e80",
X"e63883c0",
X"80088482",
X"812e9f38",
X"81b43983",
X"c0800880",
X"c082832e",
X"80f43883",
X"c0800880",
X"c086832e",
X"80e83881",
X"993983c0",
X"9c335580",
X"5674762e",
X"09810681",
X"8b387454",
X"76539152",
X"7751fbd6",
X"3f745476",
X"53905277",
X"51fbcb3f",
X"74547653",
X"84527751",
X"fbfc3f81",
X"0b83c09c",
X"3481b156",
X"80de3980",
X"54765391",
X"527751fb",
X"a93f8054",
X"76539052",
X"7751fb9e",
X"3f800b83",
X"c09c3476",
X"52871833",
X"5197963f",
X"b5398054",
X"76539452",
X"7751fb82",
X"3f805476",
X"53905277",
X"51faf73f",
X"7551ffbc",
X"db3f83c0",
X"8008892a",
X"81065376",
X"52871833",
X"5190cd3f",
X"800b83c0",
X"9c348056",
X"7583c080",
X"0c893d0d",
X"04f23d0d",
X"6090115a",
X"58800b88",
X"1a337159",
X"56567476",
X"2e82a538",
X"82ac3f84",
X"190883c0",
X"80082682",
X"95387833",
X"5a810b8e",
X"3d23903d",
X"f81155f4",
X"05539918",
X"5277518a",
X"e53f83c0",
X"800881ff",
X"06705755",
X"74772e09",
X"810681d9",
X"38863974",
X"5681d239",
X"81568257",
X"8e3d3377",
X"06557480",
X"2ebb3880",
X"0b8d3d34",
X"903df005",
X"54845375",
X"527751fa",
X"cd3f83c0",
X"800881ff",
X"0655749d",
X"387b5375",
X"527751fc",
X"e73f83c0",
X"800881ff",
X"06557481",
X"b12e818b",
X"3874ffb3",
X"38761081",
X"fc068117",
X"7081ff06",
X"58565787",
X"7627ffa8",
X"38815675",
X"7a2680eb",
X"38800b8d",
X"3d348c3d",
X"70555784",
X"53755277",
X"51f9f73f",
X"83c08008",
X"81ff0655",
X"7480c138",
X"7651ffba",
X"d73f83c0",
X"80088287",
X"06557482",
X"812e0981",
X"06aa3802",
X"ae053381",
X"07557402",
X"8405ae05",
X"347b5375",
X"527751fb",
X"eb3f83c0",
X"800881ff",
X"06557481",
X"b12e9038",
X"74feb838",
X"81167081",
X"ff065755",
X"ff913980",
X"567581ff",
X"0656973f",
X"83c08008",
X"8fd00584",
X"1a0c7557",
X"7683c080",
X"0c903d0d",
X"04049080",
X"a00883c0",
X"800c04ff",
X"3d0d7387",
X"e82951ff",
X"91d63f83",
X"3d0d0404",
X"83caf80b",
X"83c0800c",
X"04fd3d0d",
X"75775454",
X"800b83ca",
X"d834728a",
X"38909080",
X"0b84150c",
X"90397281",
X"2e098106",
X"88389098",
X"800b8415",
X"0c841408",
X"83caf00c",
X"800b8815",
X"0c800b8c",
X"150c83ca",
X"f0085382",
X"0b878014",
X"348151ff",
X"9e3f83ca",
X"f0085380",
X"0b881434",
X"83caf008",
X"53810b87",
X"80143483",
X"caf00853",
X"800b8c14",
X"3483caf0",
X"0853800b",
X"a4143491",
X"7434800b",
X"83c0a034",
X"800b83c0",
X"a434800b",
X"83c0a834",
X"80547381",
X"c42983ca",
X"fc055380",
X"0b831434",
X"81147081",
X"ff065553",
X"8f7427e6",
X"38853d0d",
X"04fe3d0d",
X"74768211",
X"3370bf06",
X"81712bff",
X"05565151",
X"52539071",
X"278338ff",
X"52765171",
X"712383ca",
X"f0085187",
X"13339012",
X"34800b83",
X"c0a43480",
X"0b83c0a8",
X"34881333",
X"8a143352",
X"5271802e",
X"aa387081",
X"ff065184",
X"52708338",
X"70527183",
X"c0a4348a",
X"13337030",
X"70802584",
X"2b708807",
X"51515253",
X"7083c0a8",
X"34903970",
X"81ff0651",
X"70833898",
X"527183c0",
X"a834800b",
X"83c0800c",
X"843d0d04",
X"f13d0d61",
X"6568028c",
X"0580cb05",
X"33029005",
X"80ce0522",
X"02940580",
X"d6052242",
X"40415a40",
X"40fd8b3f",
X"83c08008",
X"a788055b",
X"8070715b",
X"5b528394",
X"3983caf0",
X"08517d94",
X"123483c0",
X"a4338107",
X"55807054",
X"567f8626",
X"80ea387f",
X"842981d8",
X"940583ca",
X"f0085351",
X"70080480",
X"0b841334",
X"a1397733",
X"70307080",
X"25837131",
X"51515253",
X"70841334",
X"8d39810b",
X"841334b8",
X"39830b84",
X"13348170",
X"5456ad39",
X"810b8413",
X"34a23977",
X"33703070",
X"80258371",
X"31515152",
X"53708413",
X"34807833",
X"52527083",
X"38815271",
X"78348153",
X"74880755",
X"83c0a833",
X"83caf008",
X"5257810b",
X"81d01234",
X"83caf008",
X"51810b81",
X"9012347e",
X"802eae38",
X"72802ea9",
X"387eff1e",
X"52547083",
X"ffff0653",
X"7283ffff",
X"2e973873",
X"70810555",
X"3383caf0",
X"08535170",
X"81c01334",
X"ff1351de",
X"3983caf0",
X"08a81133",
X"53517688",
X"123483ca",
X"f0085174",
X"713481ff",
X"52913983",
X"caf008a0",
X"11337081",
X"06515253",
X"708f38fa",
X"fd3f7a83",
X"c0800826",
X"e6388188",
X"39810ba0",
X"143483ca",
X"f008a811",
X"3380ff06",
X"70780752",
X"53517080",
X"2e80ed38",
X"71862a70",
X"81065151",
X"70802e91",
X"38807833",
X"52537083",
X"38815372",
X"783480e0",
X"3971842a",
X"70810651",
X"5170802e",
X"9b388119",
X"7083ffff",
X"067d3070",
X"9f2a5152",
X"5a51787c",
X"2e098106",
X"af38a439",
X"71832a70",
X"81065151",
X"70802e93",
X"38811a70",
X"81ff065b",
X"5179832e",
X"09810690",
X"388a3971",
X"a3065170",
X"802e8538",
X"71519239",
X"f9e43f7a",
X"83c08008",
X"26fce238",
X"7181bf06",
X"517083c0",
X"800c913d",
X"0d04f63d",
X"0d02b305",
X"33028405",
X"b7053302",
X"8805ba05",
X"22595959",
X"800b8c3d",
X"348c3dfc",
X"05568055",
X"80547653",
X"77527851",
X"fbf23f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f33d",
X"0d7f6264",
X"028c0580",
X"c2052272",
X"22811533",
X"425f415e",
X"59598078",
X"237d5378",
X"33528151",
X"ffa03f83",
X"c0800881",
X"ff065675",
X"802e8638",
X"755481ad",
X"3983caf0",
X"08a81133",
X"821b3370",
X"862a7081",
X"0673982b",
X"5351575c",
X"56577980",
X"25833881",
X"5673762e",
X"873881f0",
X"54818239",
X"818c1733",
X"7081ff06",
X"79227d71",
X"31902b70",
X"902c7009",
X"709f2c72",
X"06705252",
X"53515357",
X"57547574",
X"24833875",
X"55748480",
X"8029fc80",
X"80057090",
X"2c515574",
X"ff2e9438",
X"83caf008",
X"81801133",
X"5154737c",
X"7081055e",
X"34db3977",
X"22760554",
X"73782379",
X"09709f2a",
X"70810682",
X"1c3381bf",
X"0671862b",
X"07515151",
X"5473821a",
X"347c7626",
X"8a387722",
X"547a7426",
X"febb3880",
X"547383c0",
X"800c8f3d",
X"0d04f93d",
X"0d7a5780",
X"0b893d23",
X"893dfc05",
X"53765279",
X"51f8da3f",
X"83c08008",
X"81ff0670",
X"57557496",
X"387c547b",
X"53883d22",
X"527651fd",
X"e53f83c0",
X"800881ff",
X"06567583",
X"c0800c89",
X"3d0d04f0",
X"3d0d6266",
X"02880580",
X"ce052241",
X"5d5e8002",
X"840580d2",
X"05227f81",
X"0533ff11",
X"5a5d5a5d",
X"81da5876",
X"bf2680e9",
X"3878802e",
X"80e1387a",
X"58787b27",
X"83387858",
X"821e3370",
X"872a585a",
X"76923d34",
X"923dfc05",
X"5677557b",
X"547e537d",
X"33528251",
X"f8de3f83",
X"c0800881",
X"ff065d80",
X"0b923d33",
X"585a7680",
X"2e833881",
X"5a821e33",
X"80ff067a",
X"872b0757",
X"76821f34",
X"7c913878",
X"78317083",
X"ffff0679",
X"1e5e5a57",
X"ff9b397c",
X"587783c0",
X"800c923d",
X"0d04f83d",
X"0d7b0284",
X"05b20522",
X"5858800b",
X"8a3d238a",
X"3dfc0553",
X"77527a51",
X"f6f73f83",
X"c0800881",
X"ff067057",
X"55749638",
X"7d547653",
X"893d2252",
X"7751feaf",
X"3f83c080",
X"0881ff06",
X"567583c0",
X"800c8a3d",
X"0d04ec3d",
X"0d666e02",
X"880580df",
X"0533028c",
X"0580e305",
X"33029005",
X"80e70533",
X"02940580",
X"eb053302",
X"980580ee",
X"05224143",
X"415f5c40",
X"570280f2",
X"0522963d",
X"23963df0",
X"05538417",
X"70537752",
X"59f6863f",
X"83c08008",
X"81ff0658",
X"7781e538",
X"777a8180",
X"06584080",
X"77258338",
X"81407994",
X"3d347b02",
X"840580c9",
X"05347c02",
X"840580ca",
X"05347d02",
X"840580cb",
X"05347a95",
X"3d347a88",
X"2a577602",
X"840580cd",
X"0534953d",
X"22577602",
X"840580ce",
X"05347688",
X"2a577602",
X"840580cf",
X"05347792",
X"3d34963d",
X"ec115757",
X"8855f417",
X"54923d22",
X"53775277",
X"51f6953f",
X"83c08008",
X"81ff0658",
X"7780ed38",
X"7e802e80",
X"cb38923d",
X"22790858",
X"587f802e",
X"9c387681",
X"80800779",
X"0c7e5496",
X"3dfc0553",
X"7783ffff",
X"06527851",
X"f9fc3f99",
X"39768280",
X"8007790c",
X"7e54953d",
X"22537783",
X"ffff0652",
X"7851fc8f",
X"3f83c080",
X"0881ff06",
X"58779d38",
X"923d2253",
X"80527f30",
X"70802584",
X"71315351",
X"57f9873f",
X"83c08008",
X"81ff0658",
X"7783c080",
X"0c963d0d",
X"04f63d0d",
X"7c028405",
X"b705335b",
X"5b805880",
X"57805680",
X"55795485",
X"5380527a",
X"51fda33f",
X"83c08008",
X"81ff0659",
X"78853879",
X"871c3478",
X"83c0800c",
X"8c3d0d04",
X"f93d0d02",
X"a7053302",
X"8405ab05",
X"33028805",
X"af053358",
X"5957800b",
X"83caff33",
X"54547274",
X"2e9f3881",
X"147081ff",
X"06555373",
X"8f2681b6",
X"387381c4",
X"2983cafc",
X"05831133",
X"515372e3",
X"387381c4",
X"2983caf8",
X"0555800b",
X"87163476",
X"88163475",
X"8a163477",
X"89163480",
X"750c83ca",
X"f0088c16",
X"0c800b84",
X"1634880b",
X"85163480",
X"0b861634",
X"841508ff",
X"a1ff06a0",
X"80078416",
X"0c811470",
X"81ff0653",
X"537451fe",
X"bc3f83c0",
X"800881ff",
X"06705553",
X"7280cd38",
X"8a397308",
X"750c7254",
X"80c23972",
X"81ddb055",
X"5681ddb0",
X"08802eb2",
X"38758429",
X"14700876",
X"53700851",
X"5454722d",
X"83c08008",
X"81ff0653",
X"72802ece",
X"38811670",
X"81ff0681",
X"ddb07184",
X"29115356",
X"57537208",
X"d0388054",
X"7383c080",
X"0c893d0d",
X"04f93d0d",
X"7957800b",
X"84180883",
X"caf00c58",
X"f0883f88",
X"170883c0",
X"80082783",
X"ed38effa",
X"3f83c080",
X"08810588",
X"180c83ca",
X"f008b811",
X"337081ff",
X"06515154",
X"73812ea4",
X"38738124",
X"88387378",
X"2e8a38b8",
X"3973822e",
X"9538b139",
X"763381f0",
X"06547390",
X"2ea63891",
X"7734a139",
X"73587633",
X"81f00654",
X"73902e09",
X"81069138",
X"efa83f83",
X"c0800881",
X"c8058c18",
X"0ca07734",
X"80567581",
X"c42983ca",
X"ff113355",
X"5573802e",
X"aa3883ca",
X"f8157008",
X"56547480",
X"2e9d3888",
X"1508802e",
X"96388c14",
X"0883caf0",
X"082e0981",
X"06893873",
X"51881508",
X"54732d81",
X"167081ff",
X"0657548f",
X"7627ffba",
X"38763354",
X"73b02e81",
X"993873b0",
X"248f3873",
X"912eab38",
X"73a02e80",
X"f53882a6",
X"397380d0",
X"2e81e438",
X"7380d024",
X"8b387380",
X"c02e8199",
X"38828f39",
X"7381802e",
X"81fb3882",
X"85398056",
X"7581c429",
X"83cafc11",
X"83113356",
X"59557380",
X"2ea83883",
X"caf81570",
X"08565474",
X"802e9b38",
X"8c140883",
X"caf0082e",
X"0981068e",
X"38735184",
X"15085473",
X"2d800b83",
X"19348116",
X"7081ff06",
X"57548f76",
X"27ffb938",
X"92773481",
X"b539edc2",
X"3f8c1708",
X"83c08008",
X"2781a738",
X"b0773481",
X"a13983ca",
X"f0085480",
X"0b8c1534",
X"83caf008",
X"54840b88",
X"153480c0",
X"7734ed96",
X"3f83c080",
X"08b2058c",
X"180c80fa",
X"39ed873f",
X"8c170883",
X"c0800827",
X"80ec3883",
X"caf00854",
X"810b8c15",
X"3483caf0",
X"0854800b",
X"88153483",
X"caf00854",
X"880ba015",
X"34ecdb3f",
X"83c08008",
X"94058c18",
X"0c80d077",
X"34bc3983",
X"caf008a0",
X"11337083",
X"2a708106",
X"51515555",
X"73802ea6",
X"38880ba0",
X"1634ecae",
X"3f8c1708",
X"83c08008",
X"279438ff",
X"8077348e",
X"39775380",
X"528051fa",
X"8b3fff90",
X"773483ca",
X"f008a011",
X"3370832a",
X"70810651",
X"51555573",
X"802e8638",
X"880ba016",
X"34893d0d",
X"04f63d0d",
X"02b30533",
X"028405b7",
X"05335b5b",
X"800b83ca",
X"fc708412",
X"72745d59",
X"575b5856",
X"83153353",
X"72802e80",
X"f3387333",
X"537a732e",
X"09810680",
X"e7388114",
X"33537973",
X"2e098106",
X"80da3880",
X"557481c4",
X"2983cb80",
X"05703383",
X"1b335855",
X"5373762e",
X"0981068a",
X"38811333",
X"527351ff",
X"9c3f8115",
X"7081ff06",
X"56538f75",
X"27d33880",
X"0b83caf8",
X"19700856",
X"54557375",
X"2e913872",
X"51841408",
X"53722d83",
X"c0800881",
X"ff065580",
X"0b831834",
X"7453a039",
X"811681c4",
X"1981c417",
X"81c41781",
X"c41d81c4",
X"1c5c5d57",
X"5759568f",
X"7625fee8",
X"38805372",
X"83c0800c",
X"8c3d0d04",
X"f83d0d02",
X"ae05227d",
X"59578056",
X"81558054",
X"86538180",
X"527a51f5",
X"953f83c0",
X"800881ff",
X"0683c080",
X"0c8a3d0d",
X"04f73d0d",
X"02b20522",
X"028405b7",
X"0533605a",
X"5b578056",
X"82557954",
X"86538180",
X"527b51f4",
X"e53f83c0",
X"800881ff",
X"0683c080",
X"0c8b3d0d",
X"04f83d0d",
X"02af0533",
X"59805880",
X"57805680",
X"55785489",
X"5380527a",
X"51f4bb3f",
X"83c08008",
X"81ff0683",
X"c0800c8a",
X"3d0d0400",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002b0a",
X"00002b4b",
X"00002b6d",
X"00002b93",
X"00002b93",
X"00002b93",
X"00002b93",
X"00002c04",
X"00002c55",
X"00004170",
X"000049b4",
X"00004a6d",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3f00",
X"0c0c4000",
X"0a0a4100",
X"0b0b4100",
X"07074100",
X"0a0b4300",
X"080b4200",
X"04044500",
X"05054400",
X"06060004",
X"08080004",
X"09090004",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"000056f9",
X"00005a00",
X"0000580c",
X"00005a00",
X"00005849",
X"0000589a",
X"000058d9",
X"000058e2",
X"00005a00",
X"00005a00",
X"00005a00",
X"00005a00",
X"000058eb",
X"000058f3",
X"000058fa",
X"00005b00",
X"00005bf9",
X"00005d0d",
X"00006003",
X"0000601e",
X"0000600a",
X"0000601e",
X"00006025",
X"00006030",
X"00006037",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"66726565",
X"7a65722e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00006c70",
X"00006c74",
X"00006c7c",
X"00006c88",
X"00006c94",
X"00006ca0",
X"00006cac",
X"00006cb0",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00006c08",
X"00006a5c",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"69383030",
X"00000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
