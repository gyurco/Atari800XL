
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f3",
X"c0738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80f7",
X"800c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f1",
X"802d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580f0bf",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80dbcb04",
X"fd3d0d75",
X"705254ae",
X"a63f83e0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83e0",
X"8008732e",
X"a13883e0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183e0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83e2c008",
X"248a38b4",
X"f73fff0b",
X"83e2c00c",
X"800b83e0",
X"800c04ff",
X"3d0d7352",
X"83e09c08",
X"722e8d38",
X"d93f7151",
X"96993f71",
X"83e09c0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"558154bc",
X"15088191",
X"387451cf",
X"3f795880",
X"7a2580f7",
X"3883e2f0",
X"0870892a",
X"5783ff06",
X"78848072",
X"31565657",
X"73782583",
X"38735575",
X"83e2c008",
X"2e8438ff",
X"893f83e2",
X"c0088025",
X"a6387589",
X"2b5198dc",
X"3f83e2f0",
X"088f3dfc",
X"11555c54",
X"8152f81b",
X"5196c63f",
X"761483e2",
X"f00c7583",
X"e2c00c74",
X"53765278",
X"51b3a83f",
X"83e08008",
X"83e2f008",
X"1683e2f0",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8b3861",
X"7a710c54",
X"75547580",
X"2e833881",
X"547383e0",
X"800c8e3d",
X"0d04fc3d",
X"0dfe9b3f",
X"7651feaf",
X"3f863dfc",
X"05537852",
X"775195e9",
X"3f797571",
X"0c5483e0",
X"80085483",
X"e0800880",
X"2e833881",
X"547383e0",
X"800c863d",
X"0d04fe3d",
X"0d7583e2",
X"c0085353",
X"80722489",
X"3871732e",
X"8438fdd6",
X"3f7451fd",
X"ea3f7251",
X"97ae3f83",
X"e0800852",
X"83e08008",
X"802e8338",
X"81527183",
X"e0800c84",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"e0800c51",
X"823d0d04",
X"80c40b83",
X"e0800c04",
X"fd3d0d75",
X"77715470",
X"535553a9",
X"fe3f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfceb3f",
X"735193ab",
X"3f7383e0",
X"9c0c83e0",
X"80085383",
X"e0800880",
X"2e833881",
X"537283e0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcbf3f",
X"72802ea5",
X"38bc1308",
X"527351a9",
X"883f83e0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"e0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83e0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83e2c0",
X"0c7483e0",
X"a00c7583",
X"e2bc0caf",
X"dc3f83e0",
X"800881ff",
X"06528153",
X"71993883",
X"e2d8518e",
X"943f83e0",
X"80085283",
X"e0800880",
X"2e833872",
X"52715372",
X"83e0800c",
X"843d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"51a6f93f",
X"83e08008",
X"557483e0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"e0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283e2bc",
X"085180df",
X"c23f83e0",
X"800857f9",
X"e13f7952",
X"83e2c451",
X"95b73f83",
X"e0800854",
X"805383e0",
X"8008732e",
X"09810682",
X"833883e0",
X"a0080b0b",
X"80f4f453",
X"705256a6",
X"b63f0b0b",
X"80f4f452",
X"80c01651",
X"a6a93f75",
X"bc170c73",
X"82c0170c",
X"810b82c4",
X"170c810b",
X"82c8170c",
X"7382cc17",
X"0cff1782",
X"d0175557",
X"81913983",
X"e0ac3370",
X"822a7081",
X"06515455",
X"72818038",
X"74812a81",
X"06587780",
X"f6387484",
X"2a810682",
X"c4150c83",
X"e0ac3381",
X"0682c815",
X"0c795273",
X"51a5d03f",
X"7351a5e7",
X"3f83e080",
X"081453af",
X"73708105",
X"553472bc",
X"150c83e0",
X"ad527251",
X"a5b13f83",
X"e0a40882",
X"c0150c83",
X"e0ba5280",
X"c01451a5",
X"9e3f7880",
X"2e8d3873",
X"51782d83",
X"e0800880",
X"2e993877",
X"82cc150c",
X"75802e86",
X"387382cc",
X"170c7382",
X"d015ff19",
X"59555676",
X"802e9b38",
X"83e0a452",
X"83e2c451",
X"94ad3f83",
X"e080088a",
X"3883e0ad",
X"335372fe",
X"d2387880",
X"2e893883",
X"e0a00851",
X"fcb83f83",
X"e0a00853",
X"7283e080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb53f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f690",
X"3f83e080",
X"08745387",
X"3d705355",
X"55f6b03f",
X"f7903f73",
X"51d33f63",
X"53745283",
X"e0800851",
X"fab83f92",
X"3d0d0471",
X"83e0800c",
X"0480c012",
X"83e0800c",
X"04803d0d",
X"7282c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"e0800c51",
X"823d0d04",
X"f93d0d79",
X"83e09008",
X"57578177",
X"27819638",
X"76881708",
X"27818e38",
X"75335574",
X"822e8938",
X"74832eb3",
X"3880fe39",
X"74547610",
X"83fe0653",
X"76882a8c",
X"17080552",
X"893dfc05",
X"51aa8a3f",
X"83e08008",
X"80df3802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d13984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"51a9da3f",
X"83e08008",
X"b038029f",
X"05330284",
X"059e0533",
X"71982b71",
X"902b0702",
X"8c059d05",
X"3370882b",
X"72078d3d",
X"337180ff",
X"fffe8006",
X"07515253",
X"57585683",
X"39815574",
X"83e0800c",
X"893d0d04",
X"fb3d0d83",
X"e09008fe",
X"19881208",
X"fe055556",
X"54805674",
X"73278d38",
X"82143375",
X"71299416",
X"08055753",
X"7583e080",
X"0c873d0d",
X"04fc3d0d",
X"7652800b",
X"83e09008",
X"70335152",
X"5370832e",
X"09810691",
X"38951233",
X"94133371",
X"982b7190",
X"2b075555",
X"519b1233",
X"9a133371",
X"882b0774",
X"0783e080",
X"0c55863d",
X"0d04fc3d",
X"0d7683e0",
X"90085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"fed63f83",
X"e0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183e080",
X"0c863d0d",
X"04fa3d0d",
X"7883e090",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fcb13f",
X"81527183",
X"e0800827",
X"a8388352",
X"83e08008",
X"88170827",
X"9c3883e0",
X"80088c16",
X"0c83e080",
X"0851fdbc",
X"3f83e080",
X"0890160c",
X"73752380",
X"527183e0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585e5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"9f269138",
X"7a51fdd2",
X"3f83e080",
X"0856807d",
X"34838139",
X"933d841c",
X"08705859",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"3880705a",
X"5c887f08",
X"5f5a7b81",
X"1d7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535e57",
X"557480e7",
X"3876ae2e",
X"09810683",
X"38815578",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675bb",
X"3888598b",
X"5affab39",
X"76982b55",
X"74802587",
X"3880f2d0",
X"173357ff",
X"9f175574",
X"99268938",
X"e0177081",
X"ff065855",
X"78811a70",
X"81ff0672",
X"1b535b57",
X"55767534",
X"fef8397b",
X"1e7f0c80",
X"5576a026",
X"83388155",
X"748b1934",
X"7a51fc82",
X"3f83e080",
X"0880f538",
X"a0547a22",
X"70852b83",
X"e0065455",
X"901b0852",
X"7c51a495",
X"3f83e080",
X"085783e0",
X"80088181",
X"387c3355",
X"74802e80",
X"f4388b1d",
X"3370832a",
X"70810651",
X"565674b4",
X"388b7d84",
X"1d0883e0",
X"8008595b",
X"5b58ff18",
X"5877ff2e",
X"9a387970",
X"81055b33",
X"79708105",
X"5b337171",
X"31525656",
X"75802ee2",
X"38863975",
X"802e9638",
X"7a51fbe5",
X"3fff8639",
X"83e08008",
X"5683e080",
X"08b63883",
X"39765684",
X"1b088b11",
X"33515574",
X"a7388b1d",
X"3370842a",
X"70810651",
X"56567489",
X"38835694",
X"39815690",
X"397c51fa",
X"943f83e0",
X"8008881c",
X"0cfd8139",
X"7583e080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"51a2da3f",
X"835683e0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"51a2ae3f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"7651a285",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583e080",
X"0c8a3d0d",
X"04eb3d0d",
X"675a800b",
X"83e0900c",
X"a1a73f83",
X"e0800881",
X"06558256",
X"7483ef38",
X"7475538f",
X"3d705357",
X"59feca3f",
X"83e08008",
X"81ff0657",
X"76812e09",
X"810680d4",
X"38905483",
X"be537452",
X"7551a199",
X"3f83e080",
X"0880c938",
X"8f3d3355",
X"74802e80",
X"c93802bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"33710770",
X"587b575e",
X"525e5759",
X"57fdee3f",
X"83e08008",
X"81ff0657",
X"76832e09",
X"81068638",
X"815682f2",
X"3976802e",
X"86388656",
X"82e839a4",
X"548d5378",
X"527551a0",
X"b03f8156",
X"83e08008",
X"82d43802",
X"be053302",
X"8405bd05",
X"3371882b",
X"07595d77",
X"ab380280",
X"ce053302",
X"840580cd",
X"05337198",
X"2b71902b",
X"07973d33",
X"70882b72",
X"07029405",
X"80cb0533",
X"71075452",
X"5e575956",
X"02b70533",
X"78712902",
X"8805b605",
X"33028c05",
X"b5053371",
X"882b0770",
X"1d707f8c",
X"050c5f59",
X"57595d8e",
X"3d33821b",
X"3402b905",
X"33903d33",
X"71882b07",
X"5a5c7884",
X"1b2302bb",
X"05330284",
X"05ba0533",
X"71882b07",
X"565c74ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"07515253",
X"575e5c74",
X"76317831",
X"79842a90",
X"3d335471",
X"71315356",
X"5680d0a7",
X"3f83e080",
X"08820570",
X"881c0c83",
X"e08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83e0900c",
X"80567583",
X"e0800c97",
X"3d0d04e9",
X"3d0d83e0",
X"90085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e53f83e0",
X"80085483",
X"e0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f489",
X"3f83e080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383e080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83e09008",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0e93f",
X"83e08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"833f83e0",
X"80085583",
X"e0800880",
X"2eff8938",
X"83e08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"519ad63f",
X"83e08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83e0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83e09008",
X"55568555",
X"73802e81",
X"e3388114",
X"33810653",
X"84557280",
X"2e81d538",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b9388214",
X"3370892b",
X"56537680",
X"2eb73874",
X"52ff1651",
X"80cba83f",
X"83e08008",
X"ff187654",
X"70535853",
X"80cb983f",
X"83e08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed63f83",
X"e0800853",
X"810b83e0",
X"8008278b",
X"38881408",
X"83e08008",
X"26883880",
X"0b811534",
X"b03983e0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc53f",
X"83e08008",
X"8c3883e0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683e0",
X"800805a8",
X"150c8055",
X"7483e080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83e09008",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1cf3f",
X"83e08008",
X"5583e080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef5",
X"3f83e080",
X"0888170c",
X"7551efa6",
X"3f83e080",
X"08557483",
X"e0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683e0",
X"9008802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f53f83e0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"96df3f83",
X"e0800841",
X"83e08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"eddf3f83",
X"e0800841",
X"83e08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"8e853f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f03f83e0",
X"80088332",
X"70307072",
X"079f2c83",
X"e0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"8c913f75",
X"83e0800c",
X"9e3d0d04",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"7751e0d2",
X"3f83e080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3380f788",
X"0b80f788",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"527751e0",
X"813f83e0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583e0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"558b983f",
X"83e08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"8114518a",
X"b03f83e0",
X"80083070",
X"83e08008",
X"07802583",
X"e0800c53",
X"863d0d04",
X"fc3d0d76",
X"705255e6",
X"ee3f83e0",
X"80085481",
X"5383e080",
X"0880c138",
X"7451e6b1",
X"3f83e080",
X"0880f584",
X"5383e080",
X"085253ff",
X"913f83e0",
X"8008a138",
X"80f58852",
X"7251ff82",
X"3f83e080",
X"08923880",
X"f58c5272",
X"51fef33f",
X"83e08008",
X"802e8338",
X"81547353",
X"7283e080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"e68d3f81",
X"5383e080",
X"08983873",
X"51e5d63f",
X"83e38808",
X"5283e080",
X"0851feba",
X"3f83e080",
X"08537283",
X"e0800c85",
X"3d0d04df",
X"3d0da43d",
X"0870525e",
X"dbfb3f83",
X"e0800833",
X"953d5654",
X"73963880",
X"fa845274",
X"5189903f",
X"9a397d52",
X"7851defc",
X"3f84cf39",
X"7d51dbe1",
X"3f83e080",
X"08527451",
X"db913f80",
X"43804280",
X"41804083",
X"e3900852",
X"943d7052",
X"5de1e43f",
X"83e08008",
X"59800b83",
X"e0800855",
X"5b83e080",
X"087b2e94",
X"38811b74",
X"525be4e6",
X"3f83e080",
X"085483e0",
X"8008ee38",
X"805aff5f",
X"7909709f",
X"2c7b065b",
X"547a7a24",
X"8438ff1b",
X"5af61a70",
X"09709f2c",
X"72067bff",
X"125a5a52",
X"55558075",
X"25953876",
X"51e4ab3f",
X"83e08008",
X"76ff1858",
X"55577380",
X"24ed3874",
X"7f2e8638",
X"a0d83f74",
X"5f78ff1b",
X"70585d58",
X"807a2595",
X"387751e4",
X"813f83e0",
X"800876ff",
X"18585558",
X"738024ed",
X"38800b83",
X"e7c00c80",
X"0b83e7e4",
X"0c80f590",
X"518d8f3f",
X"81800b83",
X"e7e40c80",
X"f598518d",
X"813fa80b",
X"83e7c00c",
X"76802e80",
X"e43883e7",
X"c0087779",
X"32703070",
X"72078025",
X"70872b83",
X"e7e40c51",
X"56785356",
X"56e3b83f",
X"83e08008",
X"802e8838",
X"80f5a051",
X"8cc83f76",
X"51e2fa3f",
X"83e08008",
X"5280f6ac",
X"518cb73f",
X"7651e382",
X"3f83e080",
X"0883e7c0",
X"08555775",
X"74258638",
X"a81656f7",
X"397583e7",
X"c00c86f0",
X"7624ff98",
X"3887980b",
X"83e7c00c",
X"77802eb1",
X"387751e2",
X"b83f83e0",
X"80087852",
X"55e2d83f",
X"80f5a854",
X"83e08008",
X"8d388739",
X"80763481",
X"d03980f5",
X"a4547453",
X"735280f4",
X"f8518bd6",
X"3f805480",
X"f580518b",
X"cd3f8114",
X"5473a82e",
X"098106ef",
X"38868da0",
X"519cdd3f",
X"8052903d",
X"70525780",
X"c0fa3f83",
X"52765180",
X"c0f23f62",
X"818f3861",
X"802e80fb",
X"387b5473",
X"ff2e9638",
X"78802e81",
X"89387851",
X"e1dc3f83",
X"e08008ff",
X"155559e7",
X"3978802e",
X"80f43878",
X"51e1d83f",
X"83e08008",
X"802efc8e",
X"387851e1",
X"a03f83e0",
X"80085280",
X"f4f45183",
X"e33f83e0",
X"8008a338",
X"7c51859b",
X"3f83e080",
X"085574ff",
X"16565480",
X"7425ae38",
X"741d7033",
X"555673af",
X"2efecd38",
X"e9397851",
X"e0e13f83",
X"e0800852",
X"7c5184d3",
X"3f8f397f",
X"88296010",
X"057a0561",
X"055afc90",
X"3962802e",
X"fbd13880",
X"527651bf",
X"d33fa33d",
X"0d04803d",
X"0d9088b8",
X"337081ff",
X"0670842a",
X"81327081",
X"06515151",
X"5170802e",
X"8d38a80b",
X"9088b834",
X"b80b9088",
X"b8347083",
X"e0800c82",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067085",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d3898",
X"0b9088b8",
X"34b80b90",
X"88b83470",
X"83e0800c",
X"823d0d04",
X"930b9088",
X"bc34ff0b",
X"9088a834",
X"04ff3d0d",
X"028f0533",
X"52800b90",
X"88bc348a",
X"519aa53f",
X"df3f80f8",
X"0b9088a0",
X"34800b90",
X"888834fa",
X"12527190",
X"88803480",
X"0b908898",
X"34719088",
X"90349088",
X"b8528072",
X"34b87234",
X"833d0d04",
X"803d0d02",
X"8b053351",
X"709088b4",
X"34febf3f",
X"83e08008",
X"802ef638",
X"823d0d04",
X"803d0d84",
X"39a3fe3f",
X"fed93f83",
X"e0800880",
X"2ef33890",
X"88b43370",
X"81ff0683",
X"e0800c51",
X"823d0d04",
X"803d0da3",
X"0b9088bc",
X"34ff0b90",
X"88a83490",
X"88b851a8",
X"7134b871",
X"34823d0d",
X"04803d0d",
X"9088bc33",
X"7081c006",
X"70307080",
X"2583e080",
X"0c515151",
X"823d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"832a8132",
X"70810651",
X"51515170",
X"802ee838",
X"b00b9088",
X"b834b80b",
X"9088b834",
X"823d0d04",
X"803d0d90",
X"80ac0881",
X"0683e080",
X"0c823d0d",
X"04fd3d0d",
X"75775454",
X"80732594",
X"38737081",
X"05553352",
X"80f5ac51",
X"87843fff",
X"1353e939",
X"853d0d04",
X"fd3d0d75",
X"77535473",
X"33517089",
X"38713351",
X"70802ea1",
X"38733372",
X"33525372",
X"71278538",
X"ff519439",
X"70732785",
X"3881518b",
X"39811481",
X"135354d3",
X"39805170",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"77545472",
X"337081ff",
X"06525270",
X"802ea338",
X"7181ff06",
X"8114ffbf",
X"12535452",
X"70992689",
X"38a01270",
X"81ff0653",
X"51717470",
X"81055634",
X"d2398074",
X"34853d0d",
X"04ffbd3d",
X"0d80c63d",
X"0852a53d",
X"705254ff",
X"b33f80c7",
X"3d085285",
X"3d705253",
X"ffa63f72",
X"527351fe",
X"df3f80c5",
X"3d0d04fe",
X"3d0d7476",
X"53537170",
X"81055333",
X"51707370",
X"81055534",
X"70f03884",
X"3d0d04fe",
X"3d0d7452",
X"80723352",
X"5370732e",
X"8d388112",
X"81147133",
X"53545270",
X"f5387283",
X"e0800c84",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"b7fd3f83",
X"e080087a",
X"27ee3874",
X"802e80dd",
X"38745275",
X"51b7e83f",
X"83e08008",
X"75537652",
X"54b7ec3f",
X"83e08008",
X"7a537552",
X"56b7d03f",
X"83e08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"e08008c5",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9f",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fc813f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd53f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbb13f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83e0940c",
X"7183e098",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383e094",
X"085283e0",
X"980851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"bdba5351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fc3d",
X"0d765574",
X"83e39808",
X"2eaf3880",
X"53745187",
X"c13f83e0",
X"800881ff",
X"06ff1470",
X"81ff0672",
X"30709f2a",
X"51525553",
X"5472802e",
X"843871dd",
X"3873fe38",
X"7483e398",
X"0c863d0d",
X"04ff3d0d",
X"ff0b83e3",
X"980c84a5",
X"3f815187",
X"853f83e0",
X"800881ff",
X"065271ee",
X"3881d33f",
X"7183e080",
X"0c833d0d",
X"04fc3d0d",
X"76028405",
X"a2052202",
X"8805a605",
X"227a5455",
X"5555ff82",
X"3f72802e",
X"a03883e3",
X"ac143375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552dd",
X"39800b83",
X"e0800c86",
X"3d0d04fc",
X"3d0d7678",
X"7a115653",
X"55805371",
X"742e9338",
X"72155170",
X"3383e3ac",
X"13348112",
X"81145452",
X"ea39800b",
X"83e0800c",
X"863d0d04",
X"fd3d0d90",
X"5483e398",
X"085186f4",
X"3f83e080",
X"0881ff06",
X"ff157130",
X"71307073",
X"079f2a72",
X"9f2a0652",
X"55525553",
X"72db3885",
X"3d0d0480",
X"3d0d83e3",
X"a4081083",
X"e39c0807",
X"9080a80c",
X"823d0d04",
X"800b83e3",
X"a40ce43f",
X"04810b83",
X"e3a40cdb",
X"3f04ed3f",
X"047183e3",
X"a00c0480",
X"3d0d8051",
X"f43f810b",
X"83e3a40c",
X"810b83e3",
X"9c0cffbb",
X"3f823d0d",
X"04803d0d",
X"72307074",
X"07802583",
X"e39c0c51",
X"ffa53f82",
X"3d0d0480",
X"3d0d028b",
X"05339080",
X"a40c9080",
X"a8087081",
X"06515170",
X"f5389080",
X"a4087081",
X"ff0683e0",
X"800c5182",
X"3d0d0480",
X"3d0d81ff",
X"51d13f83",
X"e0800881",
X"ff0683e0",
X"800c823d",
X"0d04803d",
X"0d73902b",
X"73079080",
X"b40c823d",
X"0d0404fb",
X"3d0d7802",
X"84059f05",
X"3370982b",
X"55575572",
X"80259b38",
X"7580ff06",
X"56805280",
X"f751e03f",
X"83e08008",
X"81ff0654",
X"73812680",
X"ff388051",
X"fee73fff",
X"a23f8151",
X"fedf3fff",
X"9a3f7551",
X"feed3f74",
X"982a51fe",
X"e63f7490",
X"2a7081ff",
X"065253fe",
X"da3f7488",
X"2a7081ff",
X"065253fe",
X"ce3f7481",
X"ff0651fe",
X"c63f8155",
X"7580c02e",
X"09810686",
X"38819555",
X"8d397580",
X"c82e0981",
X"06843881",
X"87557451",
X"fea53f8a",
X"55fec83f",
X"83e08008",
X"81ff0670",
X"982b5454",
X"7280258c",
X"38ff1570",
X"81ff0656",
X"5374e238",
X"7383e080",
X"0c873d0d",
X"04fa3d0d",
X"fdc53f80",
X"51fdda3f",
X"8a54fe93",
X"3fff1470",
X"81ff0655",
X"5373f338",
X"73745355",
X"80c051fe",
X"a63f83e0",
X"800881ff",
X"06547381",
X"2e098106",
X"829f3883",
X"aa5280c8",
X"51fe8c3f",
X"83e08008",
X"81ff0653",
X"72812e09",
X"810681a8",
X"38745487",
X"3d741154",
X"56fdc83f",
X"83e08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e53802",
X"9a053353",
X"72812e09",
X"810681d9",
X"38029b05",
X"335380ce",
X"90547281",
X"aa2e8d38",
X"81c73980",
X"e4518acc",
X"3fff1454",
X"73802e81",
X"b838820a",
X"5281e951",
X"fda53f83",
X"e0800881",
X"ff065372",
X"de387252",
X"80fa51fd",
X"923f83e0",
X"800881ff",
X"06537281",
X"90387254",
X"731653fc",
X"d63f83e0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e8",
X"38873d33",
X"70862a70",
X"81065154",
X"548c5572",
X"80e33884",
X"5580de39",
X"745281e9",
X"51fccc3f",
X"83e08008",
X"81ff0653",
X"825581e9",
X"56817327",
X"86387355",
X"80c15680",
X"ce90548a",
X"3980e451",
X"89be3fff",
X"14547380",
X"2ea93880",
X"527551fc",
X"9a3f83e0",
X"800881ff",
X"065372e1",
X"38848052",
X"80d051fc",
X"863f83e0",
X"800881ff",
X"06537280",
X"2e833880",
X"557483e3",
X"a8348051",
X"fb873ffb",
X"c23f883d",
X"0d04fb3d",
X"0d775480",
X"0b83e3a8",
X"3370832a",
X"70810651",
X"55575572",
X"752e0981",
X"06853873",
X"892b5473",
X"5280d151",
X"fbbd3f83",
X"e0800881",
X"ff065372",
X"bd3882b8",
X"c054fb83",
X"3f83e080",
X"0881ff06",
X"537281ff",
X"2e098106",
X"8938ff14",
X"5473e738",
X"9f397281",
X"fe2e0981",
X"06963883",
X"e7ac5283",
X"e3ac51fa",
X"ed3ffad3",
X"3ffad03f",
X"83398155",
X"8051fa89",
X"3ffac43f",
X"7481ff06",
X"83e0800c",
X"873d0d04",
X"fb3d0d77",
X"83e3ac56",
X"548151f9",
X"ec3f83e3",
X"a8337083",
X"2a708106",
X"51545672",
X"85387389",
X"2b547352",
X"80d851fa",
X"b63f83e0",
X"800881ff",
X"06537280",
X"e43881ff",
X"51f9d43f",
X"81fe51f9",
X"ce3f8480",
X"53747081",
X"05563351",
X"f9c13fff",
X"137083ff",
X"ff065153",
X"72eb3872",
X"51f9b03f",
X"7251f9ab",
X"3ff9d03f",
X"83e08008",
X"9f0653a7",
X"88547285",
X"2e8c3899",
X"3980e451",
X"86f63fff",
X"1454f9b3",
X"3f83e080",
X"0881ff2e",
X"843873e9",
X"388051f8",
X"e43ff99f",
X"3f800b83",
X"e0800c87",
X"3d0d0471",
X"83e7b00c",
X"8880800b",
X"83e7ac0c",
X"8480800b",
X"83e7b40c",
X"04fd3d0d",
X"77701755",
X"7705ff1a",
X"535371ff",
X"2e943873",
X"70810555",
X"33517073",
X"70810555",
X"34ff1252",
X"e939853d",
X"0d04fc3d",
X"0d87a681",
X"55743383",
X"e7b834a0",
X"5483a080",
X"5383e7b0",
X"085283e7",
X"ac0851ff",
X"b83fa054",
X"83a48053",
X"83e7b008",
X"5283e7ac",
X"0851ffa5",
X"3f905483",
X"a8805383",
X"e7b00852",
X"83e7ac08",
X"51ff923f",
X"a0538052",
X"83e7b408",
X"83a08005",
X"5185ce3f",
X"a0538052",
X"83e7b408",
X"83a48005",
X"5185be3f",
X"90538052",
X"83e7b408",
X"83a88005",
X"5185ae3f",
X"ff753483",
X"a0805480",
X"5383e7b0",
X"085283e7",
X"b40851fe",
X"cc3f80d0",
X"805483b0",
X"805383e7",
X"b0085283",
X"e7b40851",
X"feb73f86",
X"e13fa254",
X"805383e7",
X"b4088c80",
X"055280f7",
X"fc51fea1",
X"3f860b87",
X"a8833480",
X"0b87a882",
X"34800b87",
X"a09a34af",
X"0b87a096",
X"34bf0b87",
X"a0973480",
X"0b87a098",
X"349f0b87",
X"a0993480",
X"0b87a09b",
X"34e00b87",
X"a88934a2",
X"0b87a880",
X"34830b87",
X"a48f3482",
X"0b87a881",
X"34863d0d",
X"04fd3d0d",
X"83a08054",
X"805383e7",
X"b4085283",
X"e7b00851",
X"fdbf3f80",
X"d0805483",
X"b0805383",
X"e7b40852",
X"83e7b008",
X"51fdaa3f",
X"a05483a0",
X"805383e7",
X"b4085283",
X"e7b00851",
X"fd973fa0",
X"5483a480",
X"5383e7b4",
X"085283e7",
X"b00851fd",
X"843f9054",
X"83a88053",
X"83e7b408",
X"5283e7b0",
X"0851fcf1",
X"3f83e7b8",
X"3387a681",
X"34853d0d",
X"04803d0d",
X"90809008",
X"810683e0",
X"800c823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087081",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fd0676",
X"1007720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870822c",
X"bf0683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe830676",
X"822b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087088",
X"2c870683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f1ff06",
X"76882b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"8b2cbf06",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f88f",
X"ff06768b",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870912c",
X"bf0683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fc87ffff",
X"0676912b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70992c81",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870ff",
X"bf0a0676",
X"992b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"80087088",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"892c8106",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708a2c81",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708b2c",
X"810683e0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708c",
X"2cbf0683",
X"e0800c51",
X"823d0d04",
X"fe3d0d74",
X"81e62987",
X"2a9080a0",
X"0c843d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727081",
X"055434ff",
X"1151f039",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708405",
X"540cff11",
X"51f03984",
X"3d0d04fe",
X"3d0d8480",
X"80538052",
X"88800a51",
X"ffb33f81",
X"80805380",
X"5282800a",
X"51c63f84",
X"3d0d0480",
X"3d0d8151",
X"fbfc3f72",
X"802e9038",
X"8051fdfe",
X"3fcd3f83",
X"e7bc3351",
X"fdf43f81",
X"51fc8d3f",
X"8051fc88",
X"3f8051fb",
X"d93f823d",
X"0d04fd3d",
X"0d755280",
X"5480ff72",
X"25883881",
X"0bff8013",
X"5354ffbf",
X"12517099",
X"268638e0",
X"12529e39",
X"ff9f1251",
X"99712795",
X"38d012e0",
X"13705454",
X"51897127",
X"88388f73",
X"27833880",
X"5273802e",
X"85388180",
X"12527181",
X"ff0683e0",
X"800c853d",
X"0d04803d",
X"0d84d8c0",
X"51807170",
X"81055334",
X"7084e0c0",
X"2e098106",
X"f038823d",
X"0d04fe3d",
X"0d029705",
X"3351ff86",
X"3f83e080",
X"0881ff06",
X"83e7c008",
X"54528073",
X"249b3883",
X"e7e00813",
X"7283e7e4",
X"08075353",
X"71733483",
X"e7c00881",
X"0583e7c0",
X"0c843d0d",
X"04fa3d0d",
X"82800a1b",
X"55805788",
X"3dfc0554",
X"79537452",
X"7851ffbb",
X"893f883d",
X"0d04fe3d",
X"0d83e7d8",
X"08527451",
X"c1ed3f83",
X"e080088c",
X"38765375",
X"5283e7d8",
X"0851c63f",
X"843d0d04",
X"fe3d0d83",
X"e7d80853",
X"75527451",
X"ffbcab3f",
X"83e08008",
X"8d387753",
X"765283e7",
X"d80851ff",
X"a03f843d",
X"0d04fe3d",
X"0d83e7d8",
X"0851ffbb",
X"9e3f83e0",
X"80088180",
X"802e0981",
X"06883883",
X"c1808053",
X"9c3983e7",
X"d80851ff",
X"bb813f83",
X"e0800880",
X"d0802e09",
X"81069338",
X"83c1b080",
X"5383e080",
X"085283e7",
X"d80851fe",
X"d43f843d",
X"0d04803d",
X"0df9e03f",
X"83e08008",
X"842980f8",
X"a0057008",
X"83e0800c",
X"51823d0d",
X"04ed3d0d",
X"80448043",
X"80428041",
X"80705a5b",
X"fdcc3f80",
X"0b83e7c0",
X"0c800b83",
X"e7e40c80",
X"f5f851ea",
X"a53f8180",
X"0b83e7e4",
X"0c80f5fc",
X"51ea973f",
X"80d00b83",
X"e7c00c78",
X"30707a07",
X"80257087",
X"2b83e7e4",
X"0c5155f8",
X"d13f83e0",
X"80085280",
X"f68451e9",
X"f13f80f8",
X"0b83e7c0",
X"0c788132",
X"70307072",
X"07802570",
X"872b83e7",
X"e40c5156",
X"56feef3f",
X"83e08008",
X"5280f690",
X"51e9c73f",
X"81a00b83",
X"e7c00c78",
X"82327030",
X"70720780",
X"2570872b",
X"83e7e40c",
X"515683e7",
X"d8085256",
X"ffb6a63f",
X"83e08008",
X"5280f698",
X"51e9973f",
X"81f00b83",
X"e7c00c81",
X"0b83e7c4",
X"5b5883e7",
X"c0088219",
X"7a327030",
X"70720780",
X"2570872b",
X"83e7e40c",
X"51578e3d",
X"7055ff1b",
X"54575757",
X"99fb3f79",
X"7084055b",
X"0851ffb5",
X"dc3f7454",
X"83e08008",
X"53775280",
X"f6a051e8",
X"c93fa817",
X"83e7c00c",
X"81185877",
X"852e0981",
X"06ffaf38",
X"83900b83",
X"e7c00c78",
X"87327030",
X"70720780",
X"2570872b",
X"83e7e40c",
X"515656f7",
X"f53f80f6",
X"b05583e0",
X"8008802e",
X"8f3883e7",
X"d40851ff",
X"b5873f83",
X"e0800855",
X"745280f6",
X"b851e7f6",
X"3f83e00b",
X"83e7c00c",
X"78883270",
X"30707207",
X"80257087",
X"2b83e7e4",
X"0c515780",
X"f6c45255",
X"e7d43f86",
X"8da051f8",
X"ef3f8052",
X"913d7052",
X"559d8d3f",
X"83527451",
X"9d863f63",
X"557482fa",
X"38611959",
X"78802585",
X"38745990",
X"39887925",
X"85388859",
X"87397888",
X"2682d938",
X"78822b55",
X"80f4d015",
X"0804f5e2",
X"3f83e080",
X"08615755",
X"75812e09",
X"81068938",
X"83e08008",
X"10559039",
X"75ff2e09",
X"81068838",
X"83e08008",
X"812c5590",
X"75258538",
X"90558839",
X"74802483",
X"38815574",
X"51f5bc3f",
X"828e39f5",
X"ce3f83e0",
X"80086105",
X"55748025",
X"85388055",
X"88398775",
X"25833887",
X"557451f5",
X"c73f81ec",
X"39608738",
X"62802e81",
X"e33883e3",
X"8c0883e3",
X"880cade5",
X"0b83e390",
X"0c83e7d8",
X"0851d78b",
X"3ffadb3f",
X"81c63960",
X"56807625",
X"9838ad84",
X"0b83e390",
X"0c83e7b8",
X"15700852",
X"55d6ec3f",
X"74085292",
X"39758025",
X"923883e7",
X"b8150851",
X"ffb2f03f",
X"8052fd19",
X"51b83962",
X"802e818c",
X"3883e7b8",
X"15700883",
X"e7c40872",
X"0c83e7c4",
X"0cfd1a70",
X"5351558b",
X"f63f83e0",
X"80085680",
X"518bec3f",
X"83e08008",
X"52745188",
X"833f7552",
X"805187fc",
X"3f80d539",
X"60558075",
X"25b63883",
X"e3940883",
X"e3880cad",
X"e50b83e3",
X"900c83e7",
X"d40851d5",
X"f63f83e7",
X"d40851d3",
X"973f83e0",
X"800881ff",
X"06705255",
X"f4d53f74",
X"802e9d38",
X"8155a139",
X"74802594",
X"3883e7d4",
X"0851ffb1",
X"e23f8051",
X"f4b93f84",
X"39628738",
X"7a802efa",
X"83388055",
X"7483e080",
X"0c953d0d",
X"04fe3d0d",
X"f4e53f83",
X"e0800880",
X"2e863880",
X"51818a39",
X"f4ea3f83",
X"e0800880",
X"fe38f58a",
X"3f83e080",
X"08802eb9",
X"388151f2",
X"993f8051",
X"f4a03fef",
X"8d3f800b",
X"83e7c00c",
X"f9ab3f83",
X"e0800853",
X"ff0b83e7",
X"c00cf0f9",
X"3f7280cb",
X"3883e7bc",
X"3351f3fa",
X"3f7251f1",
X"e93f80c0",
X"39f4b23f",
X"83e08008",
X"802eb538",
X"8151f1d6",
X"3f8051f3",
X"dd3feeca",
X"3fad840b",
X"83e3900c",
X"83e7c408",
X"51d4a83f",
X"ff0b83e7",
X"c00cf0b5",
X"3f83e7c4",
X"08528051",
X"85fa3f81",
X"51f5a43f",
X"843d0d04",
X"fb3d0d80",
X"0b83e7bc",
X"34908080",
X"52868480",
X"8051ffb4",
X"9b3f83e0",
X"80088197",
X"3889c53f",
X"80f9f451",
X"ffb8da3f",
X"83e08008",
X"559c800a",
X"5480c080",
X"5380f6cc",
X"5283e080",
X"0851f6f8",
X"3f83e7d8",
X"085380f6",
X"dc527451",
X"ffb3a33f",
X"83e08008",
X"8438f786",
X"3f83e7dc",
X"085380f6",
X"e8527451",
X"ffb38b3f",
X"83e08008",
X"b638873d",
X"fc055484",
X"80805386",
X"a8808052",
X"83e7dc08",
X"51ffb196",
X"3f83e080",
X"08933875",
X"8480802e",
X"09810689",
X"38810b83",
X"e7bc3487",
X"39800b83",
X"e7bc3483",
X"e7bc3351",
X"f2843f81",
X"51f3f03f",
X"92ee3f81",
X"51f3e83f",
X"8151fda1",
X"3ffa3983",
X"e08c0802",
X"83e08c0c",
X"fb3d0d02",
X"80f6f40b",
X"83e38c0c",
X"80f6f80b",
X"83e3840c",
X"80f6fc0b",
X"83e3940c",
X"83e08c08",
X"fc050c80",
X"0b83e7c4",
X"0b83e08c",
X"08f8050c",
X"83e08c08",
X"f4050cff",
X"b1a63f83",
X"e0800886",
X"05fc0683",
X"e08c08f0",
X"050c0283",
X"e08c08f0",
X"0508310d",
X"833d7083",
X"e08c08f8",
X"05087084",
X"0583e08c",
X"08f8050c",
X"0c51ffad",
X"ee3f83e0",
X"8c08f405",
X"08810583",
X"e08c08f4",
X"050c83e0",
X"8c08f405",
X"08872e09",
X"8106ffab",
X"38869480",
X"8051eb83",
X"3fff0b83",
X"e7c00c80",
X"0b83e7e4",
X"0c84d8c0",
X"0b83e7e0",
X"0c8151ee",
X"ad3f8151",
X"eed23f80",
X"51eecd3f",
X"8151eef3",
X"3f8151ef",
X"c83f8251",
X"ef963f80",
X"51efec3f",
X"8051f096",
X"3f80d0ca",
X"528051df",
X"e23ffcdc",
X"3f83e08c",
X"08fc0508",
X"0d800b83",
X"e0800c87",
X"3d0d83e0",
X"8c0c0480",
X"3d0d81ff",
X"51800b83",
X"e7f01234",
X"ff115170",
X"f438823d",
X"0d04ff3d",
X"0d737033",
X"53518111",
X"33713471",
X"81123483",
X"3d0d04fb",
X"3d0d7779",
X"56568070",
X"71555552",
X"717525ac",
X"38721670",
X"33701470",
X"81ff0655",
X"51515171",
X"74278938",
X"81127081",
X"ff065351",
X"71811470",
X"83ffff06",
X"55525474",
X"7324d638",
X"7183e080",
X"0c873d0d",
X"04fb3d0d",
X"7756d7ac",
X"3f83e080",
X"08802ef6",
X"3883ea8c",
X"08860570",
X"81ff0652",
X"53d5ae3f",
X"810b9088",
X"d4349088",
X"d4337081",
X"ff065153",
X"728b38f9",
X"fc3f8351",
X"efca3fea",
X"39805574",
X"1675822b",
X"54549088",
X"c0133374",
X"34811555",
X"74852e09",
X"8106e838",
X"810b9088",
X"d4347533",
X"83e7f034",
X"81163383",
X"e7f13482",
X"163383e7",
X"f2348316",
X"3383e7f3",
X"34845283",
X"e7f051fe",
X"ba3f83e0",
X"800881ff",
X"06841733",
X"57537276",
X"2e098106",
X"8c38d5d5",
X"3f83e080",
X"08802e9a",
X"3883ea8c",
X"08a82e09",
X"81068938",
X"860b83ea",
X"8c0c8739",
X"a80b83ea",
X"8c0c80e4",
X"51eec53f",
X"873d0d04",
X"f43d0d7e",
X"60595580",
X"5d807582",
X"2b7183ea",
X"90120c83",
X"eaa4175b",
X"5b577679",
X"3477772e",
X"83b93876",
X"527751ff",
X"acb43f8e",
X"3dfc0554",
X"905383e9",
X"f8527751",
X"ffabef3f",
X"7c567590",
X"2e098106",
X"83953883",
X"e9f851fd",
X"953f83e9",
X"fa51fd8e",
X"3f83e9fc",
X"51fd873f",
X"7683ea88",
X"0c7751ff",
X"a9bb3f0b",
X"0b80f588",
X"5283e080",
X"0851cbd2",
X"3f83e080",
X"08812e09",
X"810680d4",
X"387683ea",
X"a00c820b",
X"83e9f834",
X"ff960b83",
X"e9f93477",
X"51ffabff",
X"3f83e080",
X"085583e0",
X"80087725",
X"883883e0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83e9fa34",
X"7483e9fb",
X"347683e9",
X"fc34ff80",
X"0b83e9fd",
X"34819039",
X"83e9f833",
X"83e9f933",
X"71882b07",
X"565b7483",
X"ffff2e09",
X"810680e8",
X"38fe800b",
X"83eaa00c",
X"810b83ea",
X"880cff0b",
X"83e9f834",
X"ff0b83e9",
X"f9347751",
X"ffab8c3f",
X"83e08008",
X"83eaa80c",
X"83e08008",
X"5583e080",
X"08802588",
X"3883e080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"e9fa3474",
X"83e9fb34",
X"7683e9fc",
X"34ff800b",
X"83e9fd34",
X"810b83ea",
X"8734a539",
X"7485962e",
X"09810680",
X"fe387583",
X"eaa00c77",
X"51ffaac0",
X"3f83ea87",
X"3383e080",
X"08075574",
X"83ea8734",
X"83ea8733",
X"81065574",
X"802e8338",
X"845783e9",
X"fc3383e9",
X"fd337188",
X"2b07565c",
X"7481802e",
X"098106a1",
X"3883e9fa",
X"3383e9fb",
X"3371882b",
X"07565bad",
X"80752787",
X"38768207",
X"579c3976",
X"81075796",
X"39748280",
X"2e098106",
X"87387683",
X"07578739",
X"7481ff26",
X"8a387783",
X"ea901b0c",
X"7679348e",
X"3d0d0480",
X"3d0d7284",
X"2983ea90",
X"05700883",
X"e0800c51",
X"823d0d04",
X"fe3d0d80",
X"0b83e9f4",
X"0c800b83",
X"e9f00cff",
X"0b83e7ec",
X"0ca80b83",
X"ea8c0cae",
X"51cff63f",
X"800b83ea",
X"90545280",
X"73708405",
X"550c8112",
X"5271842e",
X"098106ef",
X"38843d0d",
X"04fe3d0d",
X"74028405",
X"96052253",
X"5371802e",
X"96387270",
X"81055433",
X"51d0813f",
X"ff127083",
X"ffff0651",
X"52e73984",
X"3d0d04fe",
X"3d0d0292",
X"05225382",
X"ac51e9d8",
X"3f80c351",
X"cfde3f81",
X"9651e9cc",
X"3f725283",
X"e7f051ff",
X"b43f7252",
X"83e7f051",
X"f8f13f83",
X"e0800881",
X"ff0651cf",
X"bb3f843d",
X"0d04ffb1",
X"3d0d80d1",
X"3df80551",
X"f99b3f83",
X"e9f40881",
X"0583e9f4",
X"0c80cf3d",
X"33cf1170",
X"81ff0651",
X"56567483",
X"2688e238",
X"758f06ff",
X"05567583",
X"e7ec082e",
X"9b387583",
X"26963875",
X"83e7ec0c",
X"75842983",
X"ea900570",
X"08535575",
X"51fa993f",
X"80762488",
X"be387584",
X"2983ea90",
X"05557408",
X"802e88af",
X"3883e7ec",
X"08842983",
X"ea900570",
X"08028805",
X"82b90533",
X"525b5574",
X"80d22e84",
X"ac387480",
X"d2249038",
X"74bf2e9c",
X"387480d0",
X"2e81d138",
X"87ee3974",
X"80d32e80",
X"cf387480",
X"d72e81c0",
X"3887dd39",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"055656ce",
X"b73f80c1",
X"51cdf13f",
X"f6ed3f86",
X"0b83e7f0",
X"34815283",
X"e7f051cf",
X"943f8151",
X"fde93f74",
X"8938860b",
X"83ea8c0c",
X"8739a80b",
X"83ea8c0c",
X"ce863f80",
X"c151cdc0",
X"3ff6bc3f",
X"900b83ea",
X"87338106",
X"56567480",
X"2e833898",
X"5683e9fc",
X"3383e9fd",
X"3371882b",
X"07565974",
X"81802e09",
X"81069c38",
X"83e9fa33",
X"83e9fb33",
X"71882b07",
X"5657ad80",
X"75278c38",
X"75818007",
X"56853975",
X"a0075675",
X"83e7f034",
X"ff0b83e7",
X"f134e00b",
X"83e7f234",
X"800b83e7",
X"f3348452",
X"83e7f051",
X"ce8b3f84",
X"51869b39",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"055659cc",
X"fb3f7951",
X"ffa5913f",
X"83e08008",
X"802e8a38",
X"80ce51cc",
X"a73f85f1",
X"3980c151",
X"cc9e3fcd",
X"933fcbc8",
X"3f83eaa0",
X"08588375",
X"259b3883",
X"e9fc3383",
X"e9fd3371",
X"882b07fc",
X"1771297a",
X"05838005",
X"5a51578d",
X"39748180",
X"2918ff80",
X"05588180",
X"57805676",
X"762e9238",
X"cbfa3f83",
X"e0800883",
X"e7f01734",
X"811656eb",
X"39cbe93f",
X"83e08008",
X"81ff0677",
X"5383e7f0",
X"5256f4e7",
X"3f83e080",
X"0881ff06",
X"5575752e",
X"09810681",
X"95389451",
X"e59a3fcb",
X"e33f80c1",
X"51cb9d3f",
X"cc923f77",
X"527951ff",
X"a3a43f80",
X"5e80d13d",
X"fdf40554",
X"765383e7",
X"f0527951",
X"ffa1b13f",
X"0282b905",
X"33558159",
X"7480d72e",
X"09810680",
X"c5387752",
X"7951ffa2",
X"f53f80d1",
X"3dfdf005",
X"5476538f",
X"3d70537a",
X"5258ffa2",
X"ad3f8056",
X"76762ea2",
X"38751883",
X"e7f01733",
X"71337072",
X"32703070",
X"80257030",
X"7f06811d",
X"5d5f5151",
X"51525b55",
X"db3982ac",
X"51e4953f",
X"78802e86",
X"3880c351",
X"843980ce",
X"51ca913f",
X"cb863fc9",
X"bb3f83d8",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055955",
X"80705d59",
X"80e451e3",
X"df3fcaa8",
X"3f80c151",
X"c9e23f83",
X"ea880879",
X"2e82d638",
X"83eaa808",
X"80fc0555",
X"80fd5274",
X"5185a03f",
X"83e08008",
X"5b778224",
X"b238ff18",
X"70872b83",
X"ffff8006",
X"80f8c005",
X"83e7f059",
X"57558180",
X"55757081",
X"05573377",
X"70810559",
X"34ff1570",
X"81ff0651",
X"5574ea38",
X"82853977",
X"82e82e81",
X"a3387782",
X"e92e0981",
X"0681aa38",
X"78587787",
X"32703070",
X"72078025",
X"7a8a3270",
X"30707207",
X"80257307",
X"53545a51",
X"57557580",
X"2e973878",
X"78269238",
X"a00b83e7",
X"f01a3481",
X"197081ff",
X"065a55eb",
X"39811870",
X"81ff0659",
X"558a7827",
X"ffbc388f",
X"5883e7eb",
X"183383e7",
X"f01934ff",
X"187081ff",
X"06595577",
X"8426ea38",
X"9058800b",
X"83e7f019",
X"34811870",
X"81ff0670",
X"982b5259",
X"55748025",
X"e93880c6",
X"557a858f",
X"24843880",
X"c2557483",
X"e7f03480",
X"f10b83e7",
X"f334810b",
X"83e7f434",
X"7a83e7f1",
X"347a882c",
X"557483e7",
X"f23480cb",
X"3982f078",
X"2580c438",
X"7780fd29",
X"fd97d305",
X"527951ff",
X"9fd03f80",
X"d13dfdec",
X"055480fd",
X"5383e7f0",
X"527951ff",
X"9f883f7b",
X"81195956",
X"7580fc24",
X"83387858",
X"77882c55",
X"7483e8ed",
X"347783e8",
X"ee347583",
X"e8ef3481",
X"805980cc",
X"3983eaa0",
X"08578378",
X"259b3883",
X"e9fc3383",
X"e9fd3371",
X"882b07fc",
X"1a712979",
X"05838005",
X"5951598d",
X"39778180",
X"2917ff80",
X"05578180",
X"59765279",
X"51ff9ede",
X"3f80d13d",
X"fdec0554",
X"785383e7",
X"f0527951",
X"ff9e973f",
X"7851f6c3",
X"3fc7a93f",
X"c5de3f8b",
X"3983e9f0",
X"08810583",
X"e9f00c80",
X"d13d0d04",
X"f6e43ffc",
X"39fc3d0d",
X"76787184",
X"2983ea90",
X"05700851",
X"53535370",
X"9e3880ce",
X"723480cf",
X"0b811334",
X"80ce0b82",
X"133480c5",
X"0b831334",
X"70841334",
X"80e73983",
X"eaa41333",
X"5480d272",
X"3473822a",
X"70810651",
X"5180cf53",
X"70843880",
X"d7537281",
X"1334a00b",
X"82133473",
X"83065170",
X"812e9e38",
X"70812488",
X"3870802e",
X"8f389f39",
X"70822e92",
X"3870832e",
X"92389339",
X"80d8558e",
X"3980d355",
X"893980cd",
X"55843980",
X"c4557483",
X"133480c4",
X"0b841334",
X"800b8513",
X"34863d0d",
X"04fc3d0d",
X"76785354",
X"81538055",
X"87397110",
X"73105452",
X"73722651",
X"72802ea7",
X"3870802e",
X"86387180",
X"25e83872",
X"802e9838",
X"71742689",
X"38737231",
X"75740756",
X"5472812a",
X"72812a53",
X"53e53973",
X"51788338",
X"74517083",
X"e0800c86",
X"3d0d04fe",
X"3d0d8053",
X"75527451",
X"ffa33f84",
X"3d0d04fe",
X"3d0d8153",
X"75527451",
X"ff933f84",
X"3d0d04fb",
X"3d0d7779",
X"55558056",
X"74762586",
X"38743055",
X"81567380",
X"25883873",
X"30768132",
X"57548053",
X"73527451",
X"fee73f83",
X"e0800854",
X"75802e87",
X"3883e080",
X"08305473",
X"83e0800c",
X"873d0d04",
X"fa3d0d78",
X"7a575580",
X"57747725",
X"86387430",
X"55815775",
X"9f2c5481",
X"53757432",
X"74315274",
X"51feaa3f",
X"83e08008",
X"5476802e",
X"873883e0",
X"80083054",
X"7383e080",
X"0c883d0d",
X"04fd3d0d",
X"75548074",
X"0c800b84",
X"150c800b",
X"88150c80",
X"0b8c150c",
X"87a68033",
X"7081ff06",
X"5151dcc7",
X"3f70812a",
X"81327181",
X"32718106",
X"71810631",
X"84170c53",
X"5370832a",
X"81327182",
X"2a813271",
X"81067181",
X"0631760c",
X"525287a0",
X"90337009",
X"81068816",
X"0c5183e0",
X"8008802e",
X"80c23883",
X"e0800881",
X"2a708106",
X"83e08008",
X"81063184",
X"160c5183",
X"e0800883",
X"2a83e080",
X"08822a71",
X"81067181",
X"0631760c",
X"525283e0",
X"8008842a",
X"81068815",
X"0c83e080",
X"08852a81",
X"068c150c",
X"853d0d04",
X"fe3d0d74",
X"76545271",
X"51fece3f",
X"72812ea2",
X"38817326",
X"8d387282",
X"2ea83872",
X"832e9c38",
X"e6397108",
X"e2388412",
X"08dd3888",
X"1208d838",
X"a5398812",
X"08812e9e",
X"38913988",
X"1208812e",
X"95387108",
X"91388412",
X"088c388c",
X"1208812e",
X"098106ff",
X"b238843d",
X"0d040000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002b0a",
X"00002b4b",
X"00002b6d",
X"00002b93",
X"00002b93",
X"00002b93",
X"00002b93",
X"00002c04",
X"00002c55",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"66726565",
X"7a65722e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00003ab4",
X"00003ab8",
X"00003ac0",
X"00003acc",
X"00003ad8",
X"00003ae4",
X"00003af0",
X"00003af4",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
