
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f2",
X"a4738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80f5",
X"dc0c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f1",
X"e42d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580f1a3",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80da9c04",
X"f93d0d80",
X"0b83e080",
X"0c893d0d",
X"04fc3d0d",
X"76705255",
X"b3a83f83",
X"e0800815",
X"ff055473",
X"752e8e38",
X"73335372",
X"ae2e8638",
X"ff1454ef",
X"39775281",
X"1451b2c0",
X"3f83e080",
X"08307083",
X"e0800807",
X"802583e0",
X"800c5386",
X"3d0d04fc",
X"3d0d7670",
X"525599e0",
X"3f83e080",
X"08548153",
X"83e08008",
X"80c73874",
X"5199a33f",
X"83e08008",
X"0b0b80f3",
X"e45383e0",
X"80085253",
X"ff8f3f83",
X"e08008a5",
X"380b0b80",
X"f3e85272",
X"51fefe3f",
X"83e08008",
X"94380b0b",
X"80f3ec52",
X"7251feed",
X"3f83e080",
X"08802e83",
X"38815473",
X"537283e0",
X"800c863d",
X"0d04fd3d",
X"0d757052",
X"5498f93f",
X"815383e0",
X"80089838",
X"735198c2",
X"3f83e0a0",
X"085283e0",
X"800851fe",
X"b43f83e0",
X"80085372",
X"83e0800c",
X"853d0d04",
X"df3d0da4",
X"3d087052",
X"5e8ee73f",
X"83e08008",
X"33953d56",
X"54739638",
X"80f8e052",
X"7451b19a",
X"3f9a397d",
X"52785191",
X"e83f84e3",
X"397d518e",
X"cd3f83e0",
X"80085274",
X"518dfd3f",
X"80438042",
X"80418040",
X"83e0a808",
X"52943d70",
X"525d94d0",
X"3f83e080",
X"0859800b",
X"83e08008",
X"555b83e0",
X"80087b2e",
X"9438811b",
X"74525b97",
X"d23f83e0",
X"80085483",
X"e08008ee",
X"38805aff",
X"5f790970",
X"9f2c7b06",
X"5b547a7a",
X"248438ff",
X"1b5af61a",
X"7009709f",
X"2c72067b",
X"ff125a5a",
X"52555580",
X"75259538",
X"76519797",
X"3f83e080",
X"0876ff18",
X"58555773",
X"8024ed38",
X"747f2e87",
X"3880c2fa",
X"3f745f78",
X"ff1b7058",
X"5d58807a",
X"25953877",
X"5196ec3f",
X"83e08008",
X"76ff1858",
X"55587380",
X"24ed3880",
X"0b83e7c0",
X"0c800b83",
X"e7e40c0b",
X"0b80f3f0",
X"518bbe3f",
X"81800b83",
X"e7e40c0b",
X"0b80f3f8",
X"518bae3f",
X"a80b83e7",
X"c00c7680",
X"2e80e838",
X"83e7c008",
X"77793270",
X"30707207",
X"80257087",
X"2b83e7e4",
X"0c515678",
X"53565696",
X"9f3f83e0",
X"8008802e",
X"8a380b0b",
X"80f48051",
X"8af33f76",
X"5195df3f",
X"83e08008",
X"520b0b80",
X"f58c518a",
X"e03f7651",
X"95e53f83",
X"e0800883",
X"e7c00855",
X"57757425",
X"8638a816",
X"56f73975",
X"83e7c00c",
X"86f07624",
X"ff943887",
X"980b83e7",
X"c00c7780",
X"2eb73877",
X"51959b3f",
X"83e08008",
X"78525595",
X"bb3f0b0b",
X"80f48854",
X"83e08008",
X"8f388739",
X"80763481",
X"d8390b0b",
X"80f48454",
X"74537352",
X"0b0b80f3",
X"d85189f9",
X"3f80540b",
X"0b80f5d8",
X"5189ee3f",
X"81145473",
X"a82e0981",
X"06ed3886",
X"8da051be",
X"ef3f8052",
X"903d7052",
X"5780e0d7",
X"3f835276",
X"5180e0cf",
X"3f628191",
X"3861802e",
X"80fd387b",
X"5473ff2e",
X"96387880",
X"2e818c38",
X"785194b7",
X"3f83e080",
X"08ff1555",
X"59e73978",
X"802e80f7",
X"38785194",
X"b33f83e0",
X"8008802e",
X"fbfd3878",
X"5193fb3f",
X"83e08008",
X"520b0b80",
X"f3e051ab",
X"da3f83e0",
X"8008a338",
X"7c51ad92",
X"3f83e080",
X"085574ff",
X"16565480",
X"7425ae38",
X"741d7033",
X"555673af",
X"2efec538",
X"e9397851",
X"93ba3f83",
X"e0800852",
X"7c51acca",
X"3f8f397f",
X"88296010",
X"057a0561",
X"055afbfd",
X"3962802e",
X"fbbe3880",
X"52765180",
X"dfad3fa3",
X"3d0d0480",
X"3d0d9080",
X"f8337081",
X"ff067084",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d38a8",
X"0b9080f8",
X"34b80b90",
X"80f83470",
X"83e0800c",
X"823d0d04",
X"803d0d90",
X"80f83370",
X"81ff0670",
X"852a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"980b9080",
X"f834b80b",
X"9080f834",
X"7083e080",
X"0c823d0d",
X"04930b90",
X"80fc34ff",
X"0b9080e8",
X"3404ff3d",
X"0d028f05",
X"3352800b",
X"9080fc34",
X"8a51bcb4",
X"3fdf3f80",
X"f80b9080",
X"e034800b",
X"9080c834",
X"fa125271",
X"9080c034",
X"800b9080",
X"d8347190",
X"80d03490",
X"80f85280",
X"7234b872",
X"34833d0d",
X"04803d0d",
X"028b0533",
X"51709080",
X"f434febf",
X"3f83e080",
X"08802ef6",
X"38823d0d",
X"04803d0d",
X"853980c6",
X"833ffed8",
X"3f83e080",
X"08802ef2",
X"389080f4",
X"337081ff",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0da30b90",
X"80fc34ff",
X"0b9080e8",
X"349080f8",
X"51a87134",
X"b8713482",
X"3d0d0480",
X"3d0d9080",
X"fc337081",
X"c0067030",
X"70802583",
X"e0800c51",
X"5151823d",
X"0d04803d",
X"0d9080f8",
X"337081ff",
X"0670832a",
X"81327081",
X"06515151",
X"5170802e",
X"e838b00b",
X"9080f834",
X"b80b9080",
X"f834823d",
X"0d04803d",
X"0d9080ac",
X"08810683",
X"e0800c82",
X"3d0d04fd",
X"3d0d7577",
X"54548073",
X"25943873",
X"70810555",
X"335280f4",
X"8c5185a1",
X"3fff1353",
X"e939853d",
X"0d04f63d",
X"0d7c7e60",
X"625a5d5b",
X"56805981",
X"55853974",
X"7a295574",
X"52755180",
X"ddad3f83",
X"e080087a",
X"27ed3874",
X"802e80e0",
X"38745275",
X"5180dd97",
X"3f83e080",
X"08755376",
X"525480dd",
X"9a3f83e0",
X"80087a53",
X"75525680",
X"dcfd3f83",
X"e0800879",
X"30707b07",
X"9f2a7077",
X"80240751",
X"51545572",
X"873883e0",
X"8008c238",
X"768118b0",
X"16555858",
X"8974258b",
X"38b71453",
X"7a853880",
X"d7145372",
X"78348119",
X"59ff9c39",
X"8077348c",
X"3d0d04f7",
X"3d0d7b7d",
X"7f620290",
X"05bb0533",
X"5759565a",
X"5ab05872",
X"8338a058",
X"75707081",
X"05523371",
X"59545590",
X"39807425",
X"8e38ff14",
X"77708105",
X"59335454",
X"72ef3873",
X"ff155553",
X"80732589",
X"38775279",
X"51782def",
X"39753375",
X"57537280",
X"2e903872",
X"52795178",
X"2d757081",
X"05573353",
X"ed398b3d",
X"0d04ee3d",
X"0d646669",
X"69707081",
X"0552335b",
X"4a5c5e5e",
X"76802e82",
X"f93876a5",
X"2e098106",
X"82e03880",
X"70416770",
X"70810552",
X"33714a59",
X"575f76b0",
X"2e098106",
X"8c387570",
X"81055733",
X"76485781",
X"5fd01756",
X"75892680",
X"da387667",
X"5c59805c",
X"9339778a",
X"2480c338",
X"7b8a2918",
X"7b708105",
X"5d335a5c",
X"d0197081",
X"ff065858",
X"897727a4",
X"38ff9f19",
X"7081ff06",
X"ffa91b5a",
X"51568576",
X"279238ff",
X"bf197081",
X"ff065156",
X"7585268a",
X"38c91958",
X"778025ff",
X"b9387a47",
X"7b407881",
X"ff065776",
X"80e42e80",
X"e5387680",
X"e424a738",
X"7680d82e",
X"81863876",
X"80d82490",
X"3876802e",
X"81cc3876",
X"a52e81b6",
X"3881b939",
X"7680e32e",
X"818c3881",
X"af397680",
X"f52e9b38",
X"7680f524",
X"8b387680",
X"f32e8181",
X"38819939",
X"7680f82e",
X"80ca3881",
X"8f39913d",
X"70555780",
X"538a5279",
X"841b7108",
X"535b56fb",
X"fd3f7655",
X"ab397984",
X"1b710894",
X"3d705b5b",
X"525b5675",
X"80258c38",
X"753056ad",
X"78340280",
X"c1055776",
X"5480538a",
X"527551fb",
X"d13f7755",
X"7e54b839",
X"913d7055",
X"7780d832",
X"70307080",
X"25565158",
X"56905279",
X"841b7108",
X"535b57fb",
X"ad3f7555",
X"db397984",
X"1b831233",
X"545b5698",
X"3979841b",
X"7108575b",
X"5680547f",
X"537c527d",
X"51fc9c3f",
X"87397652",
X"7d517c2d",
X"66703358",
X"810547fd",
X"8339943d",
X"0d047283",
X"e0900c71",
X"83e0940c",
X"04fb3d0d",
X"883d7070",
X"84055208",
X"57547553",
X"83e09008",
X"5283e094",
X"0851fcc6",
X"3f873d0d",
X"04ff3d0d",
X"73700853",
X"51029305",
X"33723470",
X"08810571",
X"0c833d0d",
X"04fc3d0d",
X"873d8811",
X"55785498",
X"f15351fc",
X"993f8052",
X"873d51d1",
X"3f863d0d",
X"04fd3d0d",
X"75705254",
X"a3c43f83",
X"e0800814",
X"5372742e",
X"9238ff13",
X"70335353",
X"71af2e09",
X"8106ee38",
X"81135372",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"77705354",
X"54c73f83",
X"e0800873",
X"2ea13883",
X"e0800873",
X"3152ff12",
X"5271ff2e",
X"8f387270",
X"81055433",
X"74708105",
X"5634eb39",
X"ff145480",
X"7434853d",
X"0d04803d",
X"0d7251ff",
X"903f823d",
X"0d047183",
X"e0800c04",
X"803d0d72",
X"51807134",
X"810bbc12",
X"0c800b80",
X"c0120c82",
X"3d0d0480",
X"0b83e2d4",
X"08248a38",
X"a4ae3fff",
X"0b83e2d4",
X"0c800b83",
X"e0800c04",
X"ff3d0d73",
X"5283e0b0",
X"08722e8d",
X"38d93f71",
X"5196993f",
X"7183e0b0",
X"0c833d0d",
X"04f43d0d",
X"7e60625c",
X"5a558154",
X"bc150881",
X"91387451",
X"cf3f7958",
X"807a2580",
X"f73883e3",
X"84087089",
X"2a5783ff",
X"06788480",
X"72315656",
X"57737825",
X"83387355",
X"7583e2d4",
X"082e8438",
X"ff893f83",
X"e2d40880",
X"25a63875",
X"892b5198",
X"dc3f83e3",
X"84088f3d",
X"fc11555c",
X"548152f8",
X"1b5196c6",
X"3f761483",
X"e3840c75",
X"83e2d40c",
X"74537652",
X"7851a2df",
X"3f83e080",
X"0883e384",
X"081683e3",
X"840c7876",
X"31761b5b",
X"59567780",
X"24ff8b38",
X"617a710c",
X"54755475",
X"802e8338",
X"81547383",
X"e0800c8e",
X"3d0d04fc",
X"3d0dfe9b",
X"3f7651fe",
X"af3f863d",
X"fc055378",
X"52775195",
X"e93f7975",
X"710c5483",
X"e0800854",
X"83e08008",
X"802e8338",
X"81547383",
X"e0800c86",
X"3d0d04fe",
X"3d0d7583",
X"e2d40853",
X"53807224",
X"89387173",
X"2e8438fd",
X"d63f7451",
X"fdea3f72",
X"5197ae3f",
X"83e08008",
X"5283e080",
X"08802e83",
X"38815271",
X"83e0800c",
X"843d0d04",
X"803d0d72",
X"80c01108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"72bc1108",
X"83e0800c",
X"51823d0d",
X"0480c40b",
X"83e0800c",
X"04fd3d0d",
X"75777154",
X"70535553",
X"9f9c3f82",
X"c81308bc",
X"150c82c0",
X"130880c0",
X"150cfceb",
X"3f735193",
X"ab3f7383",
X"e0b00c83",
X"e0800853",
X"83e08008",
X"802e8338",
X"81537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"5553fcbf",
X"3f72802e",
X"a538bc13",
X"08527351",
X"9ea63f83",
X"e080088f",
X"38775272",
X"51ff9a3f",
X"83e08008",
X"538a3982",
X"cc130853",
X"d8398153",
X"7283e080",
X"0c853d0d",
X"04fe3d0d",
X"ff0b83e2",
X"d40c7483",
X"e0b40c75",
X"83e2d00c",
X"9f933f83",
X"e0800881",
X"ff065281",
X"53719938",
X"83e2ec51",
X"8e943f83",
X"e0800852",
X"83e08008",
X"802e8338",
X"72527153",
X"7283e080",
X"0c843d0d",
X"04fa3d0d",
X"787a82c4",
X"120882c4",
X"12087072",
X"24595656",
X"57577373",
X"2e098106",
X"913880c0",
X"165280c0",
X"17519c97",
X"3f83e080",
X"08557483",
X"e0800c88",
X"3d0d04f6",
X"3d0d7c5b",
X"807b715c",
X"54577a77",
X"2e8c3881",
X"1a82cc14",
X"08545a72",
X"f6388059",
X"80d9397a",
X"54815780",
X"707b7b31",
X"5a5755ff",
X"18537473",
X"2580c138",
X"82cc1408",
X"527351ff",
X"8c3f800b",
X"83e08008",
X"25a13882",
X"cc140882",
X"cc110882",
X"cc160c74",
X"82cc120c",
X"5375802e",
X"86387282",
X"cc170c72",
X"54805773",
X"82cc1508",
X"81175755",
X"56ffb839",
X"81195980",
X"0bff1b54",
X"54787325",
X"83388154",
X"76813270",
X"75065153",
X"72ff9038",
X"8c3d0d04",
X"f73d0d7b",
X"7d5a5a82",
X"d05283e2",
X"d0085180",
X"d0b53f83",
X"e0800857",
X"f9e13f79",
X"5283e2d8",
X"5195b53f",
X"83e08008",
X"54805383",
X"e0800873",
X"2e098106",
X"82833883",
X"e0b4080b",
X"0b80f3e0",
X"53705256",
X"9bd43f0b",
X"0b80f3e0",
X"5280c016",
X"519bc73f",
X"75bc170c",
X"7382c017",
X"0c810b82",
X"c4170c81",
X"0b82c817",
X"0c7382cc",
X"170cff17",
X"82d01755",
X"57819139",
X"83e0c033",
X"70822a70",
X"81065154",
X"55728180",
X"3874812a",
X"81065877",
X"80f63874",
X"842a8106",
X"82c4150c",
X"83e0c033",
X"810682c8",
X"150c7952",
X"73519aee",
X"3f73519b",
X"853f83e0",
X"80081453",
X"af737081",
X"05553472",
X"bc150c83",
X"e0c15272",
X"519acf3f",
X"83e0b808",
X"82c0150c",
X"83e0ce52",
X"80c01451",
X"9abc3f78",
X"802e8d38",
X"7351782d",
X"83e08008",
X"802e9938",
X"7782cc15",
X"0c75802e",
X"86387382",
X"cc170c73",
X"82d015ff",
X"19595556",
X"76802e9b",
X"3883e0b8",
X"5283e2d8",
X"5194ab3f",
X"83e08008",
X"8a3883e0",
X"c1335372",
X"fed23878",
X"802e8938",
X"83e0b408",
X"51fcb83f",
X"83e0b408",
X"537283e0",
X"800c8b3d",
X"0d04ff3d",
X"0d805273",
X"51fdb53f",
X"833d0d04",
X"f03d0d62",
X"705254f6",
X"903f83e0",
X"80087453",
X"873d7053",
X"5555f6b0",
X"3ff7903f",
X"7351d33f",
X"63537452",
X"83e08008",
X"51fab83f",
X"923d0d04",
X"7183e080",
X"0c0480c0",
X"1283e080",
X"0c04803d",
X"0d7282c0",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"cc110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"82c41108",
X"83e0800c",
X"51823d0d",
X"04f93d0d",
X"7983e098",
X"08575781",
X"77278196",
X"38768817",
X"0827818e",
X"38753355",
X"74822e89",
X"3874832e",
X"b33880fe",
X"39745476",
X"1083fe06",
X"5376882a",
X"8c170805",
X"52893dfc",
X"055199c1",
X"3f83e080",
X"0880df38",
X"029d0533",
X"893d3371",
X"882b0756",
X"5680d139",
X"84547682",
X"2b83fc06",
X"5376872a",
X"8c170805",
X"52893dfc",
X"05519991",
X"3f83e080",
X"08b03802",
X"9f053302",
X"84059e05",
X"3371982b",
X"71902b07",
X"028c059d",
X"05337088",
X"2b72078d",
X"3d337180",
X"fffffe80",
X"06075152",
X"53575856",
X"83398155",
X"7483e080",
X"0c893d0d",
X"04fb3d0d",
X"83e09808",
X"fe198812",
X"08fe0555",
X"56548056",
X"7473278d",
X"38821433",
X"75712994",
X"16080557",
X"537583e0",
X"800c873d",
X"0d04fc3d",
X"0d765280",
X"0b83e098",
X"08703351",
X"52537083",
X"2e098106",
X"91389512",
X"33941333",
X"71982b71",
X"902b0755",
X"55519b12",
X"339a1333",
X"71882b07",
X"740783e0",
X"800c5586",
X"3d0d04fc",
X"3d0d7683",
X"e0980855",
X"55807523",
X"88150853",
X"72812e88",
X"38881408",
X"73268538",
X"8152b239",
X"72903873",
X"33527183",
X"2e098106",
X"85389014",
X"0853728c",
X"160c7280",
X"2e8d3872",
X"51fed63f",
X"83e08008",
X"52853990",
X"14085271",
X"90160c80",
X"527183e0",
X"800c863d",
X"0d04fa3d",
X"0d7883e0",
X"98087122",
X"81057083",
X"ffff0657",
X"54575573",
X"802e8838",
X"90150853",
X"72863883",
X"5280e739",
X"738f0652",
X"7180da38",
X"81139016",
X"0c8c1508",
X"53729038",
X"830b8417",
X"22575273",
X"762780c6",
X"38bf3982",
X"1633ff05",
X"74842a06",
X"5271b238",
X"7251fcb1",
X"3f815271",
X"83e08008",
X"27a83883",
X"5283e080",
X"08881708",
X"279c3883",
X"e080088c",
X"160c83e0",
X"800851fd",
X"bc3f83e0",
X"80089016",
X"0c737523",
X"80527183",
X"e0800c88",
X"3d0d04f2",
X"3d0d6062",
X"64585e5b",
X"75335574",
X"a02e0981",
X"06883881",
X"16704456",
X"ef396270",
X"33565674",
X"af2e0981",
X"06843881",
X"1643800b",
X"881c0c62",
X"70335155",
X"749f2691",
X"387a51fd",
X"d23f83e0",
X"80085680",
X"7d348381",
X"39933d84",
X"1c087058",
X"595f8a55",
X"a0767081",
X"055834ff",
X"155574ff",
X"2e098106",
X"ef388070",
X"5a5c887f",
X"085f5a7b",
X"811d7081",
X"ff066013",
X"703370af",
X"327030a0",
X"73277180",
X"25075151",
X"525b535e",
X"57557480",
X"e73876ae",
X"2e098106",
X"83388155",
X"787a2775",
X"07557480",
X"2e9f3879",
X"88327030",
X"78ae3270",
X"30707307",
X"9f2a5351",
X"57515675",
X"bb388859",
X"8b5affab",
X"3976982b",
X"55748025",
X"873880f1",
X"b4173357",
X"ff9f1755",
X"74992689",
X"38e01770",
X"81ff0658",
X"5578811a",
X"7081ff06",
X"721b535b",
X"57557675",
X"34fef839",
X"7b1e7f0c",
X"805576a0",
X"26833881",
X"55748b19",
X"347a51fc",
X"823f83e0",
X"800880f5",
X"38a0547a",
X"2270852b",
X"83e00654",
X"55901b08",
X"527c5193",
X"cc3f83e0",
X"80085783",
X"e0800881",
X"81387c33",
X"5574802e",
X"80f4388b",
X"1d337083",
X"2a708106",
X"51565674",
X"b4388b7d",
X"841d0883",
X"e0800859",
X"5b5b58ff",
X"185877ff",
X"2e9a3879",
X"7081055b",
X"33797081",
X"055b3371",
X"71315256",
X"5675802e",
X"e2388639",
X"75802e96",
X"387a51fb",
X"e53fff86",
X"3983e080",
X"085683e0",
X"8008b638",
X"83397656",
X"841b088b",
X"11335155",
X"74a7388b",
X"1d337084",
X"2a708106",
X"51565674",
X"89388356",
X"94398156",
X"90397c51",
X"fa943f83",
X"e0800888",
X"1c0cfd81",
X"397583e0",
X"800c903d",
X"0d04f83d",
X"0d7a7c59",
X"57825483",
X"fe537752",
X"76519291",
X"3f835683",
X"e0800880",
X"ec388117",
X"33773371",
X"882b0756",
X"56825674",
X"82d4d52e",
X"09810680",
X"d4387554",
X"b6537752",
X"765191e5",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"ac388254",
X"80d25377",
X"52765191",
X"bc3f83e0",
X"80089838",
X"81173377",
X"3371882b",
X"0783e080",
X"08525656",
X"748182c6",
X"2e833881",
X"567583e0",
X"800c8a3d",
X"0d04eb3d",
X"0d675a80",
X"0b83e098",
X"0c90de3f",
X"83e08008",
X"81065582",
X"567483ef",
X"38747553",
X"8f3d7053",
X"5759feca",
X"3f83e080",
X"0881ff06",
X"5776812e",
X"09810680",
X"d4389054",
X"83be5374",
X"52755190",
X"d03f83e0",
X"800880c9",
X"388f3d33",
X"5574802e",
X"80c93802",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"70587b57",
X"5e525e57",
X"5957fdee",
X"3f83e080",
X"0881ff06",
X"5776832e",
X"09810686",
X"38815682",
X"f2397680",
X"2e863886",
X"5682e839",
X"a4548d53",
X"78527551",
X"8fe73f81",
X"5683e080",
X"0882d438",
X"02be0533",
X"028405bd",
X"05337188",
X"2b07595d",
X"77ab3802",
X"80ce0533",
X"02840580",
X"cd053371",
X"982b7190",
X"2b07973d",
X"3370882b",
X"72070294",
X"0580cb05",
X"33710754",
X"525e5759",
X"5602b705",
X"33787129",
X"028805b6",
X"0533028c",
X"05b50533",
X"71882b07",
X"701d707f",
X"8c050c5f",
X"5957595d",
X"8e3d3382",
X"1b3402b9",
X"0533903d",
X"3371882b",
X"075a5c78",
X"841b2302",
X"bb053302",
X"8405ba05",
X"3371882b",
X"07565c74",
X"ab380280",
X"ca053302",
X"840580c9",
X"05337198",
X"2b71902b",
X"07963d33",
X"70882b72",
X"07029405",
X"80c70533",
X"71075152",
X"53575e5c",
X"74763178",
X"3179842a",
X"903d3354",
X"71713153",
X"565680c1",
X"9a3f83e0",
X"80088205",
X"70881c0c",
X"83e08008",
X"e08a0556",
X"567483df",
X"fe268338",
X"825783ff",
X"f6762785",
X"38835789",
X"39865676",
X"802e80db",
X"38767a34",
X"76832e09",
X"8106b038",
X"0280d605",
X"33028405",
X"80d50533",
X"71982b71",
X"902b0799",
X"3d337088",
X"2b720702",
X"940580d3",
X"05337107",
X"7f90050c",
X"525e5758",
X"56863977",
X"1b901b0c",
X"841a228c",
X"1b081971",
X"842a0594",
X"1c0c5d80",
X"0b811b34",
X"7983e098",
X"0c805675",
X"83e0800c",
X"973d0d04",
X"e93d0d83",
X"e0980856",
X"85547580",
X"2e818238",
X"800b8117",
X"34993de0",
X"11466a54",
X"8a3d7054",
X"58ec0551",
X"f6e53f83",
X"e0800854",
X"83e08008",
X"80df3889",
X"3d335473",
X"802e9138",
X"02ab0533",
X"70842a81",
X"06515574",
X"802e8638",
X"835480c1",
X"397651f4",
X"893f83e0",
X"8008a017",
X"0c02bf05",
X"33028405",
X"be053371",
X"982b7190",
X"2b07028c",
X"05bd0533",
X"70882b72",
X"07953d33",
X"71079c1c",
X"0c527898",
X"1b0c5356",
X"5957810b",
X"81173474",
X"547383e0",
X"800c993d",
X"0d04f53d",
X"0d7d7f61",
X"7283e098",
X"085a5d5d",
X"595c807b",
X"0c855775",
X"802e81e0",
X"38811633",
X"81065584",
X"5774802e",
X"81d23891",
X"39748117",
X"34863980",
X"0b811734",
X"815781c0",
X"399c1608",
X"98170831",
X"55747827",
X"83387458",
X"77802e81",
X"a9389816",
X"087083ff",
X"06565774",
X"80cf3882",
X"1633ff05",
X"77892a06",
X"7081ff06",
X"5a5578a0",
X"38768738",
X"a0160855",
X"8d39a416",
X"0851f0e9",
X"3f83e080",
X"08558175",
X"27ffa838",
X"74a4170c",
X"a4160851",
X"f2833f83",
X"e0800855",
X"83e08008",
X"802eff89",
X"3883e080",
X"0819a817",
X"0c981608",
X"83ff0684",
X"80713151",
X"55777527",
X"83387755",
X"7483ffff",
X"06549816",
X"0883ff06",
X"53a81608",
X"5279577b",
X"83387b57",
X"76518a8d",
X"3f83e080",
X"08fed038",
X"98160815",
X"98170c74",
X"1a787631",
X"7c08177d",
X"0c595afe",
X"d3398057",
X"7683e080",
X"0c8d3d0d",
X"04fa3d0d",
X"7883e098",
X"08555685",
X"5573802e",
X"81e13881",
X"14338106",
X"53845572",
X"802e81d3",
X"389c1408",
X"53727627",
X"83387256",
X"98140857",
X"800b9815",
X"0c75802e",
X"81b73882",
X"14337089",
X"2b565376",
X"802eb538",
X"7452ff16",
X"51bc9c3f",
X"83e08008",
X"ff187654",
X"70535853",
X"bc8d3f83",
X"e0800873",
X"26963874",
X"30707806",
X"7098170c",
X"777131a4",
X"17085258",
X"51538939",
X"a0140870",
X"a4160c53",
X"747627b9",
X"387251ee",
X"d83f83e0",
X"80085381",
X"0b83e080",
X"08278b38",
X"88140883",
X"e0800826",
X"8838800b",
X"811534b0",
X"3983e080",
X"08a4150c",
X"98140815",
X"98150c75",
X"753156c4",
X"39981408",
X"16709816",
X"0c735256",
X"efc73f83",
X"e080088c",
X"3883e080",
X"08811534",
X"81559439",
X"821433ff",
X"0576892a",
X"0683e080",
X"0805a815",
X"0c805574",
X"83e0800c",
X"883d0d04",
X"ef3d0d63",
X"56855583",
X"e0980880",
X"2e80d238",
X"933df405",
X"84170c64",
X"53883d70",
X"53765257",
X"f1d13f83",
X"e0800855",
X"83e08008",
X"b438883d",
X"33547380",
X"2ea13802",
X"a7053370",
X"842a7081",
X"06515555",
X"83557380",
X"2e973876",
X"51eef73f",
X"83e08008",
X"88170c75",
X"51efa83f",
X"83e08008",
X"557483e0",
X"800c933d",
X"0d04e43d",
X"0d6ea13d",
X"08405e85",
X"5683e098",
X"08802e84",
X"85389e3d",
X"f405841f",
X"0c7e9838",
X"7d51eef7",
X"3f83e080",
X"085683ee",
X"39814181",
X"f6398341",
X"81f13993",
X"3d7f9605",
X"4159807f",
X"8295055e",
X"56756081",
X"ff053483",
X"41901e08",
X"762e81d3",
X"38a0547d",
X"2270852b",
X"83e00654",
X"58901e08",
X"52785186",
X"983f83e0",
X"80084183",
X"e08008ff",
X"b8387833",
X"5c7b802e",
X"ffb4388b",
X"193370bf",
X"06718106",
X"52435574",
X"802e80de",
X"387b81bf",
X"0655748f",
X"2480d338",
X"9a193355",
X"7480cb38",
X"f31d7058",
X"5d815675",
X"8b2e0981",
X"0685388e",
X"568b3975",
X"9a2e0981",
X"0683389c",
X"56751970",
X"70810552",
X"33713381",
X"1a821a5f",
X"5b525b55",
X"74863879",
X"77348539",
X"80df7734",
X"777b5757",
X"7aa02e09",
X"8106c038",
X"81567b81",
X"e5327030",
X"709f2a51",
X"51557bae",
X"2e933874",
X"802e8e38",
X"61832a70",
X"81065155",
X"74802e97",
X"387d51ed",
X"e13f83e0",
X"80084183",
X"e0800887",
X"38901e08",
X"feaf3880",
X"60347580",
X"2e88387c",
X"527f5183",
X"a53f6080",
X"2e863880",
X"0b901f0c",
X"60566083",
X"2e853860",
X"81d03889",
X"1f57901e",
X"08802e81",
X"a8388056",
X"75197033",
X"515574a0",
X"2ea03874",
X"852e0981",
X"06843881",
X"e5557477",
X"70810559",
X"34811670",
X"81ff0657",
X"55877627",
X"d7388819",
X"335574a0",
X"2ea938ae",
X"77708105",
X"59348856",
X"75197033",
X"515574a0",
X"2e953874",
X"77708105",
X"59348116",
X"7081ff06",
X"57558a76",
X"27e2388b",
X"19337f88",
X"05349f19",
X"339e1a33",
X"71982b71",
X"902b079d",
X"1c337088",
X"2b72079c",
X"1e337107",
X"640c5299",
X"1d33981e",
X"3371882b",
X"07535153",
X"57595674",
X"7f840523",
X"97193396",
X"1a337188",
X"2b075656",
X"747f8605",
X"23807734",
X"7d51ebf2",
X"3f83e080",
X"08833270",
X"30707207",
X"9f2c83e0",
X"80080652",
X"5656961f",
X"3355748a",
X"38891f52",
X"961f5181",
X"b13f7583",
X"e0800c9e",
X"3d0d04fd",
X"3d0d7577",
X"53547333",
X"51708938",
X"71335170",
X"802ea138",
X"73337233",
X"52537271",
X"278538ff",
X"51943970",
X"73278538",
X"81518b39",
X"81148113",
X"5354d339",
X"80517083",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"54547233",
X"7081ff06",
X"52527080",
X"2ea33871",
X"81ff0681",
X"14ffbf12",
X"53545270",
X"99268938",
X"a0127081",
X"ff065351",
X"71747081",
X"055634d2",
X"39807434",
X"853d0d04",
X"ffbd3d0d",
X"80c63d08",
X"52a53d70",
X"5254ffb3",
X"3f80c73d",
X"0852853d",
X"705253ff",
X"a63f7252",
X"7351fedf",
X"3f80c53d",
X"0d04fe3d",
X"0d747653",
X"53717081",
X"05533351",
X"70737081",
X"05553470",
X"f038843d",
X"0d04fe3d",
X"0d745280",
X"72335253",
X"70732e8d",
X"38811281",
X"14713353",
X"545270f5",
X"387283e0",
X"800c843d",
X"0d04fc3d",
X"0d765574",
X"83e39808",
X"2eaf3880",
X"53745187",
X"c13f83e0",
X"800881ff",
X"06ff1470",
X"81ff0672",
X"30709f2a",
X"51525553",
X"5472802e",
X"843871dd",
X"3873fe38",
X"7483e398",
X"0c863d0d",
X"04ff3d0d",
X"ff0b83e3",
X"980c84a5",
X"3f815187",
X"853f83e0",
X"800881ff",
X"065271ee",
X"3881d33f",
X"7183e080",
X"0c833d0d",
X"04fc3d0d",
X"76028405",
X"a2052202",
X"8805a605",
X"227a5455",
X"5555ff82",
X"3f72802e",
X"a03883e3",
X"ac143375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552dd",
X"39800b83",
X"e0800c86",
X"3d0d04fc",
X"3d0d7678",
X"7a115653",
X"55805371",
X"742e9338",
X"72155170",
X"3383e3ac",
X"13348112",
X"81145452",
X"ea39800b",
X"83e0800c",
X"863d0d04",
X"fd3d0d90",
X"5483e398",
X"085186f4",
X"3f83e080",
X"0881ff06",
X"ff157130",
X"71307073",
X"079f2a72",
X"9f2a0652",
X"55525553",
X"72db3885",
X"3d0d0480",
X"3d0d83e3",
X"a4081083",
X"e39c0807",
X"9080a80c",
X"823d0d04",
X"800b83e3",
X"a40ce43f",
X"04810b83",
X"e3a40cdb",
X"3f04ed3f",
X"047183e3",
X"a00c0480",
X"3d0d8051",
X"f43f810b",
X"83e3a40c",
X"810b83e3",
X"9c0cffbb",
X"3f823d0d",
X"04803d0d",
X"72307074",
X"07802583",
X"e39c0c51",
X"ffa53f82",
X"3d0d0480",
X"3d0d028b",
X"05339080",
X"a40c9080",
X"a8087081",
X"06515170",
X"f5389080",
X"a4087081",
X"ff0683e0",
X"800c5182",
X"3d0d0480",
X"3d0d81ff",
X"51d13f83",
X"e0800881",
X"ff0683e0",
X"800c823d",
X"0d04803d",
X"0d73902b",
X"73079080",
X"b40c823d",
X"0d0404fb",
X"3d0d7802",
X"84059f05",
X"3370982b",
X"55575572",
X"80259b38",
X"7580ff06",
X"56805280",
X"f751e03f",
X"83e08008",
X"81ff0654",
X"73812680",
X"ff388051",
X"fee73fff",
X"a23f8151",
X"fedf3fff",
X"9a3f7551",
X"feed3f74",
X"982a51fe",
X"e63f7490",
X"2a7081ff",
X"065253fe",
X"da3f7488",
X"2a7081ff",
X"065253fe",
X"ce3f7481",
X"ff0651fe",
X"c63f8155",
X"7580c02e",
X"09810686",
X"38819555",
X"8d397580",
X"c82e0981",
X"06843881",
X"87557451",
X"fea53f8a",
X"55fec83f",
X"83e08008",
X"81ff0670",
X"982b5454",
X"7280258c",
X"38ff1570",
X"81ff0656",
X"5374e238",
X"7383e080",
X"0c873d0d",
X"04fa3d0d",
X"fdc53f80",
X"51fdda3f",
X"8a54fe93",
X"3fff1470",
X"81ff0655",
X"5373f338",
X"73745355",
X"80c051fe",
X"a63f83e0",
X"800881ff",
X"06547381",
X"2e098106",
X"829f3883",
X"aa5280c8",
X"51fe8c3f",
X"83e08008",
X"81ff0653",
X"72812e09",
X"810681a8",
X"38745487",
X"3d741154",
X"56fdc83f",
X"83e08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e53802",
X"9a053353",
X"72812e09",
X"810681d9",
X"38029b05",
X"335380ce",
X"90547281",
X"aa2e8d38",
X"81c73980",
X"e4518acc",
X"3fff1454",
X"73802e81",
X"b838820a",
X"5281e951",
X"fda53f83",
X"e0800881",
X"ff065372",
X"de387252",
X"80fa51fd",
X"923f83e0",
X"800881ff",
X"06537281",
X"90387254",
X"731653fc",
X"d63f83e0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e8",
X"38873d33",
X"70862a70",
X"81065154",
X"548c5572",
X"80e33884",
X"5580de39",
X"745281e9",
X"51fccc3f",
X"83e08008",
X"81ff0653",
X"825581e9",
X"56817327",
X"86387355",
X"80c15680",
X"ce90548a",
X"3980e451",
X"89be3fff",
X"14547380",
X"2ea93880",
X"527551fc",
X"9a3f83e0",
X"800881ff",
X"065372e1",
X"38848052",
X"80d051fc",
X"863f83e0",
X"800881ff",
X"06537280",
X"2e833880",
X"557483e3",
X"a8348051",
X"fb873ffb",
X"c23f883d",
X"0d04fb3d",
X"0d775480",
X"0b83e3a8",
X"3370832a",
X"70810651",
X"55575572",
X"752e0981",
X"06853873",
X"892b5473",
X"5280d151",
X"fbbd3f83",
X"e0800881",
X"ff065372",
X"bd3882b8",
X"c054fb83",
X"3f83e080",
X"0881ff06",
X"537281ff",
X"2e098106",
X"8938ff14",
X"5473e738",
X"9f397281",
X"fe2e0981",
X"06963883",
X"e7ac5283",
X"e3ac51fa",
X"ed3ffad3",
X"3ffad03f",
X"83398155",
X"8051fa89",
X"3ffac43f",
X"7481ff06",
X"83e0800c",
X"873d0d04",
X"fb3d0d77",
X"83e3ac56",
X"548151f9",
X"ec3f83e3",
X"a8337083",
X"2a708106",
X"51545672",
X"85387389",
X"2b547352",
X"80d851fa",
X"b63f83e0",
X"800881ff",
X"06537280",
X"e43881ff",
X"51f9d43f",
X"81fe51f9",
X"ce3f8480",
X"53747081",
X"05563351",
X"f9c13fff",
X"137083ff",
X"ff065153",
X"72eb3872",
X"51f9b03f",
X"7251f9ab",
X"3ff9d03f",
X"83e08008",
X"9f0653a7",
X"88547285",
X"2e8c3899",
X"3980e451",
X"86f63fff",
X"1454f9b3",
X"3f83e080",
X"0881ff2e",
X"843873e9",
X"388051f8",
X"e43ff99f",
X"3f800b83",
X"e0800c87",
X"3d0d0471",
X"83e7b00c",
X"8880800b",
X"83e7ac0c",
X"8480800b",
X"83e7b40c",
X"04fd3d0d",
X"77701755",
X"7705ff1a",
X"535371ff",
X"2e943873",
X"70810555",
X"33517073",
X"70810555",
X"34ff1252",
X"e939853d",
X"0d04fc3d",
X"0d87a681",
X"55743383",
X"e7b834a0",
X"5483a080",
X"5383e7b0",
X"085283e7",
X"ac0851ff",
X"b83fa054",
X"83a48053",
X"83e7b008",
X"5283e7ac",
X"0851ffa5",
X"3f905483",
X"a8805383",
X"e7b00852",
X"83e7ac08",
X"51ff923f",
X"a0538052",
X"83e7b408",
X"83a08005",
X"5185ce3f",
X"a0538052",
X"83e7b408",
X"83a48005",
X"5185be3f",
X"90538052",
X"83e7b408",
X"83a88005",
X"5185ae3f",
X"ff753483",
X"a0805480",
X"5383e7b0",
X"085283e7",
X"b40851fe",
X"cc3f80d0",
X"805483b0",
X"805383e7",
X"b0085283",
X"e7b40851",
X"feb73f86",
X"e13fa254",
X"805383e7",
X"b4088c80",
X"055280f6",
X"d851fea1",
X"3f860b87",
X"a8833480",
X"0b87a882",
X"34800b87",
X"a09a34af",
X"0b87a096",
X"34bf0b87",
X"a0973480",
X"0b87a098",
X"349f0b87",
X"a0993480",
X"0b87a09b",
X"34e00b87",
X"a88934a2",
X"0b87a880",
X"34830b87",
X"a48f3482",
X"0b87a881",
X"34863d0d",
X"04fd3d0d",
X"83a08054",
X"805383e7",
X"b4085283",
X"e7b00851",
X"fdbf3f80",
X"d0805483",
X"b0805383",
X"e7b40852",
X"83e7b008",
X"51fdaa3f",
X"a05483a0",
X"805383e7",
X"b4085283",
X"e7b00851",
X"fd973fa0",
X"5483a480",
X"5383e7b4",
X"085283e7",
X"b00851fd",
X"843f9054",
X"83a88053",
X"83e7b408",
X"5283e7b0",
X"0851fcf1",
X"3f83e7b8",
X"3387a681",
X"34853d0d",
X"04803d0d",
X"90809008",
X"810683e0",
X"800c823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087081",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fd0676",
X"1007720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870822c",
X"bf0683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe830676",
X"822b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087088",
X"2c870683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f1ff06",
X"76882b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"8b2cbf06",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f88f",
X"ff06768b",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870912c",
X"bf0683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fc87ffff",
X"0676912b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70992c81",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870ff",
X"bf0a0676",
X"992b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"80087088",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"892c8106",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708a2c81",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708b2c",
X"810683e0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708c",
X"2cbf0683",
X"e0800c51",
X"823d0d04",
X"fe3d0d74",
X"81e62987",
X"2a9080a0",
X"0c843d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727081",
X"055434ff",
X"1151f039",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708405",
X"540cff11",
X"51f03984",
X"3d0d04fe",
X"3d0d8480",
X"80538052",
X"88800a51",
X"ffb33f81",
X"80805380",
X"5282800a",
X"51c63f84",
X"3d0d0480",
X"3d0d8151",
X"fbfc3f72",
X"802e9038",
X"8051fdfe",
X"3fcd3f83",
X"e7bc3351",
X"fdf43f81",
X"51fc8d3f",
X"8051fc88",
X"3f8051fb",
X"d93f823d",
X"0d04fd3d",
X"0d755280",
X"5480ff72",
X"25883881",
X"0bff8013",
X"5354ffbf",
X"12517099",
X"268638e0",
X"12529e39",
X"ff9f1251",
X"99712795",
X"38d012e0",
X"13705454",
X"51897127",
X"88388f73",
X"27833880",
X"5273802e",
X"85388180",
X"12527181",
X"ff0683e0",
X"800c853d",
X"0d04803d",
X"0d84d8c0",
X"51807170",
X"81055334",
X"7084e0c0",
X"2e098106",
X"f038823d",
X"0d04fe3d",
X"0d029705",
X"3351ff86",
X"3f83e080",
X"0881ff06",
X"83e7c008",
X"54528073",
X"249b3883",
X"e7e00813",
X"7283e7e4",
X"08075353",
X"71733483",
X"e7c00881",
X"0583e7c0",
X"0c843d0d",
X"04fa3d0d",
X"82800a1b",
X"55805788",
X"3dfc0554",
X"79537452",
X"7851cbd3",
X"3f883d0d",
X"04fe3d0d",
X"83e7d808",
X"527451d2",
X"b73f83e0",
X"80088c38",
X"76537552",
X"83e7d808",
X"51c73f84",
X"3d0d04fe",
X"3d0d83e7",
X"d8085375",
X"527451cc",
X"f63f83e0",
X"80088d38",
X"77537652",
X"83e7d808",
X"51ffa23f",
X"843d0d04",
X"fe3d0d83",
X"e7d80851",
X"cbea3f83",
X"e0800881",
X"80802e09",
X"81068738",
X"b1808053",
X"9a3983e7",
X"d80851cb",
X"cf3f83e0",
X"800880d0",
X"802e0981",
X"069238b1",
X"b0805383",
X"e0800852",
X"83e7d808",
X"51feda3f",
X"843d0d04",
X"803d0df9",
X"e63f83e0",
X"80088429",
X"80f6fc05",
X"700883e0",
X"800c5182",
X"3d0d04ed",
X"3d0d8043",
X"80428041",
X"80705a5b",
X"fdd43f80",
X"0b83e7c0",
X"0c800b83",
X"e7e40c80",
X"f4d851c6",
X"bc3f8180",
X"0b83e7e4",
X"0c80f4dc",
X"51c6ae3f",
X"80d00b83",
X"e7c00c78",
X"30707a07",
X"80257087",
X"2b83e7e4",
X"0c5155f8",
X"d93f83e0",
X"80085280",
X"f4e451c6",
X"883f80f8",
X"0b83e7c0",
X"0c788132",
X"70307072",
X"07802570",
X"872b83e7",
X"e40c5156",
X"56fef13f",
X"83e08008",
X"5280f4f0",
X"51c5de3f",
X"81a00b83",
X"e7c00c78",
X"82327030",
X"70720780",
X"2570872b",
X"83e7e40c",
X"515683e7",
X"d8085256",
X"c6f83f83",
X"e0800852",
X"80f4f851",
X"c5af3f81",
X"f00b83e7",
X"c00c810b",
X"83e7c45b",
X"5883e7c0",
X"0882197a",
X"32703070",
X"72078025",
X"70872b83",
X"e7e40c51",
X"578e3d70",
X"55ff1b54",
X"57575799",
X"bf3f7970",
X"84055b08",
X"51c6af3f",
X"745483e0",
X"80085377",
X"5280f580",
X"51c4e23f",
X"a81783e7",
X"c00c8118",
X"5877852e",
X"098106ff",
X"b0388390",
X"0b83e7c0",
X"0c788732",
X"70307072",
X"07802570",
X"872b83e7",
X"e40c5156",
X"56f7ff3f",
X"80f59055",
X"83e08008",
X"802e8e38",
X"83e7d408",
X"51c5db3f",
X"83e08008",
X"55745280",
X"f59851c4",
X"903f83e0",
X"0b83e7c0",
X"0c788832",
X"70307072",
X"07802570",
X"872b83e7",
X"e40c5157",
X"80f5a452",
X"55c3ee3f",
X"868da051",
X"f8fa3f80",
X"52913d70",
X"52559ae3",
X"3f835274",
X"519adc3f",
X"63557482",
X"fc386119",
X"59788025",
X"85387459",
X"90398879",
X"25853888",
X"59873978",
X"882682db",
X"3878822b",
X"5580f3b4",
X"150804f5",
X"ed3f83e0",
X"80086157",
X"5575812e",
X"09810689",
X"3883e080",
X"08105590",
X"3975ff2e",
X"09810688",
X"3883e080",
X"08812c55",
X"90752585",
X"38905588",
X"39748024",
X"83388155",
X"7451f5c7",
X"3f829039",
X"f5d93f83",
X"e0800861",
X"05557480",
X"25853880",
X"55883987",
X"75258338",
X"87557451",
X"f5d23f81",
X"ee396087",
X"3862802e",
X"81e53883",
X"e0a40883",
X"e0a00c8a",
X"ea0b83e0",
X"a80c83e7",
X"d80851ff",
X"b4f23ffa",
X"e33f81c7",
X"39605680",
X"76259938",
X"8a830b83",
X"e0a80c83",
X"e7b81570",
X"085255ff",
X"b4d23f74",
X"08529139",
X"75802591",
X"3883e7b8",
X"150851c3",
X"c33f8052",
X"fd1951b8",
X"3962802e",
X"818d3883",
X"e7b81570",
X"0883e7c4",
X"08720c83",
X"e7c40cfd",
X"1a705351",
X"558ba93f",
X"83e08008",
X"5680518b",
X"9f3f83e0",
X"80085274",
X"5187b73f",
X"75528051",
X"87b03f80",
X"d6396055",
X"807525b8",
X"3883e0ac",
X"0883e0a0",
X"0c8aea0b",
X"83e0a80c",
X"83e7d408",
X"51ffb3dc",
X"3f83e7d4",
X"0851ffb1",
X"eb3f83e0",
X"800881ff",
X"06705255",
X"f4dd3f74",
X"802e9c38",
X"8155a039",
X"74802593",
X"3883e7d4",
X"0851c2b4",
X"3f8051f4",
X"c23f8439",
X"6287387a",
X"802efa84",
X"38805574",
X"83e0800c",
X"953d0d04",
X"fe3d0df4",
X"ee3f83e0",
X"8008802e",
X"86388051",
X"818b39f4",
X"f33f83e0",
X"800880ff",
X"38f5933f",
X"83e08008",
X"802eb938",
X"8151f2a2",
X"3f8051f4",
X"a93fef96",
X"3f800b83",
X"e7c00cf9",
X"ae3f83e0",
X"800853ff",
X"0b83e7c0",
X"0cf1823f",
X"7280cc38",
X"83e7bc33",
X"51f4833f",
X"7251f1f2",
X"3f80c139",
X"f4bb3f83",
X"e0800880",
X"2eb63881",
X"51f1df3f",
X"8051f3e6",
X"3feed33f",
X"8a830b83",
X"e0a80c83",
X"e7c40851",
X"ffb28d3f",
X"ff0b83e7",
X"c00cf0bd",
X"3f83e7c4",
X"08528051",
X"85ac3f81",
X"51f5ac3f",
X"843d0d04",
X"fc3d0d80",
X"0b83e7bc",
X"34848080",
X"5284a480",
X"8051c4ed",
X"3f83e080",
X"0880cb38",
X"88f73f80",
X"f8d051c9",
X"ad3f83e0",
X"800855b0",
X"80805480",
X"c0805380",
X"f5ac5283",
X"e0800851",
X"f7813f83",
X"e7d80853",
X"80f5bc52",
X"7451c3f7",
X"3f83e080",
X"088438f7",
X"8f3f83e7",
X"bc3351f2",
X"d93f8151",
X"f4c53f92",
X"fb3f8151",
X"f4bd3ffd",
X"ef3ffc39",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"0280f5c8",
X"0b83e0a4",
X"0c80f5cc",
X"0b83e09c",
X"0c80f5d0",
X"0b83e0ac",
X"0c83e08c",
X"08fc050c",
X"800b83e7",
X"c40b83e0",
X"8c08f805",
X"0c83e08c",
X"08f4050c",
X"c2c73f83",
X"e0800886",
X"05fc0683",
X"e08c08f0",
X"050c0283",
X"e08c08f0",
X"0508310d",
X"833d7083",
X"e08c08f8",
X"05087084",
X"0583e08c",
X"08f8050c",
X"0c51ffbf",
X"8f3f83e0",
X"8c08f405",
X"08810583",
X"e08c08f4",
X"050c83e0",
X"8c08f405",
X"08872e09",
X"8106ffac",
X"3884a880",
X"8051ebdb",
X"3fff0b83",
X"e7c00c80",
X"0b83e7e4",
X"0c84d8c0",
X"0b83e7e0",
X"0c8151ef",
X"853f8151",
X"efaa3f80",
X"51efa53f",
X"8151efcb",
X"3f8151f0",
X"a03f8251",
X"efee3f80",
X"51f0c43f",
X"8051f0ee",
X"3f80cff2",
X"528051ff",
X"bcc83ffd",
X"ab3f83e0",
X"8c08fc05",
X"080d800b",
X"83e0800c",
X"873d0d83",
X"e08c0c04",
X"803d0d81",
X"ff51800b",
X"83e7f012",
X"34ff1151",
X"70f43882",
X"3d0d04ff",
X"3d0d7370",
X"33535181",
X"11337134",
X"71811234",
X"833d0d04",
X"fb3d0d77",
X"79565680",
X"70715555",
X"52717525",
X"ac387216",
X"70337014",
X"7081ff06",
X"55515151",
X"71742789",
X"38811270",
X"81ff0653",
X"51718114",
X"7083ffff",
X"06555254",
X"747324d6",
X"387183e0",
X"800c873d",
X"0d04fc3d",
X"0d7655ff",
X"b5f43f83",
X"e0800880",
X"2ef53883",
X"ea8c0886",
X"057081ff",
X"065253ff",
X"b3f43f84",
X"39fad93f",
X"ffb5d33f",
X"83e08008",
X"812ef238",
X"80547315",
X"53ffb4b9",
X"3f83e080",
X"08733481",
X"14547385",
X"2e098106",
X"e9388439",
X"faae3fff",
X"b5a83f83",
X"e0800880",
X"2ef23874",
X"3383e7f0",
X"34811533",
X"83e7f134",
X"82153383",
X"e7f23483",
X"153383e7",
X"f3348452",
X"83e7f051",
X"feba3f83",
X"e0800881",
X"ff068416",
X"33565372",
X"752e0981",
X"068d38ff",
X"b49d3f83",
X"e0800880",
X"2e9a3883",
X"ea8c08a8",
X"2e098106",
X"8938860b",
X"83ea8c0c",
X"8739a80b",
X"83ea8c0c",
X"80e451ef",
X"9b3f863d",
X"0d04f43d",
X"0d7e6059",
X"55805d80",
X"75822b71",
X"83ea9012",
X"0c83eaa4",
X"175b5b57",
X"76793477",
X"772e83b8",
X"38765277",
X"51ffbdd3",
X"3f8e3dfc",
X"05549053",
X"83e9f852",
X"7751ffbd",
X"8e3f7c56",
X"75902e09",
X"81068394",
X"3883e9f8",
X"51fd943f",
X"83e9fa51",
X"fd8d3f83",
X"e9fc51fd",
X"863f7683",
X"ea880c77",
X"51ffbada",
X"3f80f3e8",
X"5283e080",
X"0851ffaa",
X"803f83e0",
X"8008812e",
X"09810680",
X"d4387683",
X"eaa00c82",
X"0b83e9f8",
X"34ff960b",
X"83e9f934",
X"7751ffbd",
X"9f3f83e0",
X"80085583",
X"e0800877",
X"25883883",
X"e080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583e9fa",
X"347483e9",
X"fb347683",
X"e9fc34ff",
X"800b83e9",
X"fd348190",
X"3983e9f8",
X"3383e9f9",
X"3371882b",
X"07565b74",
X"83ffff2e",
X"09810680",
X"e838fe80",
X"0b83eaa0",
X"0c810b83",
X"ea880cff",
X"0b83e9f8",
X"34ff0b83",
X"e9f93477",
X"51ffbcac",
X"3f83e080",
X"0883eaa8",
X"0c83e080",
X"085583e0",
X"80088025",
X"883883e0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83e9fa34",
X"7483e9fb",
X"347683e9",
X"fc34ff80",
X"0b83e9fd",
X"34810b83",
X"ea8734a5",
X"39748596",
X"2e098106",
X"80fe3875",
X"83eaa00c",
X"7751ffbb",
X"e03f83ea",
X"873383e0",
X"80080755",
X"7483ea87",
X"3483ea87",
X"33810655",
X"74802e83",
X"38845783",
X"e9fc3383",
X"e9fd3371",
X"882b0756",
X"5c748180",
X"2e098106",
X"a13883e9",
X"fa3383e9",
X"fb337188",
X"2b07565b",
X"ad807527",
X"87387682",
X"07579c39",
X"76810757",
X"96397482",
X"802e0981",
X"06873876",
X"83075787",
X"397481ff",
X"268a3877",
X"83ea901b",
X"0c767934",
X"8e3d0d04",
X"803d0d72",
X"842983ea",
X"90057008",
X"83e0800c",
X"51823d0d",
X"04fe3d0d",
X"800b83e9",
X"f40c800b",
X"83e9f00c",
X"ff0b83e7",
X"ec0ca80b",
X"83ea8c0c",
X"ae51ffae",
X"bd3f800b",
X"83ea9054",
X"52807370",
X"8405550c",
X"81125271",
X"842e0981",
X"06ef3884",
X"3d0d04fe",
X"3d0d7402",
X"84059605",
X"22535371",
X"802e9738",
X"72708105",
X"543351ff",
X"aec73fff",
X"127083ff",
X"ff065152",
X"e639843d",
X"0d04fe3d",
X"0d029205",
X"225382ac",
X"51eaad3f",
X"80c351ff",
X"aea33f81",
X"9651eaa0",
X"3f725283",
X"e7f051ff",
X"b23f7252",
X"83e7f051",
X"f8ee3f83",
X"e0800881",
X"ff0651ff",
X"adff3f84",
X"3d0d04ff",
X"b13d0d80",
X"d13df805",
X"51f9973f",
X"83e9f408",
X"810583e9",
X"f40c80cf",
X"3d33cf11",
X"7081ff06",
X"51565674",
X"832688ed",
X"38758f06",
X"ff055675",
X"83e7ec08",
X"2e9b3875",
X"83269638",
X"7583e7ec",
X"0c758429",
X"83ea9005",
X"70085355",
X"7551fa96",
X"3f807624",
X"88c93875",
X"842983ea",
X"90055574",
X"08802e88",
X"ba3883e7",
X"ec088429",
X"83ea9005",
X"70080288",
X"0582b905",
X"33525b55",
X"7480d22e",
X"84b13874",
X"80d22490",
X"3874bf2e",
X"9c387480",
X"d02e81d7",
X"3887f839",
X"7480d32e",
X"80d23874",
X"80d72e81",
X"c63887e7",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055656",
X"ffacfb3f",
X"80c151ff",
X"acb33ff6",
X"e73f860b",
X"83e7f034",
X"815283e7",
X"f051ffad",
X"d63f8151",
X"fde43f74",
X"8938860b",
X"83ea8c0c",
X"8739a80b",
X"83ea8c0c",
X"ffacc73f",
X"80c151ff",
X"abff3ff6",
X"b33f900b",
X"83ea8733",
X"81065656",
X"74802e83",
X"38985683",
X"e9fc3383",
X"e9fd3371",
X"882b0756",
X"59748180",
X"2e098106",
X"9c3883e9",
X"fa3383e9",
X"fb337188",
X"2b075657",
X"ad807527",
X"8c387581",
X"80075685",
X"3975a007",
X"567583e7",
X"f034ff0b",
X"83e7f134",
X"e00b83e7",
X"f234800b",
X"83e7f334",
X"845283e7",
X"f051ffac",
X"ca3f8451",
X"869e3902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"5659ffab",
X"b93f7951",
X"ffb6a63f",
X"83e08008",
X"802e8b38",
X"80ce51ff",
X"aae33f85",
X"f23980c1",
X"51ffaad9",
X"3fffabce",
X"3fffaa81",
X"3f83eaa0",
X"08588375",
X"259b3883",
X"e9fc3383",
X"e9fd3371",
X"882b07fc",
X"1771297a",
X"05838005",
X"5a51578d",
X"39748180",
X"2918ff80",
X"05588180",
X"57805676",
X"762e9338",
X"ffaab23f",
X"83e08008",
X"83e7f017",
X"34811656",
X"ea39ffaa",
X"a03f83e0",
X"800881ff",
X"06775383",
X"e7f05256",
X"f4d63f83",
X"e0800881",
X"ff065575",
X"752e0981",
X"06818a38",
X"ffaa9f3f",
X"80c151ff",
X"a9d73fff",
X"aacc3f77",
X"527951ff",
X"b4b53f80",
X"5e80d13d",
X"fdf40554",
X"765383e7",
X"f0527951",
X"ffb2c23f",
X"0282b905",
X"33558158",
X"7480d72e",
X"098106bd",
X"3880d13d",
X"fdf00554",
X"76538f3d",
X"70537a52",
X"59ffb3c7",
X"3f805676",
X"762ea238",
X"751983e7",
X"f0173371",
X"33707232",
X"70307080",
X"2570307e",
X"06811d5d",
X"5e515151",
X"525b55db",
X"3982ac51",
X"e4e63f77",
X"802e8638",
X"80c35184",
X"3980ce51",
X"ffa8d23f",
X"ffa9c73f",
X"ffa7fa3f",
X"83dd3902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"59558070",
X"5d59ffa8",
X"ed3f80c1",
X"51ffa8a5",
X"3f83ea88",
X"08792e82",
X"de3883ea",
X"a80880fc",
X"055580fd",
X"52745187",
X"ae3f83e0",
X"80085b77",
X"8224b238",
X"ff187087",
X"2b83ffff",
X"800680f7",
X"9c0583e7",
X"f0595755",
X"81805575",
X"70810557",
X"33777081",
X"055934ff",
X"157081ff",
X"06515574",
X"ea38828d",
X"397782e8",
X"2e81ab38",
X"7782e92e",
X"09810681",
X"b23880f5",
X"d451ffae",
X"a83f7858",
X"77873270",
X"30707207",
X"80257a8a",
X"32703070",
X"72078025",
X"73075354",
X"5a515755",
X"75802e97",
X"38787826",
X"9238a00b",
X"83e7f01a",
X"34811970",
X"81ff065a",
X"55eb3981",
X"187081ff",
X"0659558a",
X"7827ffbc",
X"388f5883",
X"e7eb1833",
X"83e7f019",
X"34ff1870",
X"81ff0659",
X"55778426",
X"ea389058",
X"800b83e7",
X"f0193481",
X"187081ff",
X"0670982b",
X"52595574",
X"8025e938",
X"80c6557a",
X"858f2484",
X"3880c255",
X"7483e7f0",
X"3480f10b",
X"83e7f334",
X"810b83e7",
X"f4347a83",
X"e7f1347a",
X"882c5574",
X"83e7f234",
X"80cb3982",
X"f0782580",
X"c4387780",
X"fd29fd97",
X"d3055279",
X"51ffb0e3",
X"3f80d13d",
X"fdec0554",
X"80fd5383",
X"e7f05279",
X"51ffb09b",
X"3f7b8119",
X"59567580",
X"fc248338",
X"78587788",
X"2c557483",
X"e8ed3477",
X"83e8ee34",
X"7583e8ef",
X"34818059",
X"80cc3983",
X"eaa00857",
X"8378259b",
X"3883e9fc",
X"3383e9fd",
X"3371882b",
X"07fc1a71",
X"29790583",
X"80055951",
X"598d3977",
X"81802917",
X"ff800557",
X"81805976",
X"527951ff",
X"aff13f80",
X"d13dfdec",
X"05547853",
X"83e7f052",
X"7951ffaf",
X"aa3f7851",
X"f6b83fff",
X"a5e43fff",
X"a4973f8b",
X"3983e9f0",
X"08810583",
X"e9f00c80",
X"d13d0d04",
X"f6d93fea",
X"f73ff939",
X"fc3d0d76",
X"78718429",
X"83ea9005",
X"70085153",
X"5353709e",
X"3880ce72",
X"3480cf0b",
X"81133480",
X"ce0b8213",
X"3480c50b",
X"83133470",
X"84133480",
X"e73983ea",
X"a4133354",
X"80d27234",
X"73822a70",
X"81065151",
X"80cf5370",
X"843880d7",
X"53728113",
X"34a00b82",
X"13347383",
X"06517081",
X"2e9e3870",
X"81248838",
X"70802e8f",
X"389f3970",
X"822e9238",
X"70832e92",
X"38933980",
X"d8558e39",
X"80d35589",
X"3980cd55",
X"843980c4",
X"55748313",
X"3480c40b",
X"84133480",
X"0b851334",
X"863d0d04",
X"fd3d0d75",
X"5480740c",
X"800b8415",
X"0c800b88",
X"150c800b",
X"8c150c87",
X"a6803370",
X"81ff0651",
X"51defc3f",
X"70812a81",
X"32718132",
X"71810671",
X"81063184",
X"170c5353",
X"70832a81",
X"3271822a",
X"81327181",
X"06718106",
X"31760c52",
X"5287a090",
X"33700981",
X"0688160c",
X"5183e080",
X"08802e80",
X"c23883e0",
X"8008812a",
X"70810683",
X"e0800881",
X"06318416",
X"0c5183e0",
X"8008832a",
X"83e08008",
X"822a7181",
X"06718106",
X"31760c52",
X"5283e080",
X"08842a81",
X"0688150c",
X"83e08008",
X"852a8106",
X"8c150c85",
X"3d0d04fe",
X"3d0d7476",
X"54527151",
X"fece3f72",
X"812ea238",
X"8173268d",
X"3872822e",
X"a8387283",
X"2e9c38e6",
X"397108e2",
X"38841208",
X"dd388812",
X"08d838a5",
X"39881208",
X"812e9e38",
X"91398812",
X"08812e95",
X"38710891",
X"38841208",
X"8c388c12",
X"08812e09",
X"8106ffb2",
X"38843d0d",
X"04fc3d0d",
X"76785354",
X"81538055",
X"87397110",
X"73105452",
X"73722651",
X"72802ea7",
X"3870802e",
X"86387180",
X"25e83872",
X"802e9838",
X"71742689",
X"38737231",
X"75740756",
X"5472812a",
X"72812a53",
X"53e53973",
X"51788338",
X"74517083",
X"e0800c86",
X"3d0d04fe",
X"3d0d8053",
X"75527451",
X"ffa33f84",
X"3d0d04fe",
X"3d0d8153",
X"75527451",
X"ff933f84",
X"3d0d04fb",
X"3d0d7779",
X"55558056",
X"74762586",
X"38743055",
X"81567380",
X"25883873",
X"30768132",
X"57548053",
X"73527451",
X"fee73f83",
X"e0800854",
X"75802e87",
X"3883e080",
X"08305473",
X"83e0800c",
X"873d0d04",
X"fa3d0d78",
X"7a575580",
X"57747725",
X"86387430",
X"55815775",
X"9f2c5481",
X"53757432",
X"74315274",
X"51feaa3f",
X"83e08008",
X"5476802e",
X"873883e0",
X"80083054",
X"7383e080",
X"0c883d0d",
X"04000000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002aa7",
X"00002ae8",
X"00002b0a",
X"00002b31",
X"00002b31",
X"00002b31",
X"00002b31",
X"00002ba2",
X"00002bf4",
X"25732025",
X"73000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"6e616d65",
X"20000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00003a14",
X"00003a18",
X"00003a20",
X"00003a2c",
X"00003a38",
X"00003a44",
X"00003a50",
X"00003a54",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
