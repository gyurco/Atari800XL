
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81d9",
X"cc738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81e1",
X"fc0c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757580f4",
X"c12d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7580f480",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80de8f04",
X"fd3d0d75",
X"705254ae",
X"a33f83c0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"c0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83c0",
X"8008732e",
X"a13883c0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183c0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83c2d008",
X"248a38b4",
X"f43fff0b",
X"83c2d00c",
X"800b83c0",
X"800c04ff",
X"3d0d7352",
X"83c0ac08",
X"722e8d38",
X"d93f7151",
X"96993f71",
X"83c0ac0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"558154bc",
X"15088191",
X"387451cf",
X"3f795880",
X"7a2580f7",
X"3883c380",
X"0870892a",
X"5783ff06",
X"78848072",
X"31565657",
X"73782583",
X"38735575",
X"83c2d008",
X"2e8438ff",
X"893f83c2",
X"d0088025",
X"a6387589",
X"2b5198dc",
X"3f83c380",
X"088f3dfc",
X"11555c54",
X"8152f81b",
X"5196c63f",
X"761483c3",
X"800c7583",
X"c2d00c74",
X"53765278",
X"51b3a53f",
X"83c08008",
X"83c38008",
X"1683c380",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8b3861",
X"7a710c54",
X"75547580",
X"2e833881",
X"547383c0",
X"800c8e3d",
X"0d04fc3d",
X"0dfe9b3f",
X"7651feaf",
X"3f863dfc",
X"05537852",
X"775195e9",
X"3f797571",
X"0c5483c0",
X"80085483",
X"c0800880",
X"2e833881",
X"547383c0",
X"800c863d",
X"0d04fe3d",
X"0d7583c2",
X"d0085353",
X"80722489",
X"3871732e",
X"8438fdd6",
X"3f7451fd",
X"ea3f7251",
X"97ae3f83",
X"c0800852",
X"83c08008",
X"802e8338",
X"81527183",
X"c0800c84",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"c0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"c0800c51",
X"823d0d04",
X"80c40b83",
X"c0800c04",
X"fd3d0d75",
X"77715470",
X"535553a9",
X"fb3f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfceb3f",
X"735193ab",
X"3f7383c0",
X"ac0c83c0",
X"80085383",
X"c0800880",
X"2e833881",
X"537283c0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcbf3f",
X"72802ea5",
X"38bc1308",
X"527351a9",
X"853f83c0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"c0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83c0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83c2d0",
X"0c7483c0",
X"b00c7583",
X"c2cc0caf",
X"d93f83c0",
X"800881ff",
X"06528153",
X"71993883",
X"c2e8518e",
X"943f83c0",
X"80085283",
X"c0800880",
X"2e833872",
X"52715372",
X"83c0800c",
X"843d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"51a6f63f",
X"83c08008",
X"557483c0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"c0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283c2cc",
X"085180e3",
X"833f83c0",
X"800857f9",
X"e13f7952",
X"83c2d451",
X"95b73f83",
X"c0800854",
X"805383c0",
X"8008732e",
X"09810682",
X"833883c0",
X"b0080b0b",
X"81deec53",
X"705256a6",
X"b33f0b0b",
X"81deec52",
X"80c01651",
X"a6a63f75",
X"bc170c73",
X"82c0170c",
X"810b82c4",
X"170c810b",
X"82c8170c",
X"7382cc17",
X"0cff1782",
X"d0175557",
X"81913983",
X"c0bc3370",
X"822a7081",
X"06515455",
X"72818038",
X"74812a81",
X"06587780",
X"f6387484",
X"2a810682",
X"c4150c83",
X"c0bc3381",
X"0682c815",
X"0c795273",
X"51a5cd3f",
X"7351a5e4",
X"3f83c080",
X"081453af",
X"73708105",
X"553472bc",
X"150c83c0",
X"bd527251",
X"a5ae3f83",
X"c0b40882",
X"c0150c83",
X"c0ca5280",
X"c01451a5",
X"9b3f7880",
X"2e8d3873",
X"51782d83",
X"c0800880",
X"2e993877",
X"82cc150c",
X"75802e86",
X"387382cc",
X"170c7382",
X"d015ff19",
X"59555676",
X"802e9b38",
X"83c0b452",
X"83c2d451",
X"94ad3f83",
X"c080088a",
X"3883c0bd",
X"335372fe",
X"d2387880",
X"2e893883",
X"c0b00851",
X"fcb83f83",
X"c0b00853",
X"7283c080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb53f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f690",
X"3f83c080",
X"08745387",
X"3d705355",
X"55f6b03f",
X"f7903f73",
X"51d33f63",
X"53745283",
X"c0800851",
X"fab83f92",
X"3d0d0471",
X"83c0800c",
X"0480c012",
X"83c0800c",
X"04803d0d",
X"7282c011",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"c0800c51",
X"823d0d04",
X"f93d0d79",
X"83c09008",
X"57578177",
X"27819638",
X"76881708",
X"27818e38",
X"75335574",
X"822e8938",
X"74832eb3",
X"3880fe39",
X"74547610",
X"83fe0653",
X"76882a8c",
X"17080552",
X"893dfc05",
X"51aa873f",
X"83c08008",
X"80df3802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d13984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"51a9d73f",
X"83c08008",
X"b038029f",
X"05330284",
X"059e0533",
X"71982b71",
X"902b0702",
X"8c059d05",
X"3370882b",
X"72078d3d",
X"337180ff",
X"fffe8006",
X"07515253",
X"57585683",
X"39815574",
X"83c0800c",
X"893d0d04",
X"fb3d0d83",
X"c09008fe",
X"19881208",
X"fe055556",
X"54805674",
X"73278d38",
X"82143375",
X"71299416",
X"08055753",
X"7583c080",
X"0c873d0d",
X"04fc3d0d",
X"7652800b",
X"83c09008",
X"70335152",
X"5370832e",
X"09810691",
X"38951233",
X"94133371",
X"982b7190",
X"2b075555",
X"519b1233",
X"9a133371",
X"882b0774",
X"0783c080",
X"0c55863d",
X"0d04fc3d",
X"0d7683c0",
X"90085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"fed63f83",
X"c0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183c080",
X"0c863d0d",
X"04fa3d0d",
X"7883c090",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fcb13f",
X"81527183",
X"c0800827",
X"a8388352",
X"83c08008",
X"88170827",
X"9c3883c0",
X"80088c16",
X"0c83c080",
X"0851fdbc",
X"3f83c080",
X"0890160c",
X"73752380",
X"527183c0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585e5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"9f269138",
X"7a51fdd2",
X"3f83c080",
X"0856807d",
X"34838139",
X"933d841c",
X"08705859",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"3880705a",
X"5c887f08",
X"5f5a7b81",
X"1d7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535e57",
X"557480e7",
X"3876ae2e",
X"09810683",
X"38815578",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675bb",
X"3888598b",
X"5affab39",
X"76982b55",
X"74802587",
X"3881d8dc",
X"173357ff",
X"9f175574",
X"99268938",
X"e0177081",
X"ff065855",
X"78811a70",
X"81ff0672",
X"1b535b57",
X"55767534",
X"fef8397b",
X"1e7f0c80",
X"5576a026",
X"83388155",
X"748b1934",
X"7a51fc82",
X"3f83c080",
X"0880f538",
X"a0547a22",
X"70852b83",
X"e0065455",
X"901b0852",
X"7c51a492",
X"3f83c080",
X"085783c0",
X"80088181",
X"387c3355",
X"74802e80",
X"f4388b1d",
X"3370832a",
X"70810651",
X"565674b4",
X"388b7d84",
X"1d0883c0",
X"8008595b",
X"5b58ff18",
X"5877ff2e",
X"9a387970",
X"81055b33",
X"79708105",
X"5b337171",
X"31525656",
X"75802ee2",
X"38863975",
X"802e9638",
X"7a51fbe5",
X"3fff8639",
X"83c08008",
X"5683c080",
X"08b63883",
X"39765684",
X"1b088b11",
X"33515574",
X"a7388b1d",
X"3370842a",
X"70810651",
X"56567489",
X"38835694",
X"39815690",
X"397c51fa",
X"943f83c0",
X"8008881c",
X"0cfd8139",
X"7583c080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"51a2d73f",
X"835683c0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"51a2ab3f",
X"83c08008",
X"98388117",
X"33773371",
X"882b0783",
X"c0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"7651a282",
X"3f83c080",
X"08983881",
X"17337733",
X"71882b07",
X"83c08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583c080",
X"0c8a3d0d",
X"04eb3d0d",
X"675a800b",
X"83c0900c",
X"a1a43f83",
X"c0800881",
X"06558256",
X"7483ef38",
X"7475538f",
X"3d705357",
X"59feca3f",
X"83c08008",
X"81ff0657",
X"76812e09",
X"810680d4",
X"38905483",
X"be537452",
X"7551a196",
X"3f83c080",
X"0880c938",
X"8f3d3355",
X"74802e80",
X"c93802bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"33710770",
X"587b575e",
X"525e5759",
X"57fdee3f",
X"83c08008",
X"81ff0657",
X"76832e09",
X"81068638",
X"815682f2",
X"3976802e",
X"86388656",
X"82e839a4",
X"548d5378",
X"527551a0",
X"ad3f8156",
X"83c08008",
X"82d43802",
X"be053302",
X"8405bd05",
X"3371882b",
X"07595d77",
X"ab380280",
X"ce053302",
X"840580cd",
X"05337198",
X"2b71902b",
X"07973d33",
X"70882b72",
X"07029405",
X"80cb0533",
X"71075452",
X"5e575956",
X"02b70533",
X"78712902",
X"8805b605",
X"33028c05",
X"b5053371",
X"882b0770",
X"1d707f8c",
X"050c5f59",
X"57595d8e",
X"3d33821b",
X"3402b905",
X"33903d33",
X"71882b07",
X"5a5c7884",
X"1b2302bb",
X"05330284",
X"05ba0533",
X"71882b07",
X"565c74ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"07515253",
X"575e5c74",
X"76317831",
X"79842a90",
X"3d335471",
X"71315356",
X"5680d3e8",
X"3f83c080",
X"08820570",
X"881c0c83",
X"c08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83c0900c",
X"80567583",
X"c0800c97",
X"3d0d04e9",
X"3d0d83c0",
X"90085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e53f83c0",
X"80085483",
X"c0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f489",
X"3f83c080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383c080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83c09008",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0e93f",
X"83c08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"833f83c0",
X"80085583",
X"c0800880",
X"2eff8938",
X"83c08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"519ad33f",
X"83c08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83c0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83c09008",
X"55568555",
X"73802e81",
X"e3388114",
X"33810653",
X"84557280",
X"2e81d538",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b9388214",
X"3370892b",
X"56537680",
X"2eb73874",
X"52ff1651",
X"80cee93f",
X"83c08008",
X"ff187654",
X"70535853",
X"80ced93f",
X"83c08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed63f83",
X"c0800853",
X"810b83c0",
X"8008278b",
X"38881408",
X"83c08008",
X"26883880",
X"0b811534",
X"b03983c0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc53f",
X"83c08008",
X"8c3883c0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683c0",
X"800805a8",
X"150c8055",
X"7483c080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83c09008",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1cf3f",
X"83c08008",
X"5583c080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef5",
X"3f83c080",
X"0888170c",
X"7551efa6",
X"3f83c080",
X"08557483",
X"c0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683c0",
X"9008802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f53f83c0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"96dc3f83",
X"c0800841",
X"83c08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"eddf3f83",
X"c0800841",
X"83c08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"8e823f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f03f83c0",
X"80088332",
X"70307072",
X"079f2c83",
X"c0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"8c8e3f75",
X"83c0800c",
X"9e3d0d04",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"7751e0d2",
X"3f83c080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3381e284",
X"0b81e284",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"527751e0",
X"813f83c0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583c0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"558b953f",
X"83c08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"8114518a",
X"ad3f83c0",
X"80083070",
X"83c08008",
X"07802583",
X"c0800c53",
X"863d0d04",
X"fc3d0d76",
X"705255e6",
X"ee3f83c0",
X"80085481",
X"5383c080",
X"0880c138",
X"7451e6b1",
X"3f83c080",
X"0881defc",
X"5383c080",
X"085253ff",
X"913f83c0",
X"8008a138",
X"81df8052",
X"7251ff82",
X"3f83c080",
X"08923881",
X"df845272",
X"51fef33f",
X"83c08008",
X"802e8338",
X"81547353",
X"7283c080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"e68d3f81",
X"5383c080",
X"08983873",
X"51e5d63f",
X"83c39808",
X"5283c080",
X"0851feba",
X"3f83c080",
X"08537283",
X"c0800c85",
X"3d0d04df",
X"3d0da43d",
X"0870525e",
X"dbfb3f83",
X"c0800833",
X"953d5654",
X"73963881",
X"e5d45274",
X"51898d3f",
X"9a397d52",
X"7851defc",
X"3f84d039",
X"7d51dbe1",
X"3f83c080",
X"08527451",
X"db913f80",
X"43804280",
X"41804083",
X"c3a00852",
X"943d7052",
X"5de1e43f",
X"83c08008",
X"59800b83",
X"c0800855",
X"5b83c080",
X"087b2e94",
X"38811b74",
X"525be4e6",
X"3f83c080",
X"085483c0",
X"8008ee38",
X"805aff5f",
X"7909709f",
X"2c7b065b",
X"547a7a24",
X"8438ff1b",
X"5af61a70",
X"09709f2c",
X"72067bff",
X"125a5a52",
X"55558075",
X"25953876",
X"51e4ab3f",
X"83c08008",
X"76ff1858",
X"55577380",
X"24ed3874",
X"7f2e8638",
X"a1b53f74",
X"5f78ff1b",
X"70585d58",
X"807a2595",
X"387751e4",
X"813f83c0",
X"800876ff",
X"18585558",
X"738024ed",
X"38800b83",
X"c7d00c80",
X"0b83c884",
X"0c81df88",
X"518d8c3f",
X"81800b83",
X"c8840c81",
X"df90518c",
X"fe3fa80b",
X"83c7d00c",
X"76802e80",
X"e43883c7",
X"d0087779",
X"32703070",
X"72078025",
X"70872b83",
X"c8840c51",
X"56785356",
X"56e3b83f",
X"83c08008",
X"802e8838",
X"81df9851",
X"8cc53f76",
X"51e2fa3f",
X"83c08008",
X"5281e0b8",
X"518cb43f",
X"7651e382",
X"3f83c080",
X"0883c7d0",
X"08555775",
X"74258638",
X"a81656f7",
X"397583c7",
X"d00c86f0",
X"7624ff98",
X"3887980b",
X"83c7d00c",
X"77802eb1",
X"387751e2",
X"b83f83c0",
X"80087852",
X"55e2d83f",
X"81dfa054",
X"83c08008",
X"8d388739",
X"80763481",
X"d03981df",
X"9c547453",
X"735281de",
X"f0518bd3",
X"3f805481",
X"def8518b",
X"ca3f8114",
X"5473a82e",
X"098106ef",
X"38868da0",
X"519da83f",
X"8052903d",
X"70525780",
X"c4d63f83",
X"52765180",
X"c4ce3f62",
X"818f3861",
X"802e80fb",
X"387b5473",
X"ff2e9638",
X"78802e81",
X"8a387851",
X"e1dc3f83",
X"c08008ff",
X"155559e7",
X"3978802e",
X"80f53878",
X"51e1d83f",
X"83c08008",
X"802efc8e",
X"387851e1",
X"a03f83c0",
X"80085281",
X"deec5183",
X"e03f83c0",
X"8008a338",
X"7c518598",
X"3f83c080",
X"085574ff",
X"16565480",
X"7425ae38",
X"741d7033",
X"555673af",
X"2efecd38",
X"e9397851",
X"e0e13f83",
X"c0800852",
X"7c5184d0",
X"3f8f397f",
X"88296010",
X"057a0561",
X"055afc90",
X"3962802e",
X"fbd13880",
X"52765180",
X"c3ae3fa3",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067084",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d38a8",
X"0b9088b8",
X"34b80b90",
X"88b83470",
X"83c0800c",
X"823d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"852a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"980b9088",
X"b834b80b",
X"9088b834",
X"7083c080",
X"0c823d0d",
X"04930b90",
X"88bc34ff",
X"0b9088a8",
X"3404ff3d",
X"0d028f05",
X"3352800b",
X"9088bc34",
X"8a519aef",
X"3fdf3f80",
X"f80b9088",
X"a034800b",
X"90888834",
X"fa125271",
X"90888034",
X"800b9088",
X"98347190",
X"88903490",
X"88b85280",
X"7234b872",
X"34833d0d",
X"04803d0d",
X"028b0533",
X"51709088",
X"b434febf",
X"3f83c080",
X"08802ef6",
X"38823d0d",
X"04803d0d",
X"8439a6af",
X"3ffed93f",
X"83c08008",
X"802ef338",
X"9088b433",
X"7081ff06",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"a30b9088",
X"bc34ff0b",
X"9088a834",
X"9088b851",
X"a87134b8",
X"7134823d",
X"0d04803d",
X"0d9088bc",
X"3370982b",
X"70802583",
X"c0800c51",
X"51823d0d",
X"04803d0d",
X"9088b833",
X"7081ff06",
X"70832a81",
X"32708106",
X"51515151",
X"70802ee8",
X"38b00b90",
X"88b834b8",
X"0b9088b8",
X"34823d0d",
X"04803d0d",
X"9080ac08",
X"810683c0",
X"800c823d",
X"0d04fd3d",
X"0d757754",
X"54807325",
X"94387370",
X"81055533",
X"5281dfa4",
X"5187843f",
X"ff1353e9",
X"39853d0d",
X"04fd3d0d",
X"75775354",
X"73335170",
X"89387133",
X"5170802e",
X"a1387333",
X"72335253",
X"72712785",
X"38ff5194",
X"39707327",
X"85388151",
X"8b398114",
X"81135354",
X"d3398051",
X"7083c080",
X"0c853d0d",
X"04fd3d0d",
X"75775454",
X"72337081",
X"ff065252",
X"70802ea3",
X"387181ff",
X"068114ff",
X"bf125354",
X"52709926",
X"8938a012",
X"7081ff06",
X"53517174",
X"70810556",
X"34d23980",
X"7434853d",
X"0d04ffbd",
X"3d0d80c6",
X"3d0852a5",
X"3d705254",
X"ffb33f80",
X"c73d0852",
X"853d7052",
X"53ffa63f",
X"72527351",
X"fedf3f80",
X"c53d0d04",
X"fe3d0d74",
X"76535371",
X"70810553",
X"33517073",
X"70810555",
X"3470f038",
X"843d0d04",
X"fe3d0d74",
X"52807233",
X"52537073",
X"2e8d3881",
X"12811471",
X"33535452",
X"70f53872",
X"83c0800c",
X"843d0d04",
X"f63d0d7c",
X"7e60625a",
X"5d5b5680",
X"59815585",
X"39747a29",
X"55745275",
X"51bbc13f",
X"83c08008",
X"7a27ee38",
X"74802e80",
X"dd387452",
X"7551bbac",
X"3f83c080",
X"08755376",
X"5254bbb0",
X"3f83c080",
X"087a5375",
X"5256bb94",
X"3f83c080",
X"08793070",
X"7b079f2a",
X"70778024",
X"07515154",
X"55728738",
X"83c08008",
X"c5387681",
X"18b01655",
X"58588974",
X"258b38b7",
X"14537a85",
X"3880d714",
X"53727834",
X"811959ff",
X"9f398077",
X"348c3d0d",
X"04f73d0d",
X"7b7d7f62",
X"029005bb",
X"05335759",
X"565a5ab0",
X"58728338",
X"a0587570",
X"70810552",
X"33715954",
X"55903980",
X"74258e38",
X"ff147770",
X"81055933",
X"545472ef",
X"3873ff15",
X"55538073",
X"25893877",
X"52795178",
X"2def3975",
X"33755753",
X"72802e90",
X"38725279",
X"51782d75",
X"70810557",
X"3353ed39",
X"8b3d0d04",
X"ee3d0d64",
X"66696970",
X"70810552",
X"335b4a5c",
X"5e5e7680",
X"2e82f938",
X"76a52e09",
X"810682e0",
X"38807041",
X"67707081",
X"05523371",
X"4a59575f",
X"76b02e09",
X"81068c38",
X"75708105",
X"57337648",
X"57815fd0",
X"17567589",
X"2680da38",
X"76675c59",
X"805c9339",
X"778a2480",
X"c3387b8a",
X"29187b70",
X"81055d33",
X"5a5cd019",
X"7081ff06",
X"58588977",
X"27a438ff",
X"9f197081",
X"ff06ffa9",
X"1b5a5156",
X"85762792",
X"38ffbf19",
X"7081ff06",
X"51567585",
X"268a38c9",
X"19587780",
X"25ffb938",
X"7a477b40",
X"7881ff06",
X"577680e4",
X"2e80e538",
X"7680e424",
X"a7387680",
X"d82e8186",
X"387680d8",
X"24903876",
X"802e81cc",
X"3876a52e",
X"81b63881",
X"b9397680",
X"e32e818c",
X"3881af39",
X"7680f52e",
X"9b387680",
X"f5248b38",
X"7680f32e",
X"81813881",
X"99397680",
X"f82e80ca",
X"38818f39",
X"913d7055",
X"5780538a",
X"5279841b",
X"7108535b",
X"56fc813f",
X"7655ab39",
X"79841b71",
X"08943d70",
X"5b5b525b",
X"56758025",
X"8c387530",
X"56ad7834",
X"0280c105",
X"57765480",
X"538a5275",
X"51fbd53f",
X"77557e54",
X"b839913d",
X"70557780",
X"d8327030",
X"70802556",
X"51585690",
X"5279841b",
X"7108535b",
X"57fbb13f",
X"7555db39",
X"79841b83",
X"1233545b",
X"56983979",
X"841b7108",
X"575b5680",
X"547f537c",
X"527d51fc",
X"9c3f8739",
X"76527d51",
X"7c2d6670",
X"33588105",
X"47fd8339",
X"943d0d04",
X"7283c094",
X"0c7183c0",
X"980c04fb",
X"3d0d883d",
X"70708405",
X"52085754",
X"755383c0",
X"94085283",
X"c0980851",
X"fcc63f87",
X"3d0d04ff",
X"3d0d7370",
X"08535102",
X"93053372",
X"34700881",
X"05710c83",
X"3d0d04fc",
X"3d0d873d",
X"88115578",
X"54bdb753",
X"51fc993f",
X"8052873d",
X"51d13f86",
X"3d0d04fc",
X"3d0d7655",
X"7483c3ac",
X"082eaf38",
X"80537451",
X"87c13f83",
X"c0800881",
X"ff06ff14",
X"7081ff06",
X"7230709f",
X"2a515255",
X"53547280",
X"2e843871",
X"dd3873fe",
X"387483c3",
X"ac0c863d",
X"0d04ff3d",
X"0dff0b83",
X"c3ac0c84",
X"a53f8151",
X"87853f83",
X"c0800881",
X"ff065271",
X"ee3881d3",
X"3f7183c0",
X"800c833d",
X"0d04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"823f7280",
X"2ea03883",
X"c3c01433",
X"75708105",
X"57348114",
X"7083ffff",
X"06ff1570",
X"83ffff06",
X"56525552",
X"dd39800b",
X"83c0800c",
X"863d0d04",
X"fc3d0d76",
X"787a1156",
X"53558053",
X"71742e93",
X"38721551",
X"703383c3",
X"c0133481",
X"12811454",
X"52ea3980",
X"0b83c080",
X"0c863d0d",
X"04fd3d0d",
X"905483c3",
X"ac085186",
X"f43f83c0",
X"800881ff",
X"06ff1571",
X"30713070",
X"73079f2a",
X"729f2a06",
X"52555255",
X"5372db38",
X"853d0d04",
X"803d0d83",
X"c3b80810",
X"83c3b008",
X"079080a8",
X"0c823d0d",
X"04800b83",
X"c3b80ce4",
X"3f04810b",
X"83c3b80c",
X"db3f04ed",
X"3f047183",
X"c3b40c04",
X"803d0d80",
X"51f43f81",
X"0b83c3b8",
X"0c810b83",
X"c3b00cff",
X"bb3f823d",
X"0d04803d",
X"0d723070",
X"74078025",
X"83c3b00c",
X"51ffa53f",
X"823d0d04",
X"803d0d02",
X"8b053390",
X"80a40c90",
X"80a80870",
X"81065151",
X"70f53890",
X"80a40870",
X"81ff0683",
X"c0800c51",
X"823d0d04",
X"803d0d81",
X"ff51d13f",
X"83c08008",
X"81ff0683",
X"c0800c82",
X"3d0d0480",
X"3d0d7390",
X"2b730790",
X"80b40c82",
X"3d0d0404",
X"fb3d0d78",
X"0284059f",
X"05337098",
X"2b555755",
X"7280259b",
X"387580ff",
X"06568052",
X"80f751e0",
X"3f83c080",
X"0881ff06",
X"54738126",
X"80ff3880",
X"51fee73f",
X"ffa23f81",
X"51fedf3f",
X"ff9a3f75",
X"51feed3f",
X"74982a51",
X"fee63f74",
X"902a7081",
X"ff065253",
X"feda3f74",
X"882a7081",
X"ff065253",
X"fece3f74",
X"81ff0651",
X"fec63f81",
X"557580c0",
X"2e098106",
X"86388195",
X"558d3975",
X"80c82e09",
X"81068438",
X"81875574",
X"51fea53f",
X"8a55fec8",
X"3f83c080",
X"0881ff06",
X"70982b54",
X"54728025",
X"8c38ff15",
X"7081ff06",
X"565374e2",
X"387383c0",
X"800c873d",
X"0d04fa3d",
X"0dfdc53f",
X"8051fdda",
X"3f8a54fe",
X"933fff14",
X"7081ff06",
X"555373f3",
X"38737453",
X"5580c051",
X"fea63f83",
X"c0800881",
X"ff065473",
X"812e0981",
X"06829f38",
X"83aa5280",
X"c851fe8c",
X"3f83c080",
X"0881ff06",
X"5372812e",
X"09810681",
X"a8387454",
X"873d7411",
X"5456fdc8",
X"3f83c080",
X"08733481",
X"147081ff",
X"06555383",
X"7427e538",
X"029a0533",
X"5372812e",
X"09810681",
X"d938029b",
X"05335380",
X"ce905472",
X"81aa2e8d",
X"3881c739",
X"80e4518b",
X"9a3fff14",
X"5473802e",
X"81b83882",
X"0a5281e9",
X"51fda53f",
X"83c08008",
X"81ff0653",
X"72de3872",
X"5280fa51",
X"fd923f83",
X"c0800881",
X"ff065372",
X"81903872",
X"54731653",
X"fcd63f83",
X"c0800873",
X"34811470",
X"81ff0655",
X"53837427",
X"e838873d",
X"3370862a",
X"70810651",
X"54548c55",
X"7280e338",
X"845580de",
X"39745281",
X"e951fccc",
X"3f83c080",
X"0881ff06",
X"53825581",
X"e9568173",
X"27863873",
X"5580c156",
X"80ce9054",
X"8a3980e4",
X"518a8c3f",
X"ff145473",
X"802ea938",
X"80527551",
X"fc9a3f83",
X"c0800881",
X"ff065372",
X"e1388480",
X"5280d051",
X"fc863f83",
X"c0800881",
X"ff065372",
X"802e8338",
X"80557483",
X"c3bc3480",
X"51fb873f",
X"fbc23f88",
X"3d0d04fb",
X"3d0d7754",
X"800b83c3",
X"bc337083",
X"2a708106",
X"51555755",
X"72752e09",
X"81068538",
X"73892b54",
X"735280d1",
X"51fbbd3f",
X"83c08008",
X"81ff0653",
X"72bd3882",
X"b8c054fb",
X"833f83c0",
X"800881ff",
X"06537281",
X"ff2e0981",
X"068938ff",
X"145473e7",
X"389f3972",
X"81fe2e09",
X"81069638",
X"83c7c052",
X"83c3c051",
X"faed3ffa",
X"d33ffad0",
X"3f833981",
X"558051fa",
X"893ffac4",
X"3f7481ff",
X"0683c080",
X"0c873d0d",
X"04fb3d0d",
X"7783c3c0",
X"56548151",
X"f9ec3f83",
X"c3bc3370",
X"832a7081",
X"06515456",
X"72853873",
X"892b5473",
X"5280d851",
X"fab63f83",
X"c0800881",
X"ff065372",
X"80e43881",
X"ff51f9d4",
X"3f81fe51",
X"f9ce3f84",
X"80537470",
X"81055633",
X"51f9c13f",
X"ff137083",
X"ffff0651",
X"5372eb38",
X"7251f9b0",
X"3f7251f9",
X"ab3ff9d0",
X"3f83c080",
X"089f0653",
X"a7885472",
X"852e8c38",
X"993980e4",
X"5187c43f",
X"ff1454f9",
X"b33f83c0",
X"800881ff",
X"2e843873",
X"e9388051",
X"f8e43ff9",
X"9f3f800b",
X"83c0800c",
X"873d0d04",
X"7183c7c4",
X"0c888080",
X"0b83c7c0",
X"0c848080",
X"0b83c7c8",
X"0c04fd3d",
X"0d777017",
X"557705ff",
X"1a535371",
X"ff2e9438",
X"73708105",
X"55335170",
X"73708105",
X"5534ff12",
X"52e93985",
X"3d0d04fb",
X"3d0d87a6",
X"810b83c7",
X"c4085656",
X"753383a6",
X"801634a0",
X"5483a080",
X"5383c7c4",
X"085283c7",
X"c00851ff",
X"b13fa054",
X"83a48053",
X"83c7c408",
X"5283c7c0",
X"0851ff9e",
X"3f905483",
X"a8805383",
X"c7c40852",
X"83c7c008",
X"51ff8b3f",
X"a0538052",
X"83c7c808",
X"83a08005",
X"5186953f",
X"a0538052",
X"83c7c808",
X"83a48005",
X"5186853f",
X"90538052",
X"83c7c808",
X"83a88005",
X"5185f53f",
X"ff763483",
X"a0805480",
X"5383c7c4",
X"085283c7",
X"c80851fe",
X"c53f80d0",
X"805483b0",
X"805383c7",
X"c4085283",
X"c7c80851",
X"feb03f87",
X"ba3fa254",
X"805383c7",
X"c8088c80",
X"055281e2",
X"f851fe9a",
X"3f860b87",
X"a8833480",
X"0b87a882",
X"34800b87",
X"a09a34af",
X"0b87a096",
X"34bf0b87",
X"a0973480",
X"0b87a098",
X"349f0b87",
X"a0993480",
X"0b87a09b",
X"34e00b87",
X"a88934a2",
X"0b87a880",
X"34830b87",
X"a48f3482",
X"0b87a881",
X"34873d0d",
X"04fc3d0d",
X"83a08054",
X"805383c7",
X"c8085283",
X"c7c40851",
X"fdb83f80",
X"d0805483",
X"b0805383",
X"c7c80852",
X"83c7c408",
X"51fda33f",
X"a05483a0",
X"805383c7",
X"c8085283",
X"c7c40851",
X"fd903fa0",
X"5483a480",
X"5383c7c8",
X"085283c7",
X"c40851fc",
X"fd3f9054",
X"83a88053",
X"83c7c808",
X"5283c7c4",
X"0851fcea",
X"3f83c7c4",
X"085583a6",
X"80153387",
X"a6813486",
X"3d0d04fa",
X"3d0d7870",
X"5255c1e3",
X"3f83ffff",
X"0b83c080",
X"0825a938",
X"7451c1e4",
X"3f83c080",
X"089e3883",
X"c0800857",
X"883dfc05",
X"54848080",
X"5383c7c4",
X"08527451",
X"ffbf9d3f",
X"ffbee33f",
X"883d0d04",
X"fa3d0d78",
X"705255c1",
X"a23f83ff",
X"ff0b83c0",
X"80082596",
X"38805788",
X"3dfc0554",
X"84808053",
X"83c7c408",
X"527451c0",
X"953f883d",
X"0d04803d",
X"0d908090",
X"08810683",
X"c0800c82",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe067607",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"812c8106",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fd06",
X"76100772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087082",
X"2cbf0683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fe8306",
X"76822b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"882c8706",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f1ff",
X"0676882b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70912cbf",
X"0683c080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870fc",
X"87ffff06",
X"76912b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"992c8106",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870ffbf",
X"0a067699",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908080",
X"0870882c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"80087089",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8a2c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708b2c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708c2c",
X"bf0683c0",
X"800c5182",
X"3d0d04fe",
X"3d0d7481",
X"e629872a",
X"9080a00c",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d848080",
X"53805288",
X"800a51ff",
X"b33f8180",
X"80538052",
X"82800a51",
X"c63f843d",
X"0d04803d",
X"0d8151fc",
X"aa3f7280",
X"2e903880",
X"51fdfe3f",
X"cd3f83c7",
X"cc3351fd",
X"f43f8151",
X"fcbb3f80",
X"51fcb63f",
X"8051fc87",
X"3f823d0d",
X"04fd3d0d",
X"75528054",
X"80ff7225",
X"8838810b",
X"ff801353",
X"54ffbf12",
X"51709926",
X"8638e012",
X"52b039ff",
X"9f125199",
X"7127a738",
X"d012e013",
X"54517089",
X"26853872",
X"52983972",
X"8f268538",
X"72528f39",
X"71ba2e09",
X"81068538",
X"9a528339",
X"80527380",
X"2e853881",
X"80125271",
X"81ff0683",
X"c0800c85",
X"3d0d0480",
X"3d0d84d8",
X"c0518071",
X"70810553",
X"347084e0",
X"c02e0981",
X"06f03882",
X"3d0d04fe",
X"3d0d0297",
X"053351fe",
X"f43f83c0",
X"800881ff",
X"0683c7d0",
X"08545280",
X"73249b38",
X"83c88008",
X"137283c8",
X"84080753",
X"53717334",
X"83c7d008",
X"810583c7",
X"d00c843d",
X"0d04fa3d",
X"0d82800a",
X"1b558057",
X"883dfc05",
X"54795374",
X"527851ff",
X"baac3f88",
X"3d0d04fe",
X"3d0d83c7",
X"e8085274",
X"51c1903f",
X"83c08008",
X"8c387653",
X"755283c7",
X"e80851c6",
X"3f843d0d",
X"04fe3d0d",
X"83c7e808",
X"53755274",
X"51ffbbce",
X"3f83c080",
X"088d3877",
X"53765283",
X"c7e80851",
X"ffa03f84",
X"3d0d04fe",
X"3d0d83c7",
X"e80851ff",
X"bac13f83",
X"c0800881",
X"80802e09",
X"81068838",
X"83c18080",
X"539c3983",
X"c7e80851",
X"ffbaa43f",
X"83c08008",
X"80d0802e",
X"09810693",
X"3883c1b0",
X"805383c0",
X"80085283",
X"c7e80851",
X"fed43f84",
X"3d0d0480",
X"3d0df9fc",
X"3f83c080",
X"08842981",
X"e39c0570",
X"0883c080",
X"0c51823d",
X"0d04ed3d",
X"0d804480",
X"43804280",
X"4180705a",
X"5bfdcc3f",
X"800b83c7",
X"d00c800b",
X"83c8840c",
X"81dff051",
X"e9c53f81",
X"800b83c8",
X"840c81df",
X"f451e9b7",
X"3f80d00b",
X"83c7d00c",
X"7830707a",
X"07802570",
X"872b83c8",
X"840c5155",
X"f8ed3f83",
X"c0800852",
X"81dffc51",
X"e9913f80",
X"f80b83c7",
X"d00c7881",
X"32703070",
X"72078025",
X"70872b83",
X"c8840c51",
X"56569ed2",
X"3f83c080",
X"085281e0",
X"8c51e8e7",
X"3f81a00b",
X"83c7d00c",
X"78823270",
X"30707207",
X"80257087",
X"2b83c884",
X"0c515656",
X"fec53f83",
X"c0800852",
X"81e09c51",
X"e8bd3f81",
X"c80b83c7",
X"d00c7883",
X"32703070",
X"72078025",
X"70872b83",
X"c8840c51",
X"5683c7e8",
X"085256ff",
X"b59f3f83",
X"c0800852",
X"81e0a451",
X"e88d3f82",
X"980b83c7",
X"d00c810b",
X"83c7d45b",
X"5883c7d0",
X"0883197a",
X"32703070",
X"72078025",
X"70872b83",
X"c8840c51",
X"578e3d70",
X"55ff1b54",
X"5757579c",
X"943f7970",
X"84055b08",
X"51ffb4d5",
X"3f745483",
X"c0800853",
X"775281e0",
X"ac51e7bf",
X"3fa81783",
X"c7d00c81",
X"18587785",
X"2e098106",
X"ffaf3883",
X"b80b83c7",
X"d00c7888",
X"32703070",
X"72078025",
X"70872b83",
X"c8840c51",
X"5656f7b9",
X"3f81e0bc",
X"5583c080",
X"08802e8f",
X"3883c7e4",
X"0851ffb4",
X"803f83c0",
X"80085574",
X"5281e0c4",
X"51e6ec3f",
X"84880b83",
X"c7d00c78",
X"89327030",
X"70720780",
X"2570872b",
X"83c8840c",
X"515681e0",
X"d05256e6",
X"ca3f84b0",
X"0b83c7d0",
X"0c788a32",
X"70307072",
X"07802570",
X"872b83c8",
X"840c5156",
X"81e0dc52",
X"56e6a83f",
X"85800b83",
X"c7d00c78",
X"8b327030",
X"70720780",
X"2570872b",
X"83c8840c",
X"515681e0",
X"f85256e6",
X"863f868d",
X"a051f7ef",
X"3f805291",
X"3d705255",
X"9f9e3f83",
X"5274519f",
X"973f6355",
X"7483e138",
X"61195978",
X"80258538",
X"74599139",
X"8c792586",
X"388c5983",
X"c539788b",
X"2683bf38",
X"78822b55",
X"81dadc15",
X"0804f58f",
X"3f83c080",
X"08615755",
X"75812e09",
X"81068938",
X"83c08008",
X"10559039",
X"75ff2e09",
X"81068838",
X"83c08008",
X"812c5590",
X"75258538",
X"90558839",
X"74802483",
X"38815574",
X"51f4e93f",
X"82f4399a",
X"d43f83c0",
X"80086105",
X"55748025",
X"85388055",
X"88398775",
X"25833887",
X"5574518e",
X"b73f82d2",
X"39f4d93f",
X"83c08008",
X"61055574",
X"80258538",
X"80558839",
X"86752583",
X"38865574",
X"51f4d23f",
X"82b03960",
X"87386280",
X"2e82a738",
X"83c39c08",
X"83c3980c",
X"ade50b83",
X"c3a00c83",
X"c7e80851",
X"d59d3ff9",
X"ca3f828a",
X"39605680",
X"76259838",
X"ad840b83",
X"c3a00c83",
X"c7c41570",
X"085255d4",
X"fe3f7408",
X"52923975",
X"80259238",
X"83c7c415",
X"0851ffb1",
X"823f8052",
X"fc1951b8",
X"3962802e",
X"81d03883",
X"c7c41570",
X"0883c7d4",
X"08720c83",
X"c7d40cfc",
X"1a705351",
X"558d843f",
X"83c08008",
X"5680518c",
X"fa3f83c0",
X"80085274",
X"5189933f",
X"75528051",
X"898c3f81",
X"99396055",
X"807525b8",
X"3883c3a8",
X"0883c398",
X"0cade50b",
X"83c3a00c",
X"83c7e408",
X"51d4883f",
X"83c7e408",
X"51d1a93f",
X"83c08008",
X"81ff0670",
X"5255f3b2",
X"3f74802e",
X"80e03881",
X"5580e339",
X"74802580",
X"d53883c7",
X"e40851ff",
X"aff13f80",
X"51f3933f",
X"80c43962",
X"802ebf38",
X"83c3a408",
X"83c3980c",
X"ade50b83",
X"c3a00c83",
X"c7ec0851",
X"d3b53f78",
X"892e0981",
X"068b3883",
X"c7ec0851",
X"f0f63f96",
X"39788a2e",
X"0981068e",
X"3883c7ec",
X"0851f0a3",
X"3f843962",
X"87387a80",
X"2ef8ae38",
X"80557483",
X"c0800c95",
X"3d0d04fe",
X"3d0d83c7",
X"f05180f7",
X"913ff2f6",
X"3f83c080",
X"08802e86",
X"38805181",
X"8a39f2fb",
X"3f83c080",
X"0880fe38",
X"f39b3f83",
X"c0800880",
X"2eb93881",
X"51f0d83f",
X"8051f2b1",
X"3fecd03f",
X"800b83c7",
X"d00cf7ce",
X"3f83c080",
X"0853ff0b",
X"83c7d00c",
X"eec33f72",
X"80cb3883",
X"c7cc3351",
X"f28b3f72",
X"51f0a83f",
X"80c039f2",
X"c33f83c0",
X"8008802e",
X"b5388151",
X"f0953f80",
X"51f1ee3f",
X"ec8d3fad",
X"840b83c3",
X"a00c83c7",
X"d40851d1",
X"ee3fff0b",
X"83c7d00c",
X"edff3f83",
X"c7d40852",
X"805186be",
X"3f8151f3",
X"b53f843d",
X"0d04fb3d",
X"0d805283",
X"c7f05180",
X"e6a03f80",
X"0b83c7cc",
X"34908080",
X"52868480",
X"8051ffb1",
X"d73f83c0",
X"80088197",
X"388a993f",
X"81e5bc51",
X"ffb6963f",
X"83c08008",
X"559c800a",
X"5480c080",
X"5381e180",
X"5283c080",
X"0851f591",
X"3f83c7e8",
X"085381e1",
X"90527451",
X"ffb0df3f",
X"83c08008",
X"8438f59f",
X"3f83c7ec",
X"085381e1",
X"9c527451",
X"ffb0c73f",
X"83c08008",
X"b638873d",
X"fc055484",
X"80805386",
X"a8808052",
X"83c7ec08",
X"51ffaed2",
X"3f83c080",
X"08933875",
X"8480802e",
X"09810689",
X"38810b83",
X"c7cc3487",
X"39800b83",
X"c7cc3483",
X"c7cc3351",
X"f08b3f81",
X"51f1f73f",
X"93ca3f81",
X"51f1ef3f",
X"8151fd8f",
X"3ffa3983",
X"c08c0802",
X"83c08c0c",
X"fb3d0d02",
X"81e1a80b",
X"83c39c0c",
X"81e1ac0b",
X"83c3940c",
X"81e1b00b",
X"83c3a80c",
X"81e1b40b",
X"83c3a40c",
X"83c08c08",
X"fc050c80",
X"0b83c7d4",
X"0b83c08c",
X"08f8050c",
X"83c08c08",
X"f4050cff",
X"aeda3f83",
X"c0800886",
X"05fc0683",
X"c08c08f0",
X"050c0283",
X"c08c08f0",
X"0508310d",
X"833d7083",
X"c08c08f8",
X"05087084",
X"0583c08c",
X"08f8050c",
X"0c51ffab",
X"a23f83c0",
X"8c08f405",
X"08810583",
X"c08c08f4",
X"050c83c0",
X"8c08f405",
X"08872e09",
X"8106ffab",
X"38869480",
X"8051e8b4",
X"3fff0b83",
X"c7d00c80",
X"0b83c884",
X"0c84d8c0",
X"0b83c880",
X"0c8151ec",
X"da3f8151",
X"ecff3f80",
X"51ecfa3f",
X"8151eda0",
X"3f8251ed",
X"c83f8051",
X"edf03f80",
X"51ee9a3f",
X"80d1a752",
X"8051dd98",
X"3ffccf3f",
X"83c08c08",
X"fc05080d",
X"800b83c0",
X"800c873d",
X"0d83c08c",
X"0c04803d",
X"0d81ff51",
X"800b83c8",
X"941234ff",
X"115170f4",
X"38823d0d",
X"04ff3d0d",
X"73703353",
X"51811133",
X"71347181",
X"1234833d",
X"0d04ff3d",
X"0d83cab0",
X"08a82e09",
X"81068b38",
X"83cac808",
X"83cab00c",
X"8739a80b",
X"83cab00c",
X"83cab008",
X"86057081",
X"ff065252",
X"d3a03f83",
X"3d0d04fb",
X"3d0d7779",
X"56568070",
X"71555552",
X"717525ac",
X"38721670",
X"33701470",
X"81ff0655",
X"51515171",
X"74278938",
X"81127081",
X"ff065351",
X"71811470",
X"83ffff06",
X"55525474",
X"7324d638",
X"7183c080",
X"0c873d0d",
X"04fb3d0d",
X"77568939",
X"f9e13f83",
X"51edc83f",
X"d4a73f83",
X"c0800880",
X"2eee3883",
X"cab00886",
X"057081ff",
X"065253d2",
X"ad3f810b",
X"9088d434",
X"f9b93f83",
X"51eda03f",
X"9088d433",
X"7081ff06",
X"55537380",
X"2eea3873",
X"862a7081",
X"06515372",
X"ffbe3873",
X"982b5380",
X"732480de",
X"38d3973f",
X"83c08008",
X"5583c080",
X"0880cf38",
X"74167582",
X"2b545490",
X"88c01333",
X"74348115",
X"5574852e",
X"098106e8",
X"38753383",
X"c8943481",
X"163383c8",
X"95348216",
X"3383c896",
X"34831633",
X"83c89734",
X"845283c8",
X"9451fe93",
X"3f83c080",
X"0881ff06",
X"84173355",
X"5372742e",
X"8738fdce",
X"3ffed139",
X"80e451ec",
X"923f873d",
X"0d04f43d",
X"0d7e6059",
X"55805d80",
X"75822b71",
X"83cab412",
X"0c83cacc",
X"175b5b57",
X"76793477",
X"772e83b7",
X"38765277",
X"51ffa9b6",
X"3f8e3dfc",
X"05549053",
X"83ca9c52",
X"7751ffa8",
X"f13f7c56",
X"75902e09",
X"81068393",
X"3883ca9c",
X"51fcde3f",
X"83ca9e51",
X"fcd73f83",
X"caa051fc",
X"d03f7683",
X"caac0c77",
X"51ffa6bd",
X"3f81df80",
X"5283c080",
X"0851c8d6",
X"3f83c080",
X"08812e09",
X"810680d4",
X"387683ca",
X"c40c820b",
X"83ca9c34",
X"ff960b83",
X"ca9d3477",
X"51ffa983",
X"3f83c080",
X"085583c0",
X"80087725",
X"883883c0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83ca9e34",
X"7483ca9f",
X"347683ca",
X"a034ff80",
X"0b83caa1",
X"34819039",
X"83ca9c33",
X"83ca9d33",
X"71882b07",
X"565b7483",
X"ffff2e09",
X"810680e8",
X"38fe800b",
X"83cac40c",
X"810b83ca",
X"ac0cff0b",
X"83ca9c34",
X"ff0b83ca",
X"9d347751",
X"ffa8903f",
X"83c08008",
X"83cad00c",
X"83c08008",
X"5583c080",
X"08802588",
X"3883c080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"ca9e3474",
X"83ca9f34",
X"7683caa0",
X"34ff800b",
X"83caa134",
X"810b83ca",
X"ab34a539",
X"7485962e",
X"09810680",
X"fe387583",
X"cac40c77",
X"51ffa7c4",
X"3f83caab",
X"3383c080",
X"08075574",
X"83caab34",
X"83caab33",
X"81065574",
X"802e8338",
X"845783ca",
X"a03383ca",
X"a1337188",
X"2b07565c",
X"7481802e",
X"098106a1",
X"3883ca9e",
X"3383ca9f",
X"3371882b",
X"07565bad",
X"80752787",
X"38768207",
X"579c3976",
X"81075796",
X"39748280",
X"2e098106",
X"87387683",
X"07578739",
X"7481ff26",
X"8a387783",
X"cab41b0c",
X"7679348e",
X"3d0d0480",
X"3d0d7284",
X"2983cab4",
X"05700883",
X"c0800c51",
X"823d0d04",
X"803d0d72",
X"7083c88c",
X"0c708429",
X"81e4f005",
X"700883ca",
X"c80c5151",
X"823d0d04",
X"fe3d0d81",
X"51de3f80",
X"0b83ca98",
X"0c800b83",
X"ca940cff",
X"0b83c890",
X"0ca80b83",
X"cab00cae",
X"51ccdb3f",
X"800b83ca",
X"b4545280",
X"73708405",
X"550c8112",
X"5271842e",
X"098106ef",
X"38843d0d",
X"04fe3d0d",
X"74028405",
X"96052253",
X"5371802e",
X"96387270",
X"81055433",
X"51cce63f",
X"ff127083",
X"ffff0651",
X"52e73984",
X"3d0d04fe",
X"3d0d0292",
X"05225382",
X"ac51e787",
X"3f80c351",
X"ccc33f81",
X"9651e6fb",
X"3f725283",
X"c89451ff",
X"b43f7252",
X"83c89451",
X"f8cd3f83",
X"c0800881",
X"ff0651cc",
X"a03f843d",
X"0d04ffb1",
X"3d0d80d1",
X"3df80551",
X"f8f73f83",
X"ca980881",
X"0583ca98",
X"0c80cf3d",
X"33cf1170",
X"81ff0651",
X"56567483",
X"2688e638",
X"758f06ff",
X"05567583",
X"c890082e",
X"9b387583",
X"26963875",
X"83c8900c",
X"75842983",
X"cab40570",
X"08535575",
X"51f9fb3f",
X"80762488",
X"c2387584",
X"2983cab4",
X"05557408",
X"802e88b3",
X"3883c890",
X"08842983",
X"cab40570",
X"08028805",
X"82b90533",
X"525b5574",
X"80d22e84",
X"b0387480",
X"d2249038",
X"74bf2e9c",
X"387480d0",
X"2e81d538",
X"87f23974",
X"80d32e80",
X"d3387480",
X"d72e81c4",
X"3887e139",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"055656cb",
X"9c3f80c1",
X"51cad63f",
X"f6983f83",
X"cacb3383",
X"c8943481",
X"5283c894",
X"51cbf33f",
X"8151fde7",
X"3f748b38",
X"83cac808",
X"83cab00c",
X"8739a80b",
X"83cab00c",
X"cae73f80",
X"c151caa1",
X"3ff5e33f",
X"900b83ca",
X"ab338106",
X"56567480",
X"2e833898",
X"5683caa0",
X"3383caa1",
X"3371882b",
X"07565974",
X"81802e09",
X"81069c38",
X"83ca9e33",
X"83ca9f33",
X"71882b07",
X"5657ad80",
X"75278c38",
X"75818007",
X"56853975",
X"a0075675",
X"83c89434",
X"ff0b83c8",
X"9534e00b",
X"83c89634",
X"800b83c8",
X"97348452",
X"83c89451",
X"cae83f84",
X"51869b39",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"055659c9",
X"dc3f7951",
X"ffa1f13f",
X"83c08008",
X"802e8a38",
X"80ce51c9",
X"883f85f1",
X"3980c151",
X"c8ff3fc9",
X"f03fc8a9",
X"3f83cac4",
X"08588375",
X"259b3883",
X"caa03383",
X"caa13371",
X"882b07fc",
X"1771297a",
X"05838005",
X"5a51578d",
X"39748180",
X"2918ff80",
X"05588180",
X"57805676",
X"762e9238",
X"c8db3f83",
X"c0800883",
X"c8941734",
X"811656eb",
X"39c8ca3f",
X"83c08008",
X"81ff0677",
X"5383c894",
X"5256f4bf",
X"3f83c080",
X"0881ff06",
X"5575752e",
X"09810681",
X"95389451",
X"e2c53fc8",
X"c43f80c1",
X"51c7fe3f",
X"c8ef3f77",
X"527951ff",
X"a0843f80",
X"5e80d13d",
X"fdf40554",
X"765383c8",
X"94527951",
X"ff9e913f",
X"0282b905",
X"33558159",
X"7480d72e",
X"09810680",
X"c5387752",
X"7951ff9f",
X"d53f80d1",
X"3dfdf005",
X"5476538f",
X"3d70537a",
X"5258ff9f",
X"8d3f8056",
X"76762ea2",
X"38751883",
X"c8941733",
X"71337072",
X"32703070",
X"80257030",
X"7f06811d",
X"5d5f5151",
X"51525b55",
X"db3982ac",
X"51e1c03f",
X"78802e86",
X"3880c351",
X"843980ce",
X"51c6f23f",
X"c7e33fc6",
X"9c3f83d8",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055955",
X"80705d59",
X"80e451e1",
X"8a3fc789",
X"3f80c151",
X"c6c33f83",
X"caac0879",
X"2e82d638",
X"83cad008",
X"80fc0555",
X"80fd5274",
X"5185c13f",
X"83c08008",
X"5b778224",
X"b238ff18",
X"70872b83",
X"ffff8006",
X"81e3bc05",
X"83c89459",
X"57558180",
X"55757081",
X"05573377",
X"70810559",
X"34ff1570",
X"81ff0651",
X"5574ea38",
X"82853977",
X"82e82e81",
X"a3387782",
X"e92e0981",
X"0681aa38",
X"78587787",
X"32703070",
X"72078025",
X"7a8a3270",
X"30707207",
X"80257307",
X"53545a51",
X"57557580",
X"2e973878",
X"78269238",
X"a00b83c8",
X"941a3481",
X"197081ff",
X"065a55eb",
X"39811870",
X"81ff0659",
X"558a7827",
X"ffbc388f",
X"5883c88f",
X"183383c8",
X"941934ff",
X"187081ff",
X"06595577",
X"8426ea38",
X"9058800b",
X"83c89419",
X"34811870",
X"81ff0670",
X"982b5259",
X"55748025",
X"e93880c6",
X"557a858f",
X"24843880",
X"c2557483",
X"c8943480",
X"f10b83c8",
X"9734810b",
X"83c89834",
X"7a83c895",
X"347a882c",
X"557483c8",
X"963480cb",
X"3982f078",
X"2580c438",
X"7780fd29",
X"fd97d305",
X"527951ff",
X"9cb03f80",
X"d13dfdec",
X"055480fd",
X"5383c894",
X"527951ff",
X"9be83f7b",
X"81195956",
X"7580fc24",
X"83387858",
X"77882c55",
X"7483c991",
X"347783c9",
X"92347583",
X"c9933481",
X"805980cc",
X"3983cac4",
X"08578378",
X"259b3883",
X"caa03383",
X"caa13371",
X"882b07fc",
X"1a712979",
X"05838005",
X"5951598d",
X"39778180",
X"2917ff80",
X"05578180",
X"59765279",
X"51ff9bbe",
X"3f80d13d",
X"fdec0554",
X"785383c8",
X"94527951",
X"ff9af73f",
X"7851f6bf",
X"3fc4863f",
X"c2bf3f8b",
X"3983ca94",
X"08810583",
X"ca940c80",
X"d13d0d04",
X"f6e03ffc",
X"39fc3d0d",
X"76787184",
X"2983cab4",
X"05700851",
X"53535370",
X"9e3880ce",
X"723480cf",
X"0b811334",
X"80ce0b82",
X"133480c5",
X"0b831334",
X"70841334",
X"80e73983",
X"cacc1333",
X"5480d272",
X"3473822a",
X"70810651",
X"5180cf53",
X"70843880",
X"d7537281",
X"1334a00b",
X"82133473",
X"83065170",
X"812e9e38",
X"70812488",
X"3870802e",
X"8f389f39",
X"70822e92",
X"3870832e",
X"92389339",
X"80d8558e",
X"3980d355",
X"893980cd",
X"55843980",
X"c4557483",
X"133480c4",
X"0b841334",
X"800b8513",
X"34863d0d",
X"0483c88c",
X"0883c080",
X"0c04803d",
X"0d83c88c",
X"08842981",
X"e5900570",
X"0883c080",
X"0c51823d",
X"0d04fc3d",
X"0d767853",
X"54815380",
X"55873971",
X"10731054",
X"52737226",
X"5172802e",
X"a7387080",
X"2e863871",
X"8025e838",
X"72802e98",
X"38717426",
X"89387372",
X"31757407",
X"56547281",
X"2a72812a",
X"5353e539",
X"73517883",
X"38745170",
X"83c0800c",
X"863d0d04",
X"fe3d0d80",
X"53755274",
X"51ffa33f",
X"843d0d04",
X"fe3d0d81",
X"53755274",
X"51ff933f",
X"843d0d04",
X"fb3d0d77",
X"79555580",
X"56747625",
X"86387430",
X"55815673",
X"80258838",
X"73307681",
X"32575480",
X"53735274",
X"51fee73f",
X"83c08008",
X"5475802e",
X"873883c0",
X"80083054",
X"7383c080",
X"0c873d0d",
X"04fa3d0d",
X"787a5755",
X"80577477",
X"25863874",
X"30558157",
X"759f2c54",
X"81537574",
X"32743152",
X"7451feaa",
X"3f83c080",
X"08547680",
X"2e873883",
X"c0800830",
X"547383c0",
X"800c883d",
X"0d04fc3d",
X"0d765580",
X"750c800b",
X"84160c80",
X"0b88160c",
X"800b8c16",
X"0c83c7f0",
X"5180dd9a",
X"3f87a680",
X"337081ff",
X"06707184",
X"2a065151",
X"52d9c33f",
X"71812a81",
X"32728132",
X"71810671",
X"81063184",
X"180c5454",
X"71832a81",
X"3272822a",
X"81327081",
X"06727131",
X"780c5153",
X"5387a090",
X"3387a091",
X"337081ff",
X"06707306",
X"81328106",
X"88190c51",
X"535383c0",
X"8008802e",
X"80c23883",
X"c0800881",
X"2a708106",
X"83c08008",
X"81063184",
X"170c5283",
X"c0800883",
X"2a83c080",
X"08822a71",
X"81067181",
X"0631770c",
X"535383c0",
X"8008842a",
X"81068816",
X"0c83c080",
X"08852a81",
X"068c160c",
X"863d0d04",
X"fe3d0d74",
X"76545271",
X"51feb33f",
X"72812ea2",
X"38817326",
X"8d387282",
X"2ea83872",
X"832e9c38",
X"e6397108",
X"e2388412",
X"08dd3888",
X"1208d838",
X"a5398812",
X"08812e9e",
X"38913988",
X"1208812e",
X"95387108",
X"91388412",
X"088c388c",
X"1208812e",
X"098106ff",
X"b238843d",
X"0d04fb3d",
X"0d780284",
X"059f0533",
X"5556800b",
X"81dcf856",
X"5381732b",
X"74065271",
X"802e8338",
X"81527470",
X"82055622",
X"7073902b",
X"0790809c",
X"0c518113",
X"5372882e",
X"098106d9",
X"38805383",
X"cad81333",
X"517081ff",
X"2eb23870",
X"1081db98",
X"05702255",
X"51807317",
X"70337010",
X"81db9805",
X"70225151",
X"51525273",
X"712e9138",
X"81125271",
X"862e0981",
X"06f13873",
X"90809c0c",
X"81135372",
X"862e0981",
X"06ffb838",
X"80537216",
X"70335151",
X"7081ff2e",
X"94387010",
X"81db9805",
X"70227084",
X"80800790",
X"809c0c51",
X"51811353",
X"72862e09",
X"8106d738",
X"80537216",
X"51703383",
X"cad81434",
X"81135372",
X"862e0981",
X"06ec3887",
X"3d0d0404",
X"ff3d0d74",
X"0284058f",
X"05335252",
X"70883871",
X"9080940c",
X"8e397081",
X"2e098106",
X"86387190",
X"80980c83",
X"3d0d04fb",
X"3d0d029f",
X"05337998",
X"2b70982c",
X"7c982b70",
X"982c83ca",
X"f4157033",
X"70982b70",
X"982c5158",
X"5c5a5155",
X"51545470",
X"732e0981",
X"06943883",
X"cad41433",
X"70982b70",
X"982c5152",
X"5670722e",
X"b1387275",
X"347183ca",
X"d4153483",
X"cad53383",
X"caf53371",
X"982b7190",
X"2b0783ca",
X"d4337088",
X"2b720783",
X"caf43371",
X"079080b8",
X"0c525953",
X"5452873d",
X"0d04fe3d",
X"0d748111",
X"33713371",
X"882b0783",
X"c0800c53",
X"51843d0d",
X"0483cae0",
X"3383c080",
X"0c04f53d",
X"0d02bb05",
X"33028405",
X"bf053302",
X"880580c3",
X"0533028c",
X"0580c605",
X"22665c5a",
X"5e5c567a",
X"557b5489",
X"53a1527d",
X"5180d2fb",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8d3d0d04",
X"83c08c08",
X"0283c08c",
X"0cf53d0d",
X"83c08c08",
X"88050883",
X"c08c088f",
X"053383c0",
X"8c089205",
X"22028c05",
X"73900583",
X"c08c08e8",
X"050c83c0",
X"8c08f805",
X"0c83c08c",
X"08f0050c",
X"83c08c08",
X"ec050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"f0050883",
X"c08c08e0",
X"050c83c0",
X"8c08fc05",
X"0c83c08c",
X"08f00508",
X"89278a38",
X"890b83c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"860587ff",
X"fc0683c0",
X"8c08e005",
X"0c0283c0",
X"8c08e005",
X"08310d85",
X"3d705583",
X"c08c08ec",
X"05085483",
X"c08c08f0",
X"05085383",
X"c08c08f4",
X"05085283",
X"c08c08e4",
X"050c80dc",
X"d43f83c0",
X"800881ff",
X"0683c08c",
X"08e40508",
X"83c08c08",
X"ec050c83",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08802e8c",
X"3883c08c",
X"08f80508",
X"0d89c839",
X"83c08c08",
X"f0050880",
X"2e89a638",
X"83c08c08",
X"ec050881",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"842ea938",
X"840b83c0",
X"8c08e005",
X"082588c7",
X"3883c08c",
X"08e00508",
X"852e859b",
X"3883c08c",
X"08e00508",
X"a12e87ad",
X"3888ac39",
X"800b83c0",
X"8c08ec05",
X"08850533",
X"83c08c08",
X"e0050c83",
X"c08c08fc",
X"050c83c0",
X"8c08e005",
X"08832e09",
X"81068883",
X"3883c08c",
X"08e80508",
X"81053383",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08812687",
X"e638810b",
X"83c08c08",
X"e0050880",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08fc050c",
X"83c08c08",
X"ec050882",
X"053383c0",
X"8c08e005",
X"08870534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088b0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08e005",
X"088c0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088d0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08e005",
X"088e0523",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088a0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"08057094",
X"0508fcff",
X"ff067194",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08ec0508",
X"86053383",
X"c08c08e0",
X"050c83c0",
X"8c08f405",
X"0c83c08c",
X"08e00508",
X"83c08c08",
X"fc05082e",
X"098106b6",
X"3883c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08fc0508",
X"83c08c08",
X"e005088b",
X"053483c0",
X"8c08ec05",
X"08870533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508812e",
X"8f3883c0",
X"8c08e005",
X"08822eb7",
X"38848c39",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"820b83c0",
X"8c08e005",
X"088a0534",
X"83d93983",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c83",
X"c08c08fc",
X"050883c0",
X"8c08e005",
X"088a0534",
X"83a13983",
X"c08c08fc",
X"0508802e",
X"83953883",
X"c08c08ec",
X"05088305",
X"33830683",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08832e09",
X"810682f3",
X"3883c08c",
X"08ec0508",
X"82053370",
X"982b83c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"83c08c08",
X"e0050880",
X"2582cc38",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"83c08c08",
X"ec050886",
X"053383c0",
X"8c08e005",
X"0880d605",
X"3483c08c",
X"08e00508",
X"840583c0",
X"8c08ec05",
X"08820533",
X"8f0683c0",
X"8c08e405",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"e4050883",
X"c08c08e0",
X"05083483",
X"c08c08ec",
X"05088405",
X"3383c08c",
X"08e00508",
X"81053480",
X"0b83c08c",
X"08e00508",
X"82053483",
X"c08c08e0",
X"050808ff",
X"83ff0682",
X"800783c0",
X"8c08e005",
X"080c83c0",
X"8c08e805",
X"08810533",
X"810583c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"83c08c08",
X"e8050881",
X"05348183",
X"3983c08c",
X"08fc0508",
X"802e80f7",
X"3883c08c",
X"08ec0508",
X"86053383",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08a22e09",
X"810680d7",
X"3883c08c",
X"08ec0508",
X"88053383",
X"c08c08ec",
X"05088705",
X"33718280",
X"290583c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c52",
X"83c08c08",
X"e4050c83",
X"c08c08f4",
X"050c83c0",
X"8c08e405",
X"0883c08c",
X"08e00508",
X"88052383",
X"c08c08ec",
X"05083383",
X"c08c08f0",
X"05087131",
X"7083ffff",
X"0683c08c",
X"08f0050c",
X"83c08c08",
X"e0050c83",
X"c08c08ec",
X"05080583",
X"c08c08ec",
X"050cf6d0",
X"3983c08c",
X"08f80508",
X"0d83c08c",
X"08f00508",
X"83c08c08",
X"e0050c83",
X"c08c08f8",
X"05080d83",
X"c08c08e0",
X"050883c0",
X"800c8d3d",
X"0d83c08c",
X"0c0483c0",
X"8c080283",
X"c08c0ce6",
X"3d0d83c0",
X"8c088805",
X"08028405",
X"83c08c08",
X"e8050c83",
X"c08c08d4",
X"050c800b",
X"83cafc34",
X"83c08c08",
X"d4050890",
X"0583c08c",
X"08c0050c",
X"800b83c0",
X"8c08c005",
X"0834800b",
X"83c08c08",
X"c0050881",
X"0534800b",
X"83c08c08",
X"c4050c83",
X"c08c08c4",
X"050880d8",
X"2983c08c",
X"08c00508",
X"0583c08c",
X"08ffb405",
X"0c800b83",
X"c08c08ff",
X"b4050880",
X"d8050c83",
X"c08c08ff",
X"b4050884",
X"0583c08c",
X"08ffb405",
X"0c83c08c",
X"08c40508",
X"83c08c08",
X"ffb40508",
X"34880b83",
X"c08c08ff",
X"b4050881",
X"0534800b",
X"83c08c08",
X"ffb40508",
X"82053483",
X"c08c08ff",
X"b4050808",
X"ffa1ff06",
X"a0800783",
X"c08c08ff",
X"b405080c",
X"83c08c08",
X"c4050881",
X"057081ff",
X"0683c08c",
X"08c4050c",
X"83c08c08",
X"ffb4050c",
X"810b83c0",
X"8c08c405",
X"0827fedb",
X"3883c08c",
X"08ec0570",
X"5483c08c",
X"08c8050c",
X"925283c0",
X"8c08d405",
X"085180cf",
X"fb3f83c0",
X"800881ff",
X"067083c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"05088eb4",
X"3883c08c",
X"08f40551",
X"f18c3f83",
X"c0800883",
X"ffff0683",
X"c08c08f6",
X"055283c0",
X"8c08e405",
X"0cf0f33f",
X"83c08008",
X"83ffff06",
X"83c08c08",
X"fd053383",
X"c08c08ff",
X"b8050883",
X"c08c08c4",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08dc05",
X"0c83c08c",
X"08c40508",
X"83c08c08",
X"ffbc0508",
X"2780fe38",
X"83c08c08",
X"c8050854",
X"83c08c08",
X"c4050853",
X"895283c0",
X"8c08d405",
X"085180cf",
X"803f83c0",
X"800881ff",
X"0683c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"0880f238",
X"83c08c08",
X"ee0551ef",
X"f13f83c0",
X"800883ff",
X"ff065383",
X"c08c08c4",
X"05085283",
X"c08c08d4",
X"050851f0",
X"b33f83c0",
X"8c08c405",
X"08810570",
X"81ff0683",
X"c08c08c4",
X"050c83c0",
X"8c08ffb4",
X"050cfef1",
X"3983c08c",
X"08c00508",
X"81053383",
X"c08c08ff",
X"b4050c81",
X"db0b83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb4",
X"0508802e",
X"8caa3894",
X"3983c08c",
X"08ffb805",
X"0883c08c",
X"08ffbc05",
X"0c8c9539",
X"83c08c08",
X"f1053352",
X"83c08c08",
X"d4050851",
X"80cdfe3f",
X"800b83c0",
X"8c08c005",
X"08810533",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"c4050c83",
X"c08c08c4",
X"050883c0",
X"8c08ffb4",
X"0508278a",
X"b03883c0",
X"8c08c405",
X"0880d829",
X"7083c08c",
X"08c00508",
X"05708805",
X"70830533",
X"83c08c08",
X"cc050c83",
X"c08c08c8",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08d805",
X"0c83c08c",
X"08cc0508",
X"87f03883",
X"c08c08c8",
X"05082202",
X"84057186",
X"0587fffc",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"ffb8050c",
X"0283c08c",
X"08ffb405",
X"08310d89",
X"3d705983",
X"c08c08ff",
X"b8050858",
X"83c08c08",
X"ffbc0508",
X"87053357",
X"83c08c08",
X"ffb4050c",
X"a25583c0",
X"8c08cc05",
X"08548653",
X"81815283",
X"c08c08d4",
X"05085180",
X"c0cd3f83",
X"c0800881",
X"ff0683c0",
X"8c08d005",
X"0c83c08c",
X"08d00508",
X"81c13883",
X"c08c08ff",
X"bc050896",
X"055383c0",
X"8c08ffb8",
X"05085283",
X"c08c08ff",
X"b4050851",
X"a4803f83",
X"c0800881",
X"ff0683c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb4",
X"0508802e",
X"81853883",
X"c08c08ff",
X"bc050894",
X"0583c08c",
X"08ffbc05",
X"08960533",
X"70862a83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08cc",
X"050c83c0",
X"8c08ffb4",
X"0508832e",
X"09810680",
X"c63883c0",
X"8c08ffb4",
X"050883c0",
X"8c08c805",
X"08820534",
X"83cae033",
X"70810583",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b4050883",
X"cae03483",
X"c08c08ff",
X"b8050883",
X"c08c08cc",
X"05083483",
X"c08c08e0",
X"05080d83",
X"c08c08d0",
X"050881ff",
X"0683c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"08fbfe38",
X"83c08c08",
X"d8050883",
X"c08c08c0",
X"05080588",
X"05708205",
X"335183c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb4",
X"0508832e",
X"09810680",
X"e33883c0",
X"8c08ffb8",
X"050883c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb4",
X"05088105",
X"7081ff06",
X"5183c08c",
X"08ffb405",
X"0c810b83",
X"c08c08ff",
X"b4050827",
X"dd38800b",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb40508",
X"81057081",
X"ff065183",
X"c08c08ff",
X"b4050c97",
X"0b83c08c",
X"08ffb405",
X"0827dd38",
X"83c08c08",
X"e4050880",
X"f9327030",
X"70802551",
X"5183c08c",
X"08ffb405",
X"0c83c08c",
X"08dc0508",
X"912e0981",
X"0680f938",
X"83c08c08",
X"ffb40508",
X"802e80ec",
X"3883c08c",
X"08c40508",
X"80e23885",
X"0b83c08c",
X"08c00508",
X"a60534a0",
X"0b83c08c",
X"08c00508",
X"a7053485",
X"0b83c08c",
X"08c00508",
X"a8053480",
X"c00b83c0",
X"8c08c005",
X"08a90534",
X"860b83c0",
X"8c08c005",
X"08aa0534",
X"900b83c0",
X"8c08c005",
X"08ab0534",
X"860b83c0",
X"8c08c005",
X"08ac0534",
X"a00b83c0",
X"8c08c005",
X"08ad0534",
X"83c08c08",
X"e4050889",
X"d8327030",
X"70802551",
X"5183c08c",
X"08ffb405",
X"0c83c08c",
X"08dc0508",
X"83edec2e",
X"09810680",
X"f6388170",
X"83c08c08",
X"ffb40508",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb405",
X"08802e80",
X"ce3883c0",
X"8c08c405",
X"0880c438",
X"840b83c0",
X"8c08c005",
X"08aa0534",
X"80c00b83",
X"c08c08c0",
X"0508ab05",
X"34840b83",
X"c08c08c0",
X"0508ac05",
X"34900b83",
X"c08c08c0",
X"0508ad05",
X"3483c08c",
X"08ffb805",
X"0883c08c",
X"08c00508",
X"8c053483",
X"c08c08e4",
X"050880f9",
X"32703070",
X"80255151",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"dc050886",
X"2e098106",
X"80c33881",
X"7083c08c",
X"08ffb405",
X"080683c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb4",
X"0508802e",
X"9c3883c0",
X"8c08c405",
X"08933883",
X"c08c08ff",
X"b8050883",
X"c08c08c0",
X"05088d05",
X"3483c08c",
X"08e40508",
X"b4b43270",
X"30708025",
X"515183c0",
X"8c08ffb4",
X"050c83c0",
X"8c08dc05",
X"0890892e",
X"098106a2",
X"3883c08c",
X"08ffb405",
X"08802e96",
X"3883c08c",
X"08c40508",
X"8d38820b",
X"83c08c08",
X"c005088d",
X"053483c0",
X"8c08c405",
X"0880d829",
X"83c08c08",
X"c0050805",
X"70840570",
X"83053383",
X"c08c08ff",
X"b4050c83",
X"c08c08c8",
X"050c83c0",
X"8c08ffbc",
X"050c8058",
X"805783c0",
X"8c08ffb4",
X"05085680",
X"5580548a",
X"53a15283",
X"c08c08d4",
X"050851b8",
X"fe3f83c0",
X"800881ff",
X"06703070",
X"9f2a5183",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b80508a0",
X"2e8c3883",
X"c08c08ff",
X"b40508f5",
X"f83883c0",
X"8c08ffbc",
X"05088b05",
X"3383c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb405",
X"08802eb3",
X"3883c08c",
X"08c80508",
X"83053383",
X"c08c08ff",
X"b4050c80",
X"58805783",
X"c08c08ff",
X"b4050856",
X"80558054",
X"8b53a152",
X"83c08c08",
X"d4050851",
X"b7f93f83",
X"c08c08c4",
X"05088105",
X"7081ff06",
X"83c08c08",
X"c0050881",
X"05335283",
X"c08c08c4",
X"050c83c0",
X"8c08ffb4",
X"050cf5bf",
X"39800b83",
X"c08c08c4",
X"050c83c0",
X"8c08c405",
X"0880d829",
X"83c08c08",
X"d4050805",
X"709a0533",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb40508",
X"822e0981",
X"06a93883",
X"cafc5681",
X"55805483",
X"c08c08ff",
X"b4050853",
X"83c08c08",
X"ffb80508",
X"97053352",
X"83c08c08",
X"d4050851",
X"e3c03f83",
X"c08c08c4",
X"05088105",
X"7081ff06",
X"83c08c08",
X"c4050c83",
X"c08c08ff",
X"b4050c81",
X"0b83c08c",
X"08c40508",
X"27fefb38",
X"810b83c0",
X"8c08c005",
X"0834800b",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"e805080d",
X"83c08c08",
X"ffbc0508",
X"83c0800c",
X"9c3d0d83",
X"c08c0c04",
X"f43d0d90",
X"1f59800b",
X"811a3355",
X"5b7a7427",
X"81ad387a",
X"80d82919",
X"8a113355",
X"5573832e",
X"09810681",
X"88389415",
X"33578052",
X"7651e0f8",
X"3f805380",
X"527651e1",
X"963faaed",
X"3f83c080",
X"085c8058",
X"7781c429",
X"1c871133",
X"55557380",
X"2e80c038",
X"740881db",
X"8c2e0981",
X"06b53880",
X"755b5675",
X"80d8291a",
X"9a113355",
X"5573832e",
X"09810692",
X"38a41570",
X"33555576",
X"74278738",
X"ff145473",
X"75348116",
X"7081ff06",
X"57548176",
X"27d13881",
X"187081ff",
X"0659548f",
X"7827ffa4",
X"3883cae0",
X"33ff0554",
X"7383cae0",
X"34811b70",
X"81ff0681",
X"1b335f5c",
X"547c7b26",
X"fed53880",
X"0b83c080",
X"0c8e3d0d",
X"0483c08c",
X"080283c0",
X"8c0ce63d",
X"0d83c08c",
X"08880508",
X"02840571",
X"90057033",
X"7083c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"dc050c83",
X"c08c08e0",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"96963880",
X"0b83c08c",
X"08c80508",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08d0",
X"050c83c0",
X"8c08d005",
X"0883c08c",
X"08ffa405",
X"082595de",
X"3883c08c",
X"08d00508",
X"80d82983",
X"c08c08c8",
X"05080584",
X"05708605",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffa405",
X"08802e94",
X"ea38a893",
X"3f83c08c",
X"08ffbc05",
X"0880d405",
X"0883c080",
X"082694d3",
X"380283c0",
X"8c08ffbc",
X"05088105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08d8050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"fc052383",
X"c08c08ff",
X"a4050886",
X"0583fc06",
X"83c08c08",
X"ffa4050c",
X"0283c08c",
X"08ffa405",
X"08310d85",
X"3d705583",
X"c08c08fc",
X"055483c0",
X"8c08ffbc",
X"05085383",
X"c08c08e0",
X"05085283",
X"c08c08c4",
X"050cafeb",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"939c3883",
X"c08c08ff",
X"bc050887",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"80d53883",
X"c08c08ff",
X"bc050886",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508822e",
X"098106b3",
X"3883c08c",
X"08fc0522",
X"83c08c08",
X"ffa4050c",
X"870b83c0",
X"8c08ffa4",
X"05082797",
X"3883c08c",
X"08c40508",
X"82055283",
X"c08c08c4",
X"05083351",
X"dacc3f83",
X"c08c08ff",
X"bc050886",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508832e",
X"09810692",
X"853883c0",
X"8c08ffbc",
X"05089205",
X"70820533",
X"83c08c08",
X"fc052283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08c0",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffa8",
X"05082691",
X"c538800b",
X"83c08c08",
X"e4050c80",
X"0b83c08c",
X"08ffb005",
X"0c83c08c",
X"08ffb005",
X"081083c0",
X"8c0805f8",
X"0583c08c",
X"08ffb005",
X"08842983",
X"c08c08ff",
X"b0050810",
X"0583c08c",
X"08c00508",
X"05708405",
X"703383c0",
X"8c08c405",
X"08057033",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffb80508",
X"2383c08c",
X"08ffa805",
X"08810533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"902e0981",
X"06be3883",
X"c08c08ff",
X"a8050833",
X"83c08c08",
X"c4050805",
X"81057033",
X"70828029",
X"83c08c08",
X"ffb40508",
X"05515183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"b8050823",
X"83c08c08",
X"ffac0508",
X"86052283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a80508a2",
X"3883c08c",
X"08ffac05",
X"08880522",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"81ff2e80",
X"e53883c0",
X"8c08ffb8",
X"05082270",
X"83c08c08",
X"ffa80508",
X"31708280",
X"29713183",
X"c08c08ff",
X"ac050888",
X"05227083",
X"c08c08ff",
X"a8050831",
X"70733553",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffb805",
X"082383c0",
X"8c08ffb0",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa4050c",
X"810b83c0",
X"8c08ffb0",
X"050827fc",
X"e03883c0",
X"8c08f805",
X"2283c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08bf2691",
X"3883c08c",
X"08e40508",
X"820783c0",
X"8c08e405",
X"0c81c00b",
X"83c08c08",
X"ffa40508",
X"27913883",
X"c08c08e4",
X"05088107",
X"83c08c08",
X"e4050c83",
X"c08c08fa",
X"052283c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508bf26",
X"913883c0",
X"8c08e405",
X"08880783",
X"c08c08e4",
X"050c81c0",
X"0b83c08c",
X"08ffa405",
X"08279138",
X"83c08c08",
X"e4050884",
X"0783c08c",
X"08e4050c",
X"800b83c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffb0",
X"05081083",
X"c08c08c0",
X"05080570",
X"90057033",
X"83c08c08",
X"c4050805",
X"70337281",
X"05337072",
X"06515351",
X"83c08c08",
X"ffa8050c",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e9b",
X"38900b83",
X"c08c08ff",
X"b005082b",
X"83c08c08",
X"e4050807",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"b0050881",
X"057081ff",
X"0683c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa405",
X"0c970b83",
X"c08c08ff",
X"b0050827",
X"fef43883",
X"c08c08ff",
X"bc050890",
X"053383c0",
X"8c08e405",
X"0883c08c",
X"08ffa405",
X"0c83c08c",
X"08c0050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffbc0508",
X"8c05082e",
X"85e03883",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"bc05088c",
X"050c83c0",
X"8c08ffbc",
X"05088905",
X"3383c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa805",
X"08802e85",
X"9a3883c0",
X"8c08e405",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffa40508",
X"8f0683c0",
X"8c08e405",
X"0c83c08c",
X"08ffb005",
X"0c83c08c",
X"08d4050c",
X"83c08c08",
X"ffa80508",
X"822e0981",
X"0681c238",
X"800b83c0",
X"8c08ffa4",
X"0508862a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffa80508",
X"2e8c3881",
X"c00b83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffb0",
X"0508872a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9438",
X"83c08c08",
X"ffa80508",
X"81903283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"b0050884",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e94",
X"3883c08c",
X"08ffa805",
X"0880d032",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffb00508",
X"83c08c08",
X"ffa80508",
X"3283c08c",
X"08ffb005",
X"0c800b83",
X"c08c08f0",
X"050c800b",
X"83c08c08",
X"f4052380",
X"0b81dd88",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffb805",
X"082e82d3",
X"3883c08c",
X"08f00581",
X"dd880b83",
X"c08c08ff",
X"ac050c83",
X"c08c08cc",
X"050c83c0",
X"8c08ffac",
X"05083383",
X"c08c08ff",
X"ac050881",
X"05338172",
X"2b81722b",
X"077083c0",
X"8c08ffb0",
X"05080652",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffa80508",
X"2e098106",
X"81be3883",
X"c08c08ff",
X"b8050885",
X"2680f638",
X"83c08c08",
X"ffac0508",
X"82053370",
X"81ff0683",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050880",
X"2e80ca38",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"ffb80508",
X"81057081",
X"ff0683c0",
X"8c08cc05",
X"08730553",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffa40508",
X"3483c08c",
X"08ffac05",
X"08830533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9d38",
X"810b83c0",
X"8c08ffa4",
X"05082b83",
X"c08c08d4",
X"05080807",
X"83c08c08",
X"d405080c",
X"83c08c08",
X"ffac0508",
X"84057033",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa40508",
X"fdc83883",
X"c08c08f0",
X"05528051",
X"ce883f83",
X"c08c08e4",
X"05085283",
X"c08c08c0",
X"050851cf",
X"c33f83c0",
X"8c08fb05",
X"33708180",
X"0a29810a",
X"0570982c",
X"5583c08c",
X"08ffa405",
X"0c83c08c",
X"08f90533",
X"7081800a",
X"29810a05",
X"70982c55",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"c0050853",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa8050c",
X"cf993f83",
X"c08c08ff",
X"bc050888",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"84e03883",
X"c08c08ff",
X"bc050890",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"05088126",
X"84c03880",
X"7081ddc8",
X"0b81ddc8",
X"0b810533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffb40508",
X"2e81ae38",
X"83c08c08",
X"ffac0508",
X"842983c0",
X"8c08ffa8",
X"05080570",
X"3383c08c",
X"08c40508",
X"05703372",
X"81053370",
X"72065153",
X"5183c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802eaa",
X"38810b83",
X"c08c08ff",
X"ac05082b",
X"83c08c08",
X"ffb40508",
X"077083ff",
X"ff0683c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffac",
X"05088105",
X"7081ff06",
X"81ddc871",
X"84297105",
X"70810533",
X"515383c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508fed4",
X"3883c08c",
X"08ffbc05",
X"088a0522",
X"83c08c08",
X"c0050c83",
X"c08c08ff",
X"b4050883",
X"c08c08c0",
X"05082e82",
X"ad38800b",
X"83c08c08",
X"e8050c80",
X"0b83c08c",
X"08ec0523",
X"807083c0",
X"8c08e805",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffb0050c",
X"81af3983",
X"c08c08ff",
X"b4050883",
X"c08c08ff",
X"ac05082c",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e80e7",
X"3883c08c",
X"08ffb005",
X"0883c08c",
X"08ffb005",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"b8050873",
X"0583c08c",
X"08ffbc05",
X"08900533",
X"83c08c08",
X"ffac0508",
X"84290553",
X"5383c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa805",
X"0881ddca",
X"053383c0",
X"8c08ffa4",
X"05083483",
X"c08c08ff",
X"ac050881",
X"057081ff",
X"0683c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa405",
X"0c8f0b83",
X"c08c08ff",
X"ac050827",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb00508",
X"85268c38",
X"83c08c08",
X"ffa40508",
X"fea93883",
X"c08c08e8",
X"05528051",
X"c8b83f83",
X"c08c08ff",
X"b4050883",
X"c08c08ff",
X"bc05088a",
X"052383c0",
X"8c08ffbc",
X"050880d2",
X"053383c0",
X"8c08ffbc",
X"050880d4",
X"05080583",
X"c08c08ff",
X"bc050880",
X"d4050c83",
X"c08c08d8",
X"05080d83",
X"c08c08d0",
X"05088180",
X"0a298180",
X"0a057098",
X"2c83c08c",
X"08c80508",
X"81053383",
X"c08c08ff",
X"a8050c51",
X"83c08c08",
X"d0050c83",
X"c08c08ff",
X"a8050883",
X"c08c08d0",
X"050824ea",
X"a438800b",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"dc05080d",
X"83c08c08",
X"ffa80508",
X"83c0800c",
X"9c3d0d83",
X"c08c0c04",
X"f33d0d02",
X"bf053302",
X"840580c3",
X"053383ca",
X"fc335a5b",
X"5979802e",
X"8d387878",
X"06577680",
X"2e8e3881",
X"89397878",
X"06577680",
X"2e80ff38",
X"83cafc33",
X"707a0758",
X"58798838",
X"78097079",
X"06515776",
X"83cafc34",
X"92973f83",
X"c080085e",
X"805c8f5d",
X"7d1c8711",
X"33585876",
X"802e80c1",
X"38770881",
X"db8c2e09",
X"8106b638",
X"805b815a",
X"7d1c701c",
X"9a113359",
X"59597682",
X"2e098106",
X"943883ca",
X"fc568155",
X"80547653",
X"97183352",
X"7851c98a",
X"3fff1a80",
X"d81c5c5a",
X"798025d0",
X"38ff1d81",
X"c41d5d5d",
X"7c8025ff",
X"a7388f3d",
X"0d04e93d",
X"0d696c02",
X"880580ea",
X"05225c5a",
X"5b807071",
X"415e58ff",
X"78797a7b",
X"7c7d464c",
X"4a45405d",
X"4362993d",
X"34620284",
X"0580dd05",
X"34777922",
X"80ffff06",
X"54457279",
X"2379782e",
X"8887387a",
X"7081055c",
X"3370842a",
X"718c0670",
X"822a5a56",
X"568306ff",
X"1b7083ff",
X"ff065c54",
X"56805475",
X"742e9138",
X"7a708105",
X"5c33ff1b",
X"7083ffff",
X"065c5454",
X"8176279b",
X"387381ff",
X"067b7081",
X"055d3355",
X"74828029",
X"05ff1b70",
X"83ffff06",
X"5c545482",
X"7627aa38",
X"7383ffff",
X"067b7081",
X"055d3370",
X"902b7207",
X"7d708105",
X"5f337098",
X"2b7207fe",
X"1f7083ff",
X"ff064052",
X"52525254",
X"547e802e",
X"80c43876",
X"86f73874",
X"8a2e0981",
X"06943881",
X"1f7081ff",
X"06811e70",
X"81ff065f",
X"52405386",
X"dc39748c",
X"2e098106",
X"86d338ff",
X"1f7081ff",
X"06ff1e70",
X"81ff065f",
X"5240537b",
X"632586bd",
X"38ff4386",
X"b8397681",
X"2e83bb38",
X"76812489",
X"3876802e",
X"8d3886a5",
X"3976822e",
X"84a63886",
X"9c39f815",
X"53728426",
X"84953872",
X"842981de",
X"88055372",
X"08046480",
X"2e80cd38",
X"78228380",
X"80065372",
X"8380802e",
X"098106bc",
X"38805675",
X"6427a438",
X"751e7083",
X"ffff0677",
X"101b9011",
X"72832a58",
X"51575153",
X"73753472",
X"87068171",
X"2b515372",
X"81163481",
X"167081ff",
X"06575397",
X"7627cc38",
X"7f840740",
X"800b993d",
X"43566116",
X"70337098",
X"2b70982c",
X"51515153",
X"80732480",
X"fb386073",
X"291e7083",
X"ffff067a",
X"22838080",
X"06525853",
X"72838080",
X"2e098106",
X"80de3860",
X"88327030",
X"70720780",
X"25639032",
X"70307072",
X"07802573",
X"07535458",
X"51555373",
X"802ebd38",
X"76870653",
X"72b63875",
X"84297610",
X"05791184",
X"1179832a",
X"57575153",
X"73753460",
X"81163465",
X"86142366",
X"88142375",
X"87387f81",
X"07408d39",
X"75812e09",
X"81068538",
X"7f820740",
X"81167081",
X"ff065753",
X"817627fe",
X"e5386361",
X"291e7083",
X"ffff065f",
X"53807046",
X"42ff0284",
X"0580dd05",
X"34ff0b99",
X"3d3483f5",
X"39811c70",
X"81ff065d",
X"53804273",
X"812e0981",
X"068e3877",
X"81800a29",
X"81800a05",
X"5880d339",
X"73802e89",
X"3873822e",
X"0981068d",
X"387c8180",
X"0a298180",
X"0a055da4",
X"39815f83",
X"b839ff1c",
X"7081ff06",
X"5d537b63",
X"258338ff",
X"437c802e",
X"92387c81",
X"800a2981",
X"ff0a055d",
X"7c982c5d",
X"83933977",
X"802e9238",
X"7781800a",
X"2981ff0a",
X"05587798",
X"2c5882fd",
X"39775383",
X"9e397489",
X"2680f438",
X"74842981",
X"de9c0553",
X"72080473",
X"872e82e1",
X"3873852e",
X"82db3873",
X"882e82d5",
X"38738c2e",
X"82cf3873",
X"892e0981",
X"06863881",
X"4582c239",
X"73812e09",
X"810682b9",
X"38628025",
X"82b3387b",
X"982b7098",
X"2c514382",
X"a8397383",
X"ffff0646",
X"829f3973",
X"83ffff06",
X"47829639",
X"7381ff06",
X"41828e39",
X"73811a34",
X"82873973",
X"81ff0644",
X"81ff397e",
X"5382a039",
X"74812e81",
X"e3387481",
X"24893874",
X"802e8d38",
X"81e73974",
X"822e81d8",
X"3881de39",
X"74567b83",
X"38815674",
X"5373862e",
X"09810697",
X"38758106",
X"5372802e",
X"8e387822",
X"82ffff06",
X"fe808007",
X"53b6397b",
X"83388153",
X"73822e09",
X"81069738",
X"72810653",
X"72802e8e",
X"38782281",
X"ffff0681",
X"80800753",
X"93397b96",
X"38fc1453",
X"7281268e",
X"387822ff",
X"80800753",
X"72792380",
X"e5398055",
X"73812e09",
X"81068338",
X"73557753",
X"77802e89",
X"38748106",
X"537280ca",
X"3872d015",
X"54557281",
X"26833881",
X"5577802e",
X"b9387481",
X"06537280",
X"2eb03878",
X"22838080",
X"06537283",
X"80802e09",
X"81069f38",
X"73b02e09",
X"81068738",
X"61993d34",
X"913973b1",
X"2e098106",
X"89386102",
X"840580dd",
X"05346181",
X"05538c39",
X"61743181",
X"05538439",
X"61145372",
X"83ffff06",
X"4279f7fb",
X"387d832a",
X"5372821a",
X"34782283",
X"80800653",
X"72838080",
X"2e098106",
X"88388153",
X"7f872e83",
X"38805372",
X"83c0800c",
X"993d0d04",
X"fd3d0d75",
X"83113382",
X"12337198",
X"2b71902b",
X"07811433",
X"70882b72",
X"07753371",
X"0783c080",
X"0c525354",
X"56545285",
X"3d0d04f6",
X"3d0d02b7",
X"05330284",
X"05bb0533",
X"028805bf",
X"05335b5b",
X"5b805880",
X"5778882b",
X"7a075680",
X"557a5481",
X"53a3527c",
X"5192cc3f",
X"83c08008",
X"81ff0683",
X"c0800c8c",
X"3d0d04f6",
X"3d0d02b7",
X"05330284",
X"05bb0533",
X"028805bf",
X"05335b5b",
X"5b805880",
X"5778882b",
X"7a075680",
X"557a5483",
X"53a3527c",
X"5192903f",
X"83c08008",
X"81ff0683",
X"c0800c8c",
X"3d0d04f7",
X"3d0d02b3",
X"05330284",
X"05b60522",
X"605a5856",
X"80558054",
X"805381a3",
X"527b5191",
X"e23f83c0",
X"800881ff",
X"0683c080",
X"0c8b3d0d",
X"04ee3d0d",
X"6490115c",
X"5c807b34",
X"800b841c",
X"0c800b88",
X"1c34810b",
X"891c3488",
X"0b8a1c34",
X"800b8b1c",
X"34881b08",
X"c1068107",
X"881c0c8f",
X"3d70545d",
X"88527b51",
X"9c923f83",
X"c0800881",
X"ff06705b",
X"597881a9",
X"38903d33",
X"5e81db5a",
X"7d892e09",
X"81068199",
X"387c5392",
X"527b519b",
X"eb3f83c0",
X"800881ff",
X"06705b59",
X"78818238",
X"7c588857",
X"7856a955",
X"78548653",
X"81a0527b",
X"5190d03f",
X"83c08008",
X"81ff0670",
X"5b597880",
X"e03802ba",
X"05337b34",
X"7c547853",
X"7d527b51",
X"9bd33f83",
X"c0800881",
X"ff06705b",
X"597880c1",
X"3802bd05",
X"33527b51",
X"9beb3f83",
X"c0800881",
X"ff06705b",
X"5978aa38",
X"817b335a",
X"5a797926",
X"99388054",
X"79538852",
X"7b51fdbb",
X"3f811a70",
X"81ff067c",
X"33525b59",
X"e439810b",
X"881c3480",
X"5a7983c0",
X"800c943d",
X"0d04800b",
X"83c0800c",
X"04f93d0d",
X"79028405",
X"ab05338e",
X"3d705458",
X"5858ffbb",
X"f53f8a3d",
X"8a0551ff",
X"bbec3f75",
X"51fc8d3f",
X"83c08008",
X"8486812e",
X"be3883c0",
X"80088486",
X"81269938",
X"83c08008",
X"8482802e",
X"80e63883",
X"c0800884",
X"82812e9f",
X"3881b439",
X"83c08008",
X"80c08283",
X"2e80f438",
X"83c08008",
X"80c08683",
X"2e80e838",
X"81993983",
X"c09c3355",
X"80567476",
X"2e098106",
X"818b3874",
X"54765391",
X"527751fb",
X"d63f7454",
X"76539052",
X"7751fbcb",
X"3f745476",
X"53845277",
X"51fbfc3f",
X"810b83c0",
X"9c3481b1",
X"5680de39",
X"80547653",
X"91527751",
X"fba93f80",
X"54765390",
X"527751fb",
X"9e3f800b",
X"83c09c34",
X"76528718",
X"33519796",
X"3fb53980",
X"54765394",
X"527751fb",
X"823f8054",
X"76539052",
X"7751faf7",
X"3f7551ff",
X"baa03f83",
X"c0800889",
X"2a810653",
X"76528718",
X"335190cd",
X"3f800b83",
X"c09c3480",
X"567583c0",
X"800c893d",
X"0d04f23d",
X"0d609011",
X"5a58800b",
X"881a3371",
X"59565674",
X"762e82a5",
X"3882ac3f",
X"84190883",
X"c0800826",
X"82953878",
X"335a810b",
X"8e3d2390",
X"3df81155",
X"f4055399",
X"18527751",
X"8ae53f83",
X"c0800881",
X"ff067057",
X"5574772e",
X"09810681",
X"d9388639",
X"745681d2",
X"39815682",
X"578e3d33",
X"77065574",
X"802ebb38",
X"800b8d3d",
X"34903df0",
X"05548453",
X"75527751",
X"facd3f83",
X"c0800881",
X"ff065574",
X"9d387b53",
X"75527751",
X"fce73f83",
X"c0800881",
X"ff065574",
X"81b12e81",
X"8b3874ff",
X"b3387610",
X"81fc0681",
X"177081ff",
X"06585657",
X"877627ff",
X"a8388156",
X"757a2680",
X"eb38800b",
X"8d3d348c",
X"3d705557",
X"84537552",
X"7751f9f7",
X"3f83c080",
X"0881ff06",
X"557480c1",
X"387651ff",
X"b89c3f83",
X"c0800882",
X"87065574",
X"82812e09",
X"8106aa38",
X"02ae0533",
X"81075574",
X"028405ae",
X"05347b53",
X"75527751",
X"fbeb3f83",
X"c0800881",
X"ff065574",
X"81b12e90",
X"3874feb8",
X"38811670",
X"81ff0657",
X"55ff9139",
X"80567581",
X"ff065697",
X"3f83c080",
X"088fd005",
X"841a0c75",
X"577683c0",
X"800c903d",
X"0d040490",
X"80a00883",
X"c0800c04",
X"ff3d0d73",
X"87e82951",
X"ff8ca43f",
X"833d0d04",
X"0483cb80",
X"0b83c080",
X"0c04fd3d",
X"0d757754",
X"54800b83",
X"cae03472",
X"8a389090",
X"800b8415",
X"0c903972",
X"812e0981",
X"06883890",
X"98800b84",
X"150c8414",
X"0883caf8",
X"0c800b88",
X"150c800b",
X"8c150c83",
X"caf80853",
X"820b8780",
X"14348151",
X"ff9e3f83",
X"caf80853",
X"800b8814",
X"3483caf8",
X"0853810b",
X"87801434",
X"83caf808",
X"53800b8c",
X"143483ca",
X"f8085380",
X"0ba41434",
X"91743480",
X"0b83c0a0",
X"34800b83",
X"c0a43480",
X"0b83c0a8",
X"34805473",
X"81c42983",
X"cb840553",
X"800b8314",
X"34811470",
X"81ff0655",
X"538f7427",
X"e638853d",
X"0d04fe3d",
X"0d747682",
X"113370bf",
X"0681712b",
X"ff055651",
X"51525390",
X"71278338",
X"ff527651",
X"71712383",
X"caf80851",
X"87133390",
X"1234800b",
X"83c0a434",
X"800b83c0",
X"a8348813",
X"338a1433",
X"52527180",
X"2eaa3870",
X"81ff0651",
X"84527083",
X"38705271",
X"83c0a434",
X"8a133370",
X"30708025",
X"842b7088",
X"07515152",
X"537083c0",
X"a8349039",
X"7081ff06",
X"51708338",
X"98527183",
X"c0a83480",
X"0b83c080",
X"0c843d0d",
X"04f13d0d",
X"61656802",
X"8c0580cb",
X"05330290",
X"0580ce05",
X"22029405",
X"80d60522",
X"4240415a",
X"4040fd8b",
X"3f83c080",
X"08a78805",
X"5b807071",
X"5b5b5283",
X"943983ca",
X"f808517d",
X"94123483",
X"c0a43381",
X"07558070",
X"54567f86",
X"2680ea38",
X"7f842981",
X"ded00583",
X"caf80853",
X"51700804",
X"800b8413",
X"34a13977",
X"33703070",
X"80258371",
X"31515152",
X"53708413",
X"348d3981",
X"0b841334",
X"b839830b",
X"84133481",
X"705456ad",
X"39810b84",
X"1334a239",
X"77337030",
X"70802583",
X"71315151",
X"52537084",
X"13348078",
X"33525270",
X"83388152",
X"71783481",
X"53748807",
X"5583c0a8",
X"3383caf8",
X"08525781",
X"0b81d012",
X"3483caf8",
X"0851810b",
X"81901234",
X"7e802eae",
X"3872802e",
X"a9387eff",
X"1e525470",
X"83ffff06",
X"537283ff",
X"ff2e9738",
X"73708105",
X"553383ca",
X"f8085351",
X"7081c013",
X"34ff1351",
X"de3983ca",
X"f808a811",
X"33535176",
X"88123483",
X"caf80851",
X"74713481",
X"ff529139",
X"83caf808",
X"a0113370",
X"81065152",
X"53708f38",
X"fafd3f7a",
X"83c08008",
X"26e63881",
X"8839810b",
X"a0143483",
X"caf808a8",
X"113380ff",
X"06707807",
X"52535170",
X"802e80ed",
X"3871862a",
X"70810651",
X"5170802e",
X"91388078",
X"33525370",
X"83388153",
X"72783480",
X"e0397184",
X"2a708106",
X"51517080",
X"2e9b3881",
X"197083ff",
X"ff067d30",
X"709f2a51",
X"525a5178",
X"7c2e0981",
X"06af38a4",
X"3971832a",
X"70810651",
X"5170802e",
X"9338811a",
X"7081ff06",
X"5b517983",
X"2e098106",
X"90388a39",
X"71a30651",
X"70802e85",
X"38715192",
X"39f9e43f",
X"7a83c080",
X"0826fce2",
X"387181bf",
X"06517083",
X"c0800c91",
X"3d0d04f6",
X"3d0d02b3",
X"05330284",
X"05b70533",
X"028805ba",
X"05225959",
X"59800b8c",
X"3d348c3d",
X"fc055680",
X"55805476",
X"53775278",
X"51fbf23f",
X"83c08008",
X"81ff0683",
X"c0800c8c",
X"3d0d04f3",
X"3d0d7f62",
X"64028c05",
X"80c20522",
X"72228115",
X"33425f41",
X"5e595980",
X"78237d53",
X"78335281",
X"51ffa03f",
X"83c08008",
X"81ff0656",
X"75802e86",
X"38755481",
X"ad3983ca",
X"f808a811",
X"33821b33",
X"70862a70",
X"81067398",
X"2b535157",
X"5c565779",
X"80258338",
X"81567376",
X"2e873881",
X"f0548182",
X"39818c17",
X"337081ff",
X"0679227d",
X"7131902b",
X"70902c70",
X"09709f2c",
X"72067052",
X"52535153",
X"57575475",
X"74248338",
X"75557484",
X"808029fc",
X"80800570",
X"902c5155",
X"74ff2e94",
X"3883caf8",
X"08818011",
X"33515473",
X"7c708105",
X"5e34db39",
X"77227605",
X"54737823",
X"7909709f",
X"2a708106",
X"821c3381",
X"bf067186",
X"2b075151",
X"51547382",
X"1a347c76",
X"268a3877",
X"22547a74",
X"26febb38",
X"80547383",
X"c0800c8f",
X"3d0d04f9",
X"3d0d7a57",
X"800b893d",
X"23893dfc",
X"05537652",
X"7951f8da",
X"3f83c080",
X"0881ff06",
X"70575574",
X"96387c54",
X"7b53883d",
X"22527651",
X"fde53f83",
X"c0800881",
X"ff065675",
X"83c0800c",
X"893d0d04",
X"f03d0d62",
X"66028805",
X"80ce0522",
X"415d5e80",
X"02840580",
X"d205227f",
X"810533ff",
X"115a5d5a",
X"5d81da58",
X"76bf2680",
X"e9387880",
X"2e80e138",
X"7a58787b",
X"27833878",
X"58821e33",
X"70872a58",
X"5a76923d",
X"34923dfc",
X"05567755",
X"7b547e53",
X"7d335282",
X"51f8de3f",
X"83c08008",
X"81ff065d",
X"800b923d",
X"33585a76",
X"802e8338",
X"815a821e",
X"3380ff06",
X"7a872b07",
X"5776821f",
X"347c9138",
X"78783170",
X"83ffff06",
X"791e5e5a",
X"57ff9b39",
X"7c587783",
X"c0800c92",
X"3d0d04f8",
X"3d0d7b02",
X"8405b205",
X"22585880",
X"0b8a3d23",
X"8a3dfc05",
X"5377527a",
X"51f6f73f",
X"83c08008",
X"81ff0670",
X"57557496",
X"387d5476",
X"53893d22",
X"527751fe",
X"af3f83c0",
X"800881ff",
X"06567583",
X"c0800c8a",
X"3d0d04ec",
X"3d0d666e",
X"02880580",
X"df053302",
X"8c0580e3",
X"05330290",
X"0580e705",
X"33029405",
X"80eb0533",
X"02980580",
X"ee052241",
X"43415f5c",
X"40570280",
X"f2052296",
X"3d23963d",
X"f0055384",
X"17705377",
X"5259f686",
X"3f83c080",
X"0881ff06",
X"587781e5",
X"38777a81",
X"80065840",
X"80772583",
X"38814079",
X"943d347b",
X"02840580",
X"c905347c",
X"02840580",
X"ca05347d",
X"02840580",
X"cb05347a",
X"953d347a",
X"882a5776",
X"02840580",
X"cd053495",
X"3d225776",
X"02840580",
X"ce053476",
X"882a5776",
X"02840580",
X"cf053477",
X"923d3496",
X"3dec1157",
X"578855f4",
X"1754923d",
X"22537752",
X"7751f695",
X"3f83c080",
X"0881ff06",
X"587780ed",
X"387e802e",
X"80cb3892",
X"3d227908",
X"58587f80",
X"2e9c3876",
X"81808007",
X"790c7e54",
X"963dfc05",
X"537783ff",
X"ff065278",
X"51f9fc3f",
X"99397682",
X"80800779",
X"0c7e5495",
X"3d225377",
X"83ffff06",
X"527851fc",
X"8f3f83c0",
X"800881ff",
X"0658779d",
X"38923d22",
X"5380527f",
X"30708025",
X"84713153",
X"5157f987",
X"3f83c080",
X"0881ff06",
X"587783c0",
X"800c963d",
X"0d04f63d",
X"0d7c0284",
X"05b70533",
X"5b5b8058",
X"80578056",
X"80557954",
X"85538052",
X"7a51fda3",
X"3f83c080",
X"0881ff06",
X"59788538",
X"79871c34",
X"7883c080",
X"0c8c3d0d",
X"04f93d0d",
X"02a70533",
X"028405ab",
X"05330288",
X"05af0533",
X"58595780",
X"0b83cb87",
X"33545472",
X"742e9f38",
X"81147081",
X"ff065553",
X"738f2681",
X"b6387381",
X"c42983cb",
X"84058311",
X"33515372",
X"e3387381",
X"c42983cb",
X"80055580",
X"0b871634",
X"76881634",
X"758a1634",
X"77891634",
X"80750c83",
X"caf8088c",
X"160c800b",
X"84163488",
X"0b851634",
X"800b8616",
X"34841508",
X"ffa1ff06",
X"a0800784",
X"160c8114",
X"7081ff06",
X"53537451",
X"febc3f83",
X"c0800881",
X"ff067055",
X"537280cd",
X"388a3973",
X"08750c72",
X"5480c239",
X"7281e5b0",
X"555681e5",
X"b008802e",
X"b2387584",
X"29147008",
X"76537008",
X"51545472",
X"2d83c080",
X"0881ff06",
X"5372802e",
X"ce388116",
X"7081ff06",
X"81e5b071",
X"84291153",
X"56575372",
X"08d03880",
X"547383c0",
X"800c893d",
X"0d04f93d",
X"0d795780",
X"0b841808",
X"83caf80c",
X"58f0883f",
X"88170883",
X"c0800827",
X"83ed38ef",
X"fa3f83c0",
X"80088105",
X"88180c83",
X"caf808b8",
X"11337081",
X"ff065151",
X"5473812e",
X"a4387381",
X"24883873",
X"782e8a38",
X"b8397382",
X"2e9538b1",
X"39763381",
X"f0065473",
X"902ea638",
X"917734a1",
X"39735876",
X"3381f006",
X"5473902e",
X"09810691",
X"38efa83f",
X"83c08008",
X"81c8058c",
X"180ca077",
X"34805675",
X"81c42983",
X"cb871133",
X"55557380",
X"2eaa3883",
X"cb801570",
X"08565474",
X"802e9d38",
X"88150880",
X"2e96388c",
X"140883ca",
X"f8082e09",
X"81068938",
X"73518815",
X"0854732d",
X"81167081",
X"ff065754",
X"8f7627ff",
X"ba387633",
X"5473b02e",
X"81993873",
X"b0248f38",
X"73912eab",
X"3873a02e",
X"80f53882",
X"a6397380",
X"d02e81e4",
X"387380d0",
X"248b3873",
X"80c02e81",
X"9938828f",
X"39738180",
X"2e81fb38",
X"82853980",
X"567581c4",
X"2983cb84",
X"11831133",
X"56595573",
X"802ea838",
X"83cb8015",
X"70085654",
X"74802e9b",
X"388c1408",
X"83caf808",
X"2e098106",
X"8e387351",
X"84150854",
X"732d800b",
X"83193481",
X"167081ff",
X"0657548f",
X"7627ffb9",
X"38927734",
X"81b539ed",
X"c23f8c17",
X"0883c080",
X"082781a7",
X"38b07734",
X"81a13983",
X"caf80854",
X"800b8c15",
X"3483caf8",
X"0854840b",
X"88153480",
X"c07734ed",
X"963f83c0",
X"8008b205",
X"8c180c80",
X"fa39ed87",
X"3f8c1708",
X"83c08008",
X"2780ec38",
X"83caf808",
X"54810b8c",
X"153483ca",
X"f8085480",
X"0b881534",
X"83caf808",
X"54880ba0",
X"1534ecdb",
X"3f83c080",
X"0894058c",
X"180c80d0",
X"7734bc39",
X"83caf808",
X"a0113370",
X"832a7081",
X"06515155",
X"5573802e",
X"a638880b",
X"a01634ec",
X"ae3f8c17",
X"0883c080",
X"08279438",
X"ff807734",
X"8e397753",
X"80528051",
X"fa8b3fff",
X"90773483",
X"caf808a0",
X"11337083",
X"2a708106",
X"51515555",
X"73802e86",
X"38880ba0",
X"1634893d",
X"0d04f43d",
X"0d02bb05",
X"33028405",
X"bf05335d",
X"5d800b83",
X"cb840b83",
X"cb800b8c",
X"11727188",
X"14755c5a",
X"5b5f5c59",
X"5b588315",
X"33537280",
X"2e818838",
X"7333537c",
X"732e0981",
X"0680fc38",
X"81143353",
X"7b732e09",
X"810680ef",
X"38750883",
X"caf8082e",
X"09810680",
X"e2388056",
X"7581c429",
X"83cb8811",
X"7033831e",
X"335b5755",
X"5374782e",
X"09810697",
X"3883cb8c",
X"13087908",
X"2e098106",
X"8a388114",
X"33527451",
X"fef83f81",
X"167081ff",
X"0657538f",
X"7627c538",
X"80770854",
X"5472742e",
X"91387651",
X"84130853",
X"722d83c0",
X"800881ff",
X"0654800b",
X"831b3473",
X"53a93981",
X"1881c416",
X"81c41681",
X"c41981c4",
X"1f81c41e",
X"81c41d60",
X"81c40541",
X"5d5e5f59",
X"5656588f",
X"7825feca",
X"38805372",
X"83c0800c",
X"8e3d0d04",
X"f83d0d02",
X"ae05227d",
X"59578056",
X"81558054",
X"86538180",
X"527a51f4",
X"ee3f83c0",
X"800881ff",
X"0683c080",
X"0c8a3d0d",
X"04f73d0d",
X"02b20522",
X"028405b7",
X"0533605a",
X"5b578056",
X"82557954",
X"86538180",
X"527b51f4",
X"be3f83c0",
X"800881ff",
X"0683c080",
X"0c8b3d0d",
X"04f83d0d",
X"02af0533",
X"59805880",
X"57805680",
X"55785489",
X"5380527a",
X"51f4943f",
X"83c08008",
X"81ff0683",
X"c0800c8a",
X"3d0d0400",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002bd6",
X"00002c17",
X"00002c39",
X"00002c5b",
X"00002c81",
X"00002c81",
X"00002c81",
X"00002c81",
X"00002cf2",
X"00002d47",
X"00002d47",
X"00002d87",
X"00004332",
X"00004bc0",
X"00004c89",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3f00",
X"0c0c4000",
X"0a0a4100",
X"0b0b4100",
X"07074100",
X"0a0b4300",
X"080b4200",
X"04044500",
X"05054400",
X"0e0f2900",
X"06060004",
X"08080004",
X"09090004",
X"080f4300",
X"090f4200",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"000059f6",
X"00005cfd",
X"00005b09",
X"00005cfd",
X"00005b46",
X"00005b97",
X"00005bd6",
X"00005bdf",
X"00005cfd",
X"00005cfd",
X"00005cfd",
X"00005cfd",
X"00005be8",
X"00005bf0",
X"00005bf7",
X"00005dfd",
X"00005ef6",
X"0000600a",
X"00006300",
X"0000631b",
X"00006307",
X"0000631b",
X"00006322",
X"0000632d",
X"00006334",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"43505520",
X"54757262",
X"6f3a2564",
X"78000000",
X"44726976",
X"65205475",
X"72626f3a",
X"25730000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"4c6f6164",
X"206d656d",
X"6f727900",
X"53617665",
X"206d656d",
X"6f727920",
X"28666f72",
X"20646562",
X"75676769",
X"6e672900",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"66726565",
X"7a65722e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"4d454d00",
X"5374616e",
X"64617264",
X"00000000",
X"46617374",
X"28362900",
X"46617374",
X"28352900",
X"46617374",
X"28342900",
X"46617374",
X"28332900",
X"46617374",
X"28322900",
X"46617374",
X"28312900",
X"46617374",
X"28302900",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00006fac",
X"00006fb0",
X"00006fb8",
X"00006fc4",
X"00006fd0",
X"00006fdc",
X"00006fe8",
X"00006fec",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00000028",
X"00000006",
X"00000005",
X"00000004",
X"00000003",
X"00000002",
X"00000001",
X"00000000",
X"000070b8",
X"000070c4",
X"000070cc",
X"000070d4",
X"000070dc",
X"000070e4",
X"000070ec",
X"000070f4",
X"00006f44",
X"00006d8c",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"69383030",
X"00000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
