
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f8",
X"c4738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80fb",
X"980c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f2",
X"f42d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580f188",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"96ea0480",
X"3d0d80fc",
X"dc087008",
X"810683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d80fc",
X"dc087008",
X"70fe0676",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80fcdc08",
X"70087081",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80fcdc08",
X"700870fd",
X"06761007",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"fcdc0870",
X"0870822c",
X"bf0683e0",
X"800c5151",
X"823d0d04",
X"ff3d0d80",
X"fcdc0870",
X"0870fe83",
X"0676822b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80fcdc08",
X"70087088",
X"2c870683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80fcdc08",
X"700870f1",
X"ff067688",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d80fcdc",
X"08700870",
X"8b2cbf06",
X"83e0800c",
X"5151823d",
X"0d04ff3d",
X"0d80fcdc",
X"08700870",
X"f88fff06",
X"768b2b07",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"fcec0870",
X"0870882c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fcec0870",
X"0870892c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fcec0870",
X"08708a2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fcec0870",
X"08708b2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"fd3d0d75",
X"81e62987",
X"2a80fccc",
X"0854730c",
X"853d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d848080",
X"53805288",
X"800a51ff",
X"b33f8180",
X"80538052",
X"82800a51",
X"c63f843d",
X"0d04803d",
X"0d8151fc",
X"ce3f7280",
X"2e8338d2",
X"3f8151fc",
X"f03f8051",
X"fceb3f80",
X"51fcb83f",
X"823d0d04",
X"fd3d0d75",
X"52805480",
X"ff722588",
X"38810bff",
X"80135354",
X"ffbf1251",
X"70992686",
X"38e01252",
X"9e39ff9f",
X"12519971",
X"279538d0",
X"12e01370",
X"54545189",
X"71278838",
X"8f732783",
X"38805273",
X"802e8538",
X"81801252",
X"7181ff06",
X"83e0800c",
X"853d0d04",
X"803d0d86",
X"b8c05180",
X"71708105",
X"53347086",
X"c0c02e09",
X"8106f038",
X"823d0d04",
X"fe3d0d02",
X"97053351",
X"ff863f83",
X"e0800881",
X"ff0683e0",
X"9c085452",
X"8073249b",
X"3883e0b8",
X"08137283",
X"e0bc0807",
X"53537173",
X"3483e09c",
X"08810583",
X"e09c0c84",
X"3d0d04fa",
X"3d0d8280",
X"0a1b5580",
X"57883dfc",
X"05547953",
X"74527851",
X"b4f93f88",
X"3d0d04fe",
X"3d0d83e0",
X"b0085274",
X"51bbdb3f",
X"83e08008",
X"8c387653",
X"755283e0",
X"b00851c7",
X"3f843d0d",
X"04fe3d0d",
X"83e0b008",
X"53755274",
X"51b69b3f",
X"83e08008",
X"8d387753",
X"765283e0",
X"b00851ff",
X"a23f843d",
X"0d04fe3d",
X"0d83e0b4",
X"0851b58f",
X"3f83e080",
X"08818080",
X"2e098106",
X"883883c1",
X"8080539b",
X"3983e0b4",
X"0851b4f3",
X"3f83e080",
X"0880d080",
X"2e098106",
X"933883c1",
X"b0805383",
X"e0800852",
X"83e0b408",
X"51fed83f",
X"843d0d04",
X"803d0dfa",
X"cc3f83e0",
X"80088429",
X"80fba005",
X"700883e0",
X"800c5182",
X"3d0d04ee",
X"3d0d8043",
X"80428041",
X"80705a5b",
X"fdd23f80",
X"0b83e09c",
X"0c800b83",
X"e0bc0c0b",
X"0b80f9e0",
X"51afdd3f",
X"81800b83",
X"e0bc0c0b",
X"0b80f9e4",
X"51afcd3f",
X"80d00b83",
X"e09c0c78",
X"30707a07",
X"80257087",
X"2b83e0bc",
X"0c5155f9",
X"b73f83e0",
X"8008520b",
X"0b80f9ec",
X"51afa53f",
X"80f80b83",
X"e09c0c78",
X"81327030",
X"70720780",
X"2570872b",
X"83e0bc0c",
X"515656fe",
X"eb3f83e0",
X"8008520b",
X"0b80f9f8",
X"51aef93f",
X"81a00b83",
X"e09c0c78",
X"82327030",
X"70720780",
X"2570872b",
X"83e0bc0c",
X"515683e0",
X"b4085256",
X"b0943f83",
X"e0800852",
X"0b0b80fa",
X"8051aec8",
X"3f81f00b",
X"83e09c0c",
X"810b83e0",
X"a05b5883",
X"e09c0882",
X"197a3270",
X"30707207",
X"80257087",
X"2b83e0bc",
X"0c51578e",
X"3d7055ff",
X"1b545757",
X"57a4a63f",
X"79708405",
X"5b0851af",
X"c93f7454",
X"83e08008",
X"5377520b",
X"0b80fa88",
X"51adf93f",
X"a81783e0",
X"9c0c8118",
X"5877852e",
X"098106ff",
X"ae388390",
X"0b83e09c",
X"0c788732",
X"70307072",
X"07802570",
X"872b83e0",
X"bc0c5156",
X"0b0b80fa",
X"985256ad",
X"c33f83e0",
X"0b83e09c",
X"0c788832",
X"70307072",
X"07802570",
X"872b83e0",
X"bc0c5156",
X"0b0b80fa",
X"ac5256ad",
X"9f3f868d",
X"a051f990",
X"3f805291",
X"3d705255",
X"8ba53f83",
X"5274518b",
X"9e3f6119",
X"59788025",
X"85388059",
X"90398879",
X"25853888",
X"59873978",
X"882682ae",
X"3878822b",
X"5580f8d4",
X"150804f6",
X"e33f83e0",
X"80086157",
X"5575812e",
X"09810689",
X"3883e080",
X"08105590",
X"3975ff2e",
X"09810688",
X"3883e080",
X"08812c55",
X"90752585",
X"38905588",
X"39748024",
X"83388155",
X"7451f6c0",
X"3f81e339",
X"f6d33f83",
X"e0800861",
X"05557480",
X"25853880",
X"55883987",
X"75258338",
X"87557451",
X"f6cf3f81",
X"c1396087",
X"3862802e",
X"81b838a0",
X"990b83e0",
X"d00c83e0",
X"b408518c",
X"a93ffafe",
X"3f81a339",
X"60568076",
X"2598389f",
X"b80b83e0",
X"d00c83e0",
X"94157008",
X"52558c8a",
X"3f740852",
X"91397580",
X"25913883",
X"e0941508",
X"51ad853f",
X"8052fd19",
X"51b83962",
X"802e80ea",
X"3883e094",
X"15700883",
X"e0a00872",
X"0c83e0a0",
X"0cfd1a70",
X"53515596",
X"dc3f83e0",
X"80085680",
X"5196d23f",
X"83e08008",
X"52745192",
X"f13f7552",
X"805192ea",
X"3fb43962",
X"802eaf38",
X"a0990b83",
X"e0d00c83",
X"e0b00851",
X"8ba03f83",
X"e0b00851",
X"ac943f9c",
X"800a5380",
X"c0805283",
X"e0800851",
X"f9993f81",
X"558c3962",
X"87387a80",
X"2efac538",
X"80557483",
X"e0800c94",
X"3d0d04fe",
X"3d0df5c0",
X"3f83e080",
X"08802e86",
X"38805180",
X"f639f5c8",
X"3f83e080",
X"0880ea38",
X"f5ee3f83",
X"e0800880",
X"2eaa3881",
X"51f3c03f",
X"839b3f80",
X"0b83e09c",
X"0cf9f43f",
X"83e08008",
X"53ff0b83",
X"e09c0c85",
X"ee3f72bd",
X"387251f3",
X"9e3fbb39",
X"f5a23f83",
X"e0800880",
X"2eb03881",
X"51f38c3f",
X"82e73f9f",
X"b80b83e0",
X"d00c83e0",
X"a0085189",
X"fd3fff0b",
X"83e09c0c",
X"85b93f83",
X"e0a00852",
X"8051919e",
X"3f8151f6",
X"8d3f843d",
X"0d0483e0",
X"8c080283",
X"e08c0cfa",
X"3d0d800b",
X"83e0a00b",
X"83e08c08",
X"fc050c83",
X"e08c08f8",
X"050cadd0",
X"3f83e080",
X"088605fc",
X"0683e08c",
X"08f4050c",
X"0283e08c",
X"08f40508",
X"310d853d",
X"7083e08c",
X"08fc0508",
X"70840583",
X"e08c08fc",
X"050c0c51",
X"aa9a3f83",
X"e08c08f8",
X"05088105",
X"83e08c08",
X"f8050c83",
X"e08c08f8",
X"0508862e",
X"098106ff",
X"ad388688",
X"80805181",
X"aa3fff0b",
X"83e09c0c",
X"800b83e0",
X"bc0c86b8",
X"c00b83e0",
X"b80c8151",
X"f1c93f81",
X"51f1f23f",
X"8051f1ed",
X"3f8151f2",
X"973f8151",
X"f2f43f82",
X"51f2be3f",
X"8e845280",
X"51a7de3f",
X"84808052",
X"86848080",
X"51adb93f",
X"83e08008",
X"80d33893",
X"b53f80fe",
X"a451b1f8",
X"3f83e080",
X"0883e0b4",
X"08540b0b",
X"80fab453",
X"83e08008",
X"5283e08c",
X"08f4050c",
X"accc3f83",
X"e0800884",
X"38f6bf3f",
X"9c800a54",
X"80c08053",
X"0b0b80fa",
X"c05283e0",
X"8c08f405",
X"0851f681",
X"3f8151f3",
X"f13f9d8d",
X"3f8151f3",
X"e93ffccf",
X"3ffc3971",
X"83e0c40c",
X"8880800b",
X"83e0c00c",
X"8480800b",
X"83e0c80c",
X"04f03d0d",
X"80fbd408",
X"54733383",
X"e0cc3483",
X"a0805683",
X"e0c40816",
X"83e0c008",
X"17565474",
X"33743483",
X"e0c80816",
X"54807434",
X"81165675",
X"83a0a02e",
X"098106db",
X"3883a480",
X"5683e0c4",
X"081683e0",
X"c0081756",
X"54743374",
X"3483e0c8",
X"08165480",
X"74348116",
X"567583a4",
X"a02e0981",
X"06db3883",
X"a8805683",
X"e0c40816",
X"83e0c008",
X"17565474",
X"33743483",
X"e0c80816",
X"54807434",
X"81165675",
X"83a8902e",
X"098106db",
X"3880fbd4",
X"0854ff74",
X"34805683",
X"e0c40816",
X"83e0c808",
X"17555573",
X"33753481",
X"16567583",
X"a0802e09",
X"8106e438",
X"83b08056",
X"83e0c408",
X"1683e0c8",
X"08175555",
X"73337534",
X"81165675",
X"8480802e",
X"098106e4",
X"38f2ed3f",
X"893d58a2",
X"5380f8f8",
X"52775180",
X"dc9f3f80",
X"578c8056",
X"83e0c808",
X"16771955",
X"55733375",
X"34811681",
X"18585676",
X"a22e0981",
X"06e63880",
X"fbf80854",
X"86743480",
X"fbfc0854",
X"80743480",
X"fbf40854",
X"80743480",
X"fbe40854",
X"af743480",
X"fbf00854",
X"bf743480",
X"fbec0854",
X"80743480",
X"fbe80854",
X"9f743480",
X"fbe00854",
X"80743480",
X"fbcc0854",
X"e0743480",
X"fbc40854",
X"76743480",
X"fbc00854",
X"83743480",
X"fbc80854",
X"82743492",
X"3d0d04fe",
X"3d0d8053",
X"83e0c808",
X"1383e0c4",
X"08145252",
X"70337234",
X"81135372",
X"83a0802e",
X"098106e4",
X"3883b080",
X"5383e0c8",
X"081383e0",
X"c4081452",
X"52703372",
X"34811353",
X"72848080",
X"2e098106",
X"e43883a0",
X"805383e0",
X"c8081383",
X"e0c40814",
X"52527033",
X"72348113",
X"537283a0",
X"a02e0981",
X"06e43883",
X"a4805383",
X"e0c80813",
X"83e0c408",
X"14525270",
X"33723481",
X"13537283",
X"a4a02e09",
X"8106e438",
X"83a88053",
X"83e0c808",
X"1383e0c4",
X"08145252",
X"70337234",
X"81135372",
X"83a8902e",
X"098106e4",
X"3880fbd4",
X"085183e0",
X"cc337134",
X"843d0d04",
X"fd3d0d75",
X"5480740c",
X"800b8415",
X"0c800b88",
X"150c80fb",
X"d8087033",
X"7081ff06",
X"70812a81",
X"32718132",
X"71810671",
X"81063184",
X"1a0c5656",
X"70832a81",
X"3271822a",
X"81327181",
X"06718106",
X"31790c52",
X"55515151",
X"80fbd008",
X"70337009",
X"81068817",
X"0c515185",
X"3d0d04fe",
X"3d0d7476",
X"54527151",
X"ff9a3f72",
X"812ea238",
X"8173268d",
X"3872822e",
X"ab387283",
X"2e9f38e6",
X"397108e2",
X"38841208",
X"dd388812",
X"08d838a0",
X"39881208",
X"812e0981",
X"06cc3894",
X"39881208",
X"812e8d38",
X"71088938",
X"84120880",
X"2effb738",
X"843d0d04",
X"fc3d0d76",
X"70525580",
X"c6f63f83",
X"e0800815",
X"ff055473",
X"752e8e38",
X"73335372",
X"ae2e8638",
X"ff1454ef",
X"39775281",
X"145180c6",
X"8d3f83e0",
X"80083070",
X"83e08008",
X"07802583",
X"e0800c53",
X"863d0d04",
X"fc3d0d76",
X"705255ab",
X"e13f83e0",
X"80085481",
X"5383e080",
X"0880c138",
X"7451aba4",
X"3f83e080",
X"0880fadc",
X"5383e080",
X"085253ff",
X"8f3f83e0",
X"8008a138",
X"80fae052",
X"7251ff80",
X"3f83e080",
X"08923880",
X"fae45272",
X"51fef13f",
X"83e08008",
X"802e8338",
X"81547353",
X"7283e080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"ab803f81",
X"5383e080",
X"08973873",
X"51aac93f",
X"80fae852",
X"83e08008",
X"51feb93f",
X"83e08008",
X"537283e0",
X"800c853d",
X"0d04e03d",
X"0da33d08",
X"70525ea0",
X"f13f83e0",
X"80083394",
X"3d565473",
X"943880fe",
X"bc527451",
X"84b3397d",
X"527851a3",
X"f33f84be",
X"397d51a0",
X"d93f83e0",
X"80085274",
X"51a0893f",
X"83e0d008",
X"52933d70",
X"525da6e3",
X"3f83e080",
X"0859800b",
X"83e08008",
X"555b83e0",
X"80087b2e",
X"9438811b",
X"74525ba9",
X"e43f83e0",
X"80085483",
X"e08008ee",
X"38805aff",
X"7a437a42",
X"7a415f79",
X"09709f2c",
X"7b065b54",
X"7a7a2484",
X"38ff1b5a",
X"f61a7009",
X"709f2c72",
X"067bff12",
X"5a5a5255",
X"55807525",
X"95387651",
X"a9a33f83",
X"e0800876",
X"ff185855",
X"57738024",
X"ed38747f",
X"2e8638eb",
X"e33f745f",
X"78ff1b70",
X"585d5880",
X"7a259538",
X"7751a8f9",
X"3f83e080",
X"0876ff18",
X"58555873",
X"8024ed38",
X"800b83e0",
X"9c0c800b",
X"83e0bc0c",
X"80faec51",
X"9dce3f81",
X"800b83e0",
X"bc0c80fa",
X"f4519dc0",
X"3fa80b83",
X"e09c0c76",
X"802e80e4",
X"3883e09c",
X"08777932",
X"70307072",
X"07802570",
X"872b83e0",
X"bc0c5156",
X"78535656",
X"a8b03f83",
X"e0800880",
X"2e883880",
X"fafc519d",
X"873f7651",
X"a7f23f83",
X"e0800852",
X"80fa9451",
X"9cf63f76",
X"51a7fa3f",
X"83e08008",
X"83e09c08",
X"55577574",
X"258638a8",
X"1656f739",
X"7583e09c",
X"0c86f076",
X"24ff9838",
X"87980b83",
X"e09c0c77",
X"802eb138",
X"7751a7b0",
X"3f83e080",
X"08785255",
X"a7d03f80",
X"fb845483",
X"e080088d",
X"38873980",
X"7634fda0",
X"3980fb80",
X"54745373",
X"5280fad0",
X"519c953f",
X"805480fb",
X"8c519c8c",
X"3f811454",
X"73a82e09",
X"8106ef38",
X"868da051",
X"e7f23f80",
X"52903d70",
X"5254fa87",
X"3f835273",
X"51fa803f",
X"61802e80",
X"ff387b54",
X"73ff2e96",
X"3878802e",
X"81803878",
X"51a6da3f",
X"83e08008",
X"ff155559",
X"e7397880",
X"2e80eb38",
X"7851a6d6",
X"3f83e080",
X"08802efc",
X"96387851",
X"a69e3f83",
X"e0800852",
X"80fad851",
X"bfcb3f83",
X"e08008a5",
X"387c5180",
X"c1823f83",
X"e0800855",
X"74ff1656",
X"54807425",
X"fc823874",
X"1d703355",
X"5673af2e",
X"fed138e8",
X"397851a5",
X"dd3f83e0",
X"8008527c",
X"5180c0b8",
X"3ffbe139",
X"7f882960",
X"10057a05",
X"61055afc",
X"9239a23d",
X"0d04803d",
X"0d81ff51",
X"800b83e0",
X"dc1234ff",
X"115170f4",
X"38823d0d",
X"04ff3d0d",
X"73703353",
X"51811133",
X"71347181",
X"1234833d",
X"0d04fb3d",
X"0d777956",
X"56807071",
X"55555271",
X"7525ac38",
X"72167033",
X"70147081",
X"ff065551",
X"51517174",
X"27893881",
X"127081ff",
X"06535171",
X"81147083",
X"ffff0655",
X"52547473",
X"24d63871",
X"83e0800c",
X"873d0d04",
X"fd3d0d75",
X"54948f3f",
X"83e08008",
X"802ef638",
X"83e2f808",
X"86057081",
X"ff065253",
X"91e83f84",
X"39ef903f",
X"93f03f83",
X"e0800881",
X"2ef33892",
X"cb3f83e0",
X"80087434",
X"92c23f83",
X"e0800881",
X"153492b8",
X"3f83e080",
X"08821534",
X"92ae3f83",
X"e0800883",
X"153492a4",
X"3f83e080",
X"08841534",
X"8439eecf",
X"3f93af3f",
X"83e08008",
X"802ef338",
X"733383e0",
X"dc348114",
X"3383e0dd",
X"34821433",
X"83e0de34",
X"83143383",
X"e0df3484",
X"5283e0dc",
X"51fea73f",
X"83e08008",
X"81ff0684",
X"15335553",
X"72742e09",
X"81068c38",
X"92a03f83",
X"e0800880",
X"2e9a3883",
X"e2f808a8",
X"2e098106",
X"8938860b",
X"83e2f80c",
X"8739a80b",
X"83e2f80c",
X"80e451e4",
X"873f853d",
X"0d04f43d",
X"0d7e6059",
X"55805d80",
X"75822b71",
X"83e2fc12",
X"0c83e390",
X"175b5b57",
X"76793477",
X"772e83b1",
X"38765277",
X"519be13f",
X"8e3dfc05",
X"54905383",
X"e2e45277",
X"519b983f",
X"7c567590",
X"2e098106",
X"838f3883",
X"e2e451fd",
X"843f83e2",
X"e651fcfd",
X"3f83e2e8",
X"51fcf63f",
X"7683e2f4",
X"0c775198",
X"e53f80fa",
X"e05283e0",
X"800851f6",
X"873f83e0",
X"8008812e",
X"09810680",
X"d3387683",
X"e38c0c82",
X"0b83e2e4",
X"34ff960b",
X"83e2e534",
X"77519bab",
X"3f83e080",
X"085583e0",
X"80087725",
X"883883e0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83e2e634",
X"7483e2e7",
X"347683e2",
X"e834ff80",
X"0b83e2e9",
X"34818f39",
X"83e2e433",
X"83e2e533",
X"71882b07",
X"565b7483",
X"ffff2e09",
X"810680e7",
X"38fe800b",
X"83e38c0c",
X"810b83e2",
X"f40cff0b",
X"83e2e434",
X"ff0b83e2",
X"e5347751",
X"9ab93f83",
X"e0800883",
X"e3940c83",
X"e0800855",
X"83e08008",
X"80258838",
X"83e08008",
X"8f055574",
X"842c7083",
X"ffff0670",
X"882a5851",
X"557583e2",
X"e6347483",
X"e2e73476",
X"83e2e834",
X"ff800b83",
X"e2e93481",
X"0b83e2f3",
X"34a43974",
X"85962e09",
X"810680fd",
X"387583e3",
X"8c0c7751",
X"99ee3f83",
X"e2f33383",
X"e0800807",
X"557483e2",
X"f33483e2",
X"f3338106",
X"5574802e",
X"83388457",
X"83e2e833",
X"83e2e933",
X"71882b07",
X"565c7481",
X"802e0981",
X"06a13883",
X"e2e63383",
X"e2e73371",
X"882b0756",
X"5bad8075",
X"27873876",
X"8207579c",
X"39768107",
X"57963974",
X"82802e09",
X"81068738",
X"76830757",
X"87397481",
X"ff268a38",
X"7783e2fc",
X"1b0c7679",
X"348e3d0d",
X"04803d0d",
X"72842983",
X"e2fc0570",
X"0883e080",
X"0c51823d",
X"0d04fe3d",
X"0d800b83",
X"e2e00c80",
X"0b83e2dc",
X"0cff0b83",
X"e0d80ca8",
X"0b83e2f8",
X"0cae518c",
X"a53f800b",
X"83e2fc54",
X"52807370",
X"8405550c",
X"81125271",
X"842e0981",
X"06ef3884",
X"3d0d04fe",
X"3d0d7402",
X"84059605",
X"22535371",
X"802e9638",
X"72708105",
X"5433518c",
X"c43fff12",
X"7083ffff",
X"065152e7",
X"39843d0d",
X"04fe3d0d",
X"02920522",
X"5382ac51",
X"dfa23f80",
X"c3518ca1",
X"3f819651",
X"df963f72",
X"5283e0dc",
X"51ffb43f",
X"725283e0",
X"dc51f8e6",
X"3f83e080",
X"0881ff06",
X"518bfe3f",
X"843d0d04",
X"ffb13d0d",
X"80d13df8",
X"0551f990",
X"3f83e2e0",
X"08810583",
X"e2e00c80",
X"cf3d33cf",
X"117081ff",
X"06515656",
X"74832688",
X"cd38758f",
X"06ff0556",
X"7583e0d8",
X"082e9b38",
X"75832696",
X"387583e0",
X"d80c7584",
X"2983e2fc",
X"05700853",
X"557551fa",
X"a13f8076",
X"2488a938",
X"75842983",
X"e2fc0555",
X"7408802e",
X"889a3883",
X"e0d80884",
X"2983e2fc",
X"05700802",
X"880582b9",
X"0533525b",
X"557480d2",
X"2e849a38",
X"7480d224",
X"903874bf",
X"2e9c3874",
X"80d02e81",
X"d13887d9",
X"397480d3",
X"2e80cf38",
X"7480d72e",
X"81c03887",
X"c8390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290556",
X"568b803f",
X"80c1518a",
X"b43ff6e2",
X"3f860b83",
X"e0dc3481",
X"5283e0dc",
X"518bef3f",
X"8151fde9",
X"3f748938",
X"860b83e2",
X"f80c8739",
X"a80b83e2",
X"f80c8acf",
X"3f80c151",
X"8a833ff6",
X"b13f900b",
X"83e2f333",
X"81065656",
X"74802e83",
X"38985683",
X"e2e83383",
X"e2e93371",
X"882b0756",
X"59748180",
X"2e098106",
X"9c3883e2",
X"e63383e2",
X"e7337188",
X"2b075657",
X"ad807527",
X"8c387581",
X"80075685",
X"3975a007",
X"567583e0",
X"dc34ff0b",
X"83e0dd34",
X"e00b83e0",
X"de34800b",
X"83e0df34",
X"845283e0",
X"dc518ae6",
X"3f845186",
X"86390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290556",
X"5989c43f",
X"795194c0",
X"3f83e080",
X"08802e8a",
X"3880ce51",
X"88eb3f85",
X"dd3980c1",
X"5188e23f",
X"89ea3f87",
X"ee3f83e3",
X"8c085883",
X"75259b38",
X"83e2e833",
X"83e2e933",
X"71882b07",
X"fc177129",
X"7a058380",
X"055a5157",
X"8d397481",
X"802918ff",
X"80055881",
X"80578056",
X"76762e92",
X"3888c13f",
X"83e08008",
X"83e0dc17",
X"34811656",
X"eb3988b0",
X"3f83e080",
X"0881ff06",
X"775383e0",
X"dc5256f4",
X"dd3f83e0",
X"800881ff",
X"06557575",
X"2e098106",
X"81843888",
X"b23f80c1",
X"5187e63f",
X"88ee3f77",
X"52795192",
X"df3f805e",
X"80d13dfd",
X"f4055476",
X"5383e0dc",
X"52795190",
X"e83f0282",
X"b9053355",
X"81587480",
X"d72e0981",
X"06bc3880",
X"d13dfdf0",
X"05547653",
X"8f3d7053",
X"7a525991",
X"ee3f8056",
X"76762ea2",
X"38751983",
X"e0dc1733",
X"71337072",
X"32703070",
X"80257030",
X"7e06811d",
X"5d5e5151",
X"51525b55",
X"db3982ac",
X"51d9f13f",
X"77802e86",
X"3880c351",
X"843980ce",
X"5186e63f",
X"87ee3f85",
X"f23f83d5",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055955",
X"80705d59",
X"87893f80",
X"c15186bd",
X"3f83e2f4",
X"08792e82",
X"db3883e3",
X"940880fc",
X"055580fd",
X"527451bd",
X"c13f83e0",
X"80085b77",
X"8224b238",
X"ff187087",
X"2b83ffff",
X"800680fc",
X"f00583e0",
X"dc595755",
X"81805575",
X"70810557",
X"33777081",
X"055934ff",
X"157081ff",
X"06515574",
X"ea38828a",
X"397782e8",
X"2e81aa38",
X"7782e92e",
X"09810681",
X"b13880fb",
X"88518cd4",
X"3f785877",
X"87327030",
X"70720780",
X"257a8a32",
X"70307072",
X"07802573",
X"0753545a",
X"51575575",
X"802e9738",
X"78782692",
X"38a00b83",
X"e0dc1a34",
X"81197081",
X"ff065a55",
X"eb398118",
X"7081ff06",
X"59558a78",
X"27ffbc38",
X"8f5883e0",
X"d7183383",
X"e0dc1934",
X"ff187081",
X"ff065955",
X"778426ea",
X"38905880",
X"0b83e0dc",
X"19348118",
X"7081ff06",
X"70982b52",
X"59557480",
X"25e93880",
X"c6557a85",
X"8f248438",
X"80c25574",
X"83e0dc34",
X"80f10b83",
X"e0df3481",
X"0b83e0e0",
X"347a83e0",
X"dd347a88",
X"2c557483",
X"e0de3480",
X"c93982f0",
X"782580c2",
X"387780fd",
X"29fd97d3",
X"05527951",
X"8f963f80",
X"d13dfdec",
X"055480fd",
X"5383e0dc",
X"5279518e",
X"ca3f7b81",
X"19595675",
X"80fc2483",
X"38785877",
X"882c5574",
X"83e1d934",
X"7783e1da",
X"347583e1",
X"db348180",
X"5980ca39",
X"83e38c08",
X"57837825",
X"9b3883e2",
X"e83383e2",
X"e9337188",
X"2b07fc1a",
X"71297905",
X"83800559",
X"51598d39",
X"77818029",
X"17ff8005",
X"57818059",
X"76527951",
X"8ea63f80",
X"d13dfdec",
X"05547853",
X"83e0dc52",
X"79518ddb",
X"3f7851f6",
X"d83f8494",
X"3f82983f",
X"8b3983e2",
X"dc088105",
X"83e2dc0c",
X"80d13d0d",
X"04f6f93f",
X"dfc53ff9",
X"39fc3d0d",
X"76787184",
X"2983e2fc",
X"05700851",
X"53535370",
X"9e3880ce",
X"723480cf",
X"0b811334",
X"80ce0b82",
X"133480c5",
X"0b831334",
X"70841334",
X"80e73983",
X"e3901333",
X"5480d272",
X"3473822a",
X"70810651",
X"5180cf53",
X"70843880",
X"d7537281",
X"1334a00b",
X"82133473",
X"83065170",
X"812e9e38",
X"70812488",
X"3870802e",
X"8f389f39",
X"70822e92",
X"3870832e",
X"92389339",
X"80d8558e",
X"3980d355",
X"893980cd",
X"55843980",
X"c4557483",
X"133480c4",
X"0b841334",
X"800b8513",
X"34863d0d",
X"04fe3d0d",
X"80fc8808",
X"70337081",
X"ff067084",
X"2a813281",
X"06555152",
X"5371802e",
X"8c38a873",
X"3480fc88",
X"0851b871",
X"347183e0",
X"800c843d",
X"0d04fe3d",
X"0d80fc88",
X"08703370",
X"81ff0670",
X"852a8132",
X"81065551",
X"52537180",
X"2e8c3898",
X"733480fc",
X"880851b8",
X"71347183",
X"e0800c84",
X"3d0d0480",
X"3d0d80fc",
X"84085193",
X"713480fc",
X"900851ff",
X"7134823d",
X"0d04fe3d",
X"0d029305",
X"3380fc84",
X"08535380",
X"72348a51",
X"d3be3fd3",
X"3f80fc94",
X"085280f8",
X"723480fc",
X"ac085280",
X"7234fa13",
X"80fcb408",
X"53537272",
X"3480fc9c",
X"08528072",
X"3480fca4",
X"08527272",
X"3480fc88",
X"08528072",
X"3480fc88",
X"0852b872",
X"34843d0d",
X"04ff3d0d",
X"028f0533",
X"80fc8c08",
X"52527171",
X"34fe9e3f",
X"83e08008",
X"802ef638",
X"833d0d04",
X"803d0d84",
X"39dcb03f",
X"feb83f83",
X"e0800880",
X"2ef33880",
X"fc8c0870",
X"337081ff",
X"0683e080",
X"0c515182",
X"3d0d0480",
X"3d0d80fc",
X"840851a3",
X"713480fc",
X"900851ff",
X"713480fc",
X"880851a8",
X"713480fc",
X"880851b8",
X"7134823d",
X"0d04803d",
X"0d80fc84",
X"08703370",
X"81c00670",
X"30708025",
X"83e0800c",
X"51515151",
X"823d0d04",
X"ff3d0d80",
X"fc880870",
X"337081ff",
X"0670832a",
X"81327081",
X"06515151",
X"52527080",
X"2ee538b0",
X"723480fc",
X"880851b8",
X"7134833d",
X"0d04803d",
X"0d80fcc0",
X"08700881",
X"0683e080",
X"0c51823d",
X"0d04fd3d",
X"0d757754",
X"54807325",
X"94387370",
X"81055533",
X"5280fb90",
X"51859d3f",
X"ff1353e9",
X"39853d0d",
X"04f63d0d",
X"7c7e6062",
X"5a5d5b56",
X"80598155",
X"8539747a",
X"29557452",
X"7551b592",
X"3f83e080",
X"087a27ee",
X"3874802e",
X"80dd3874",
X"527551b4",
X"fd3f83e0",
X"80087553",
X"765254b5",
X"a43f83e0",
X"80087a53",
X"755256b4",
X"e53f83e0",
X"80087930",
X"707b079f",
X"2a707780",
X"24075151",
X"54557287",
X"3883e080",
X"08c53876",
X"8118b016",
X"55585889",
X"74258b38",
X"b714537a",
X"853880d7",
X"14537278",
X"34811959",
X"ff9f3980",
X"77348c3d",
X"0d04f73d",
X"0d7b7d7f",
X"62029005",
X"bb053357",
X"59565a5a",
X"b0587283",
X"38a05875",
X"70708105",
X"52337159",
X"54559039",
X"8074258e",
X"38ff1477",
X"70810559",
X"33545472",
X"ef3873ff",
X"15555380",
X"73258938",
X"77527951",
X"782def39",
X"75337557",
X"5372802e",
X"90387252",
X"7951782d",
X"75708105",
X"573353ed",
X"398b3d0d",
X"04ee3d0d",
X"64666969",
X"70708105",
X"52335b4a",
X"5c5e5e76",
X"802e82f9",
X"3876a52e",
X"09810682",
X"e0388070",
X"41677070",
X"81055233",
X"714a5957",
X"5f76b02e",
X"0981068c",
X"38757081",
X"05573376",
X"4857815f",
X"d0175675",
X"892680da",
X"3876675c",
X"59805c93",
X"39778a24",
X"80c3387b",
X"8a29187b",
X"7081055d",
X"335a5cd0",
X"197081ff",
X"06585889",
X"7727a438",
X"ff9f1970",
X"81ff06ff",
X"a91b5a51",
X"56857627",
X"9238ffbf",
X"197081ff",
X"06515675",
X"85268a38",
X"c9195877",
X"8025ffb9",
X"387a477b",
X"407881ff",
X"06577680",
X"e42e80e5",
X"387680e4",
X"24a73876",
X"80d82e81",
X"86387680",
X"d8249038",
X"76802e81",
X"cc3876a5",
X"2e81b638",
X"81b93976",
X"80e32e81",
X"8c3881af",
X"397680f5",
X"2e9b3876",
X"80f5248b",
X"387680f3",
X"2e818138",
X"81993976",
X"80f82e80",
X"ca38818f",
X"39913d70",
X"55578053",
X"8a527984",
X"1b710853",
X"5b56fc81",
X"3f7655ab",
X"3979841b",
X"7108943d",
X"705b5b52",
X"5b567580",
X"258c3875",
X"3056ad78",
X"340280c1",
X"05577654",
X"80538a52",
X"7551fbd5",
X"3f77557e",
X"54b83991",
X"3d705577",
X"80d83270",
X"30708025",
X"56515856",
X"90527984",
X"1b710853",
X"5b57fbb1",
X"3f7555db",
X"3979841b",
X"83123354",
X"5b569839",
X"79841b71",
X"08575b56",
X"80547f53",
X"7c527d51",
X"fc9c3f87",
X"3976527d",
X"517c2d66",
X"70335881",
X"0547fd83",
X"39943d0d",
X"047283e0",
X"900c7183",
X"e0940c04",
X"fb3d0d88",
X"3d707084",
X"05520857",
X"54755383",
X"e0900852",
X"83e09408",
X"51fcc63f",
X"873d0d04",
X"ff3d0d73",
X"70085351",
X"02930533",
X"72347008",
X"8105710c",
X"833d0d04",
X"fc3d0d87",
X"3d881155",
X"785480c0",
X"a85351fc",
X"983f8052",
X"873d51d0",
X"3f863d0d",
X"04fd3d0d",
X"75705254",
X"a58e3f83",
X"e0800814",
X"5372742e",
X"9238ff13",
X"70335353",
X"71af2e09",
X"8106ee38",
X"81135372",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"77705354",
X"54c73f83",
X"e0800873",
X"2ea13883",
X"e0800873",
X"3152ff12",
X"5271ff2e",
X"8f387270",
X"81055433",
X"74708105",
X"5634eb39",
X"ff145480",
X"7434853d",
X"0d04803d",
X"0d7251ff",
X"903f823d",
X"0d047183",
X"e0800c04",
X"803d0d72",
X"51807134",
X"810bbc12",
X"0c800b80",
X"c0120c82",
X"3d0d0480",
X"0b83e5bc",
X"08248a38",
X"a5f83fff",
X"0b83e5bc",
X"0c800b83",
X"e0800c04",
X"ff3d0d73",
X"5283e398",
X"08722e8d",
X"38d93f71",
X"5197853f",
X"7183e398",
X"0c833d0d",
X"04f43d0d",
X"7e60625c",
X"5a558154",
X"bc150881",
X"91387451",
X"cf3f7958",
X"807a2580",
X"f73883e5",
X"ec087089",
X"2a5783ff",
X"06788480",
X"72315656",
X"57737825",
X"83387355",
X"7583e5bc",
X"082e8438",
X"ff893f83",
X"e5bc0880",
X"25a63875",
X"892b5199",
X"f13f83e5",
X"ec088f3d",
X"fc11555c",
X"548152f8",
X"1b5197d6",
X"3f761483",
X"e5ec0c75",
X"83e5bc0c",
X"74537652",
X"7851a4a9",
X"3f83e080",
X"0883e5ec",
X"081683e5",
X"ec0c7876",
X"31761b5b",
X"59567780",
X"24ff8b38",
X"617a710c",
X"54755475",
X"802e8338",
X"81547383",
X"e0800c8e",
X"3d0d04fc",
X"3d0dfe9b",
X"3f7651fe",
X"af3f863d",
X"fc055302",
X"a2052252",
X"775196f6",
X"3f79863d",
X"22710c54",
X"83e08008",
X"5483e080",
X"08802e83",
X"38815473",
X"83e0800c",
X"863d0d04",
X"fd3d0d76",
X"83e5bc08",
X"53538072",
X"24893871",
X"732e8438",
X"fdd13f75",
X"51fde53f",
X"725198be",
X"3f735273",
X"802e8338",
X"81527183",
X"e0800c85",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"e0800c51",
X"823d0d04",
X"80c40b83",
X"e0800c04",
X"fd3d0d75",
X"77715470",
X"535553a0",
X"e73f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfcec3f",
X"73519498",
X"3f7383e3",
X"980c83e0",
X"80085383",
X"e0800880",
X"2e833881",
X"537283e0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcc03f",
X"72802ea5",
X"38bc1308",
X"5273519f",
X"f13f83e0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"e0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83e0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83e5bc",
X"0c7483e3",
X"9c0c7583",
X"e5b80ca0",
X"de3f83e0",
X"800881ff",
X"06528153",
X"71993883",
X"e5d4518f",
X"903f83e0",
X"80085283",
X"e0800880",
X"2e833872",
X"52715372",
X"83e0800c",
X"843d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"519de23f",
X"83e08008",
X"557483e0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"e0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283e5b8",
X"0851a89e",
X"3f83e080",
X"0857f9e3",
X"3f795283",
X"e5c05196",
X"c73f83e0",
X"80085380",
X"5483e080",
X"08742e09",
X"81068283",
X"3883e39c",
X"080b0b80",
X"fad85370",
X"52559da0",
X"3f0b0b80",
X"fad85280",
X"c015519d",
X"933f74bc",
X"160c7282",
X"c0160c81",
X"0b82c416",
X"0c810b82",
X"c8160cff",
X"17735757",
X"81973983",
X"e3a83370",
X"822a7081",
X"06515454",
X"72818638",
X"73812a81",
X"06587780",
X"fc387680",
X"2e819038",
X"82d015ff",
X"1875842a",
X"810682c4",
X"130c83e3",
X"a8338106",
X"82c8130c",
X"7b547153",
X"58569cb4",
X"3f75519c",
X"cb3f83e0",
X"80081653",
X"af737081",
X"05553472",
X"bc170c83",
X"e3a95272",
X"519c953f",
X"83e3a008",
X"82c0170c",
X"83e3b652",
X"83901551",
X"9c823f77",
X"82cc170c",
X"78802e8d",
X"38755178",
X"2d83e080",
X"08802e8d",
X"3874802e",
X"86387582",
X"cc160c75",
X"5583e3a0",
X"5283e5c0",
X"5195e73f",
X"83e08008",
X"8a3883e3",
X"a9335372",
X"fed13880",
X"0b82cc17",
X"0c78802e",
X"893883e3",
X"9c0851fc",
X"b93f83e3",
X"9c085473",
X"83e0800c",
X"8b3d0d04",
X"ff3d0d80",
X"527351fd",
X"b63f833d",
X"0d04f03d",
X"0d627052",
X"54f6923f",
X"83e08008",
X"7453873d",
X"70535555",
X"f6b23ff7",
X"923f7351",
X"d33f6353",
X"745283e0",
X"800851fa",
X"b93f923d",
X"0d047183",
X"e0800c04",
X"80c01283",
X"e0800c04",
X"803d0d72",
X"82c01108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"7282cc11",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282c4",
X"110883e0",
X"800c5182",
X"3d0d04f6",
X"3d0d7c83",
X"e0980859",
X"59817927",
X"82a93878",
X"88190827",
X"82a13877",
X"33567582",
X"2e819b38",
X"75822489",
X"3875812e",
X"8d38828b",
X"3975832e",
X"81b73882",
X"82397883",
X"ffff0670",
X"812a1170",
X"83ffff06",
X"7083ff06",
X"71892a90",
X"3d5f525a",
X"51515576",
X"83ff2e8e",
X"38825476",
X"538c1808",
X"15527951",
X"a9397554",
X"76538c18",
X"08155279",
X"519ad83f",
X"83e08008",
X"81bd3875",
X"5483e080",
X"08538c18",
X"08158105",
X"528c3dfd",
X"05519abb",
X"3f83e080",
X"0881a038",
X"02a90533",
X"8c3d3371",
X"882b077a",
X"81067184",
X"2a535758",
X"56748638",
X"769fff06",
X"56755581",
X"80397554",
X"781083fe",
X"06537888",
X"2a8c1908",
X"05528c3d",
X"fc055199",
X"fa3f83e0",
X"800880df",
X"3802a905",
X"338c3d33",
X"71882b07",
X"565780d1",
X"39845478",
X"822b83fc",
X"06537887",
X"2a8c1908",
X"05528c3d",
X"fc055199",
X"ca3f83e0",
X"8008b038",
X"02ab0533",
X"028405aa",
X"05337198",
X"2b71902b",
X"07028c05",
X"a9053370",
X"882b7207",
X"903d3371",
X"80fffffe",
X"80060751",
X"52535758",
X"56833981",
X"557483e0",
X"800c8c3d",
X"0d04fb3d",
X"0d83e098",
X"08fe1988",
X"1208fe05",
X"55565480",
X"56747327",
X"8d388214",
X"33757129",
X"94160805",
X"57537583",
X"e0800c87",
X"3d0d04fc",
X"3d0d7683",
X"e0980855",
X"55807523",
X"88150853",
X"72812e88",
X"38881408",
X"73268538",
X"8152b239",
X"72903873",
X"33527183",
X"2e098106",
X"85389014",
X"0853728c",
X"160c7280",
X"2e8d3872",
X"51ff933f",
X"83e08008",
X"52853990",
X"14085271",
X"90160c80",
X"527183e0",
X"800c863d",
X"0d04fa3d",
X"0d7883e0",
X"98087122",
X"81057083",
X"ffff0657",
X"54575573",
X"802e8838",
X"90150853",
X"72863883",
X"5280e739",
X"738f0652",
X"7180da38",
X"81139016",
X"0c8c1508",
X"53729038",
X"830b8417",
X"22575273",
X"762780c6",
X"38bf3982",
X"1633ff05",
X"74842a06",
X"5271b238",
X"7251fbdb",
X"3f815271",
X"83e08008",
X"27a83883",
X"5283e080",
X"08881708",
X"279c3883",
X"e080088c",
X"160c83e0",
X"800851fd",
X"f93f83e0",
X"80089016",
X"0c737523",
X"80527183",
X"e0800c88",
X"3d0d04f2",
X"3d0d6062",
X"64585d5b",
X"75335574",
X"a02e0981",
X"06883881",
X"16704456",
X"ef396270",
X"33565674",
X"af2e0981",
X"06843881",
X"1643800b",
X"881c0c62",
X"70335155",
X"74a02691",
X"387a51fd",
X"d23f83e0",
X"80085680",
X"7c3483a8",
X"39933d84",
X"1c087058",
X"5a5f8a55",
X"a0767081",
X"055834ff",
X"155574ff",
X"2e098106",
X"ef388070",
X"595d887f",
X"085f5a7c",
X"811e7081",
X"ff066013",
X"703370af",
X"327030a0",
X"73277180",
X"25075151",
X"525b535f",
X"57557480",
X"d83876ae",
X"2e098106",
X"83388155",
X"777a2775",
X"07557480",
X"2e9f3879",
X"88327030",
X"78ae3270",
X"30707307",
X"9f2a5351",
X"57515675",
X"ac388858",
X"8b5affab",
X"39ff9f17",
X"55749926",
X"8938e017",
X"7081ff06",
X"58557781",
X"197081ff",
X"06721c53",
X"5a575576",
X"7534ff87",
X"397c1e7f",
X"0c805576",
X"a0268338",
X"8155748b",
X"1a347a51",
X"fc913f83",
X"e0800880",
X"f538a054",
X"7a227085",
X"2b83e006",
X"5455901b",
X"08527b51",
X"94d13f83",
X"e0800857",
X"83e08008",
X"8182387b",
X"33557480",
X"2e80f538",
X"8b1c3370",
X"832a7081",
X"06515656",
X"74b4388b",
X"7c841d08",
X"83e08008",
X"595b5b58",
X"ff185877",
X"ff2e9a38",
X"79708105",
X"5b337970",
X"81055b33",
X"71713152",
X"56567580",
X"2ee23886",
X"3975802e",
X"bc387a51",
X"fbf43fff",
X"863983e0",
X"80085683",
X"e0800880",
X"2ea93883",
X"e0800883",
X"2e098106",
X"80de3884",
X"1b088b11",
X"33515574",
X"80d23884",
X"5680cd39",
X"8356ec39",
X"815680c4",
X"39765684",
X"1b088b11",
X"33515574",
X"b7388b1c",
X"3370842a",
X"70810651",
X"56577480",
X"2ed53895",
X"1c33941d",
X"3371982b",
X"71902b07",
X"9b1f337f",
X"9a053371",
X"882b0772",
X"077f8805",
X"0c5a5856",
X"58fcda39",
X"7583e080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"5192e03f",
X"835683e0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"5192b43f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"7651928b",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583e080",
X"0c8a3d0d",
X"04ec3d0d",
X"6659800b",
X"83e0980c",
X"78567880",
X"2e83e838",
X"91a53f83",
X"e0800881",
X"06558256",
X"7483d838",
X"7475538e",
X"3d705358",
X"58fec23f",
X"83e08008",
X"81ff0656",
X"75812e09",
X"810680d4",
X"38905483",
X"be537452",
X"76519197",
X"3f83e080",
X"0880c938",
X"8e3d3355",
X"74802e80",
X"c93802bb",
X"05330284",
X"05ba0533",
X"71982b71",
X"902b0702",
X"8c05b905",
X"3370882b",
X"7207943d",
X"33710770",
X"587c5754",
X"525d5759",
X"56fde63f",
X"83e08008",
X"81ff0656",
X"75832e09",
X"81068638",
X"815682db",
X"3975802e",
X"86388756",
X"82d139a4",
X"548d5377",
X"52765190",
X"ae3f8156",
X"83e08008",
X"82bd3802",
X"ba053302",
X"8405b905",
X"3371882b",
X"07585c76",
X"ab380280",
X"ca053302",
X"840580c9",
X"05337198",
X"2b71902b",
X"07963d33",
X"70882b72",
X"07029405",
X"80c70533",
X"71075452",
X"5d575856",
X"02b30533",
X"77712902",
X"8805b205",
X"33028c05",
X"b1053371",
X"882b0770",
X"1c708c1f",
X"0c5e5957",
X"585c8d3d",
X"33821a34",
X"02b50533",
X"8f3d3371",
X"882b0759",
X"5b77841a",
X"2302b705",
X"33028405",
X"b6053371",
X"882b0756",
X"5b74ab38",
X"0280c605",
X"33028405",
X"80c50533",
X"71982b71",
X"902b0795",
X"3d337088",
X"2b720702",
X"940580c3",
X"05337107",
X"51525357",
X"5d5b7476",
X"31773178",
X"842a8f3d",
X"33547171",
X"31535656",
X"98803f83",
X"e0800882",
X"0570881b",
X"0c709ff6",
X"26810557",
X"5583fff6",
X"75278338",
X"83567579",
X"3475832e",
X"098106af",
X"380280d2",
X"05330284",
X"0580d105",
X"3371982b",
X"71902b07",
X"983d3370",
X"882b7207",
X"02940580",
X"cf053371",
X"07901f0c",
X"525d5759",
X"56863976",
X"1a901a0c",
X"8419228c",
X"1a081871",
X"842a0594",
X"1b0c5c80",
X"0b811a34",
X"7883e098",
X"0c805675",
X"83e0800c",
X"963d0d04",
X"e93d0d83",
X"e0980856",
X"86547580",
X"2e81a638",
X"800b8117",
X"34993de0",
X"11466a54",
X"c01153ec",
X"0551f6cf",
X"3f83e080",
X"085483e0",
X"80088185",
X"38893d33",
X"5473802e",
X"933802ab",
X"05337084",
X"2a708106",
X"51555573",
X"802e8638",
X"835480e5",
X"3902b505",
X"338f3d33",
X"71982b71",
X"902b0702",
X"8c05bb05",
X"33029005",
X"ba053371",
X"882b0772",
X"07a01b0c",
X"029005bf",
X"05330294",
X"05be0533",
X"71982b71",
X"902b0702",
X"9c05bd05",
X"3370882b",
X"7207993d",
X"3371077f",
X"9c050c52",
X"83e08008",
X"981f0c56",
X"5a525253",
X"57595781",
X"0b811734",
X"83e08008",
X"547383e0",
X"800c993d",
X"0d04f53d",
X"0d7d6002",
X"8805ba05",
X"227283e0",
X"98085b5d",
X"5a5c5c80",
X"7b238656",
X"76802e81",
X"e0388117",
X"33810655",
X"85567480",
X"2e81d238",
X"9c170898",
X"18083155",
X"74782787",
X"387483ff",
X"ff065877",
X"802e81ae",
X"38981708",
X"7083ff06",
X"56567480",
X"ca388217",
X"33ff0576",
X"892a0670",
X"81ff065a",
X"5578a038",
X"758738a0",
X"1708558d",
X"39a41708",
X"51efe03f",
X"83e08008",
X"55817527",
X"80f83874",
X"a4180ca4",
X"170851f2",
X"8d3f83e0",
X"8008802e",
X"80e43883",
X"e0800819",
X"a8180c98",
X"170883ff",
X"06848071",
X"317083ff",
X"ff065851",
X"55777627",
X"83387756",
X"75549817",
X"0883ff06",
X"53a81708",
X"5279557b",
X"83387b55",
X"74518ad3",
X"3f83e080",
X"08a43898",
X"17081698",
X"180c751a",
X"78773170",
X"83ffff06",
X"7d227905",
X"525a565a",
X"747b23fe",
X"ce398056",
X"8839800b",
X"81183481",
X"567583e0",
X"800c8d3d",
X"0d04fa3d",
X"0d7883e0",
X"98085556",
X"86557380",
X"2e81dc38",
X"81143381",
X"06538555",
X"72802e81",
X"ce389c14",
X"08537276",
X"27833872",
X"56981408",
X"57800b98",
X"150c7580",
X"2e81a938",
X"82143370",
X"892b5653",
X"76802eb5",
X"387452ff",
X"165192ee",
X"3f83e080",
X"08ff1876",
X"54705358",
X"5392df3f",
X"83e08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b4387251",
X"edc13f83",
X"e0800853",
X"810b83e0",
X"80082780",
X"cb3883e0",
X"80088815",
X"082780c0",
X"3883e080",
X"08a4150c",
X"98140815",
X"98150c75",
X"753156c9",
X"39981408",
X"16709816",
X"0c735256",
X"efc83f83",
X"e0800880",
X"2e963882",
X"1433ff05",
X"76892a06",
X"83e08008",
X"05a8150c",
X"80558839",
X"800b8115",
X"34815574",
X"83e0800c",
X"883d0d04",
X"ee3d0d64",
X"56865583",
X"e0980880",
X"2e80f638",
X"943df411",
X"84180c66",
X"54d40552",
X"7551f197",
X"3f83e080",
X"085583e0",
X"800880cf",
X"38893d33",
X"5473802e",
X"bc3802ab",
X"05337084",
X"2a708106",
X"51555584",
X"5573802e",
X"bc3802b5",
X"05338f3d",
X"3371982b",
X"71902b07",
X"028c05bb",
X"05330290",
X"05ba0533",
X"71882b07",
X"7207881b",
X"0c535759",
X"577551ee",
X"d23f83e0",
X"80085574",
X"832e0981",
X"06833884",
X"557483e0",
X"800c943d",
X"0d04e43d",
X"0d6ea13d",
X"08405d86",
X"5683e098",
X"08802e84",
X"9b389e3d",
X"f405841e",
X"0c7e9838",
X"7c51ee97",
X"3f83e080",
X"08568484",
X"39814182",
X"80398341",
X"81fb3993",
X"3d7f9605",
X"4159807f",
X"8295055f",
X"56756081",
X"ff053483",
X"41901d08",
X"762e81dd",
X"38a0547c",
X"2270852b",
X"83e00654",
X"58901d08",
X"52785186",
X"ae3f83e0",
X"80084183",
X"e08008ff",
X"b8387833",
X"5c7b802e",
X"ffb4388b",
X"193370bf",
X"06718106",
X"52435574",
X"802e80e8",
X"387b81bf",
X"0655748f",
X"2480dd38",
X"9a193355",
X"7480d538",
X"9c193355",
X"74802e80",
X"cb38f31e",
X"70585e81",
X"56758b2e",
X"09810685",
X"388e568b",
X"39759a2e",
X"09810683",
X"389c5675",
X"19707081",
X"05523371",
X"33811a82",
X"1a5f5b52",
X"5b557486",
X"38797734",
X"853980df",
X"7734777b",
X"57577aa0",
X"2e098106",
X"c0388156",
X"7b81e532",
X"7030709f",
X"2a515155",
X"7bae2e93",
X"3874802e",
X"8e386183",
X"2a708106",
X"51557480",
X"2e97387c",
X"51ecf73f",
X"83e08008",
X"4183e080",
X"08873890",
X"1d08fea5",
X"38806034",
X"75802e88",
X"387d527f",
X"5183b13f",
X"60802e86",
X"38800b90",
X"1e0c6056",
X"60832e09",
X"81068838",
X"800b901e",
X"0c853960",
X"81d23889",
X"1f57901d",
X"08802e81",
X"a8388056",
X"75197033",
X"515574a0",
X"2ea03874",
X"852e0981",
X"06843881",
X"e5557477",
X"70810559",
X"34811670",
X"81ff0657",
X"55877627",
X"d7388819",
X"335574a0",
X"2ea938ae",
X"77708105",
X"59348856",
X"75197033",
X"515574a0",
X"2e953874",
X"77708105",
X"59348116",
X"7081ff06",
X"57558a76",
X"27e2388b",
X"19337f88",
X"05349f19",
X"339e1a33",
X"71982b71",
X"902b079d",
X"1c337088",
X"2b72079c",
X"1e337107",
X"640c5299",
X"1d33981e",
X"3371882b",
X"07535153",
X"57595674",
X"7f840523",
X"97193396",
X"1a337188",
X"2b075656",
X"747f8605",
X"23807734",
X"7c51eafe",
X"3f83e080",
X"085683e0",
X"8008832e",
X"09810688",
X"38800b90",
X"1e0c8056",
X"961f3355",
X"748a3889",
X"1f52961f",
X"5181b13f",
X"7583e080",
X"0c9e3d0d",
X"04fd3d0d",
X"75775354",
X"73335170",
X"89387133",
X"5170802e",
X"a1387333",
X"72335253",
X"72712785",
X"38ff5194",
X"39707327",
X"85388151",
X"8b398114",
X"81135354",
X"d3398051",
X"7083e080",
X"0c853d0d",
X"04fd3d0d",
X"75775454",
X"72337081",
X"ff065252",
X"70802ea3",
X"387181ff",
X"068114ff",
X"bf125354",
X"52709926",
X"8938a012",
X"7081ff06",
X"53517174",
X"70810556",
X"34d23980",
X"7434853d",
X"0d04ffbd",
X"3d0d80c6",
X"3d0852a5",
X"3d705254",
X"ffb33f80",
X"c73d0852",
X"853d7052",
X"53ffa63f",
X"72527351",
X"fedf3f80",
X"c53d0d04",
X"fe3d0d74",
X"76535371",
X"70810553",
X"33517073",
X"70810555",
X"3470f038",
X"843d0d04",
X"fe3d0d74",
X"52807233",
X"52537073",
X"2e8d3881",
X"12811471",
X"33535452",
X"70f53872",
X"83e0800c",
X"843d0d04",
X"fc3d0d76",
X"557483e6",
X"80082eaf",
X"38805374",
X"5187cd3f",
X"83e08008",
X"81ff06ff",
X"147081ff",
X"06723070",
X"9f2a5152",
X"55535472",
X"802e8438",
X"71dd3873",
X"fe387483",
X"e6800c86",
X"3d0d04ff",
X"3d0dff0b",
X"83e6800c",
X"84af3f81",
X"5187913f",
X"83e08008",
X"81ff0652",
X"71ee3881",
X"d63f7183",
X"e0800c83",
X"3d0d04fc",
X"3d0d7602",
X"8405a205",
X"22028805",
X"a605227a",
X"54555555",
X"ff823f72",
X"802ea038",
X"83e69414",
X"33757081",
X"05573481",
X"147083ff",
X"ff06ff15",
X"7083ffff",
X"06565255",
X"52dd3980",
X"0b83e080",
X"0c863d0d",
X"04fc3d0d",
X"76787a11",
X"56535580",
X"5371742e",
X"93387215",
X"51703383",
X"e6941334",
X"81128114",
X"5452ea39",
X"800b83e0",
X"800c863d",
X"0d04fd3d",
X"0d905483",
X"e6800851",
X"87803f83",
X"e0800881",
X"ff06ff15",
X"71307130",
X"7073079f",
X"2a729f2a",
X"06525552",
X"555372db",
X"38853d0d",
X"04ff3d0d",
X"83e68c08",
X"1083e684",
X"080780fc",
X"c4085271",
X"0c833d0d",
X"04800b83",
X"e68c0ce1",
X"3f04810b",
X"83e68c0c",
X"d83f04ed",
X"3f047183",
X"e6880c04",
X"803d0d80",
X"51f43f81",
X"0b83e68c",
X"0c810b83",
X"e6840cff",
X"b83f823d",
X"0d04803d",
X"0d723070",
X"74078025",
X"83e6840c",
X"51ffa23f",
X"823d0d04",
X"fe3d0d02",
X"93053380",
X"fcc80854",
X"730c80fc",
X"c4085271",
X"08708106",
X"515170f7",
X"38720870",
X"81ff0683",
X"e0800c51",
X"843d0d04",
X"803d0d81",
X"ff51cd3f",
X"83e08008",
X"81ff0683",
X"e0800c82",
X"3d0d04ff",
X"3d0d7490",
X"2b740780",
X"fcb80852",
X"710c833d",
X"0d0404fb",
X"3d0d7802",
X"84059f05",
X"3370982b",
X"55575572",
X"80259b38",
X"7580ff06",
X"56805280",
X"f751e03f",
X"83e08008",
X"81ff0654",
X"73812680",
X"ff388051",
X"fee03fff",
X"9f3f8151",
X"fed83fff",
X"973f7551",
X"fee63f74",
X"982a51fe",
X"df3f7490",
X"2a7081ff",
X"065253fe",
X"d33f7488",
X"2a7081ff",
X"065253fe",
X"c73f7481",
X"ff0651fe",
X"bf3f8155",
X"7580c02e",
X"09810686",
X"38819555",
X"8d397580",
X"c82e0981",
X"06843881",
X"87557451",
X"fe9e3f8a",
X"55fec53f",
X"83e08008",
X"81ff0670",
X"982b5454",
X"7280258c",
X"38ff1570",
X"81ff0656",
X"5374e238",
X"7383e080",
X"0c873d0d",
X"04fa3d0d",
X"fdbe3f80",
X"51fdd33f",
X"8a54fe90",
X"3fff1470",
X"81ff0655",
X"5373f338",
X"73745355",
X"80c051fe",
X"a63f83e0",
X"800881ff",
X"06547381",
X"2e098106",
X"82a13883",
X"aa5280c8",
X"51fe8c3f",
X"83e08008",
X"81ff0653",
X"72812e09",
X"810681a9",
X"38745487",
X"3d741154",
X"56fdc53f",
X"83e08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e53802",
X"9a053353",
X"72812e09",
X"810681db",
X"38029b05",
X"335380ce",
X"90547281",
X"aa2e8e38",
X"81c93980",
X"e451ff9f",
X"db3fff14",
X"5473802e",
X"81b93882",
X"0a5281e9",
X"51fda43f",
X"83e08008",
X"81ff0653",
X"72dd3872",
X"5280fa51",
X"fd913f83",
X"e0800881",
X"ff065372",
X"81913872",
X"54731653",
X"fcd23f83",
X"e0800873",
X"34811470",
X"81ff0655",
X"53837427",
X"e838873d",
X"3370862a",
X"70810651",
X"54548c55",
X"7280e438",
X"845580df",
X"39745281",
X"e951fccb",
X"3f83e080",
X"0881ff06",
X"53825581",
X"e9568173",
X"27863873",
X"5580c156",
X"80ce9054",
X"8b3980e4",
X"51ff9ecc",
X"3fff1454",
X"73802ea9",
X"38805275",
X"51fc983f",
X"83e08008",
X"81ff0653",
X"72e03884",
X"805280d0",
X"51fc843f",
X"83e08008",
X"81ff0653",
X"72802e83",
X"38805574",
X"83e69034",
X"8051fafe",
X"3ffbbd3f",
X"883d0d04",
X"fb3d0d77",
X"54800b83",
X"e6903370",
X"832a7081",
X"06515557",
X"5572752e",
X"09810685",
X"3873892b",
X"54735280",
X"d151fbbb",
X"3f83e080",
X"0881ff06",
X"5372bd38",
X"82b8c054",
X"fafe3f83",
X"e0800881",
X"ff065372",
X"81ff2e09",
X"81068938",
X"ff145473",
X"e7389f39",
X"7281fe2e",
X"09810696",
X"3883ea94",
X"5283e694",
X"51fae83f",
X"face3ffa",
X"cb3f8339",
X"81558051",
X"fa803ffa",
X"bf3f7481",
X"ff0683e0",
X"800c873d",
X"0d04fb3d",
X"0d7783e6",
X"94565481",
X"51f9e33f",
X"83e69033",
X"70832a70",
X"81065154",
X"56728538",
X"73892b54",
X"735280d8",
X"51fab43f",
X"83e08008",
X"81ff0653",
X"7280e538",
X"81ff51f9",
X"cb3f81fe",
X"51f9c53f",
X"84805374",
X"70810556",
X"3351f9b8",
X"3fff1370",
X"83ffff06",
X"515372eb",
X"387251f9",
X"a73f7251",
X"f9a23ff9",
X"cb3f83e0",
X"80089f06",
X"53a78854",
X"72852e8d",
X"389a3980",
X"e451ff9c",
X"833fff14",
X"54f9ad3f",
X"83e08008",
X"81ff2e84",
X"3873e838",
X"8051f8da",
X"3ff9993f",
X"800b83e0",
X"800c873d",
X"0d0483e0",
X"8c080283",
X"e08c0cfd",
X"3d0d8053",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"83d43f83",
X"e0800870",
X"83e0800c",
X"54853d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cfd3d",
X"0d815383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"05085183",
X"a13f83e0",
X"80087083",
X"e0800c54",
X"853d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cf93d0d",
X"800b83e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"8025b938",
X"83e08c08",
X"88050830",
X"83e08c08",
X"88050c80",
X"0b83e08c",
X"08f4050c",
X"83e08c08",
X"fc05088a",
X"38810b83",
X"e08c08f4",
X"050c83e0",
X"8c08f405",
X"0883e08c",
X"08fc050c",
X"83e08c08",
X"8c050880",
X"25b93883",
X"e08c088c",
X"05083083",
X"e08c088c",
X"050c800b",
X"83e08c08",
X"f0050c83",
X"e08c08fc",
X"05088a38",
X"810b83e0",
X"8c08f005",
X"0c83e08c",
X"08f00508",
X"83e08c08",
X"fc050c80",
X"5383e08c",
X"088c0508",
X"5283e08c",
X"08880508",
X"5181df3f",
X"83e08008",
X"7083e08c",
X"08f8050c",
X"5483e08c",
X"08fc0508",
X"802e9038",
X"83e08c08",
X"f8050830",
X"83e08c08",
X"f8050c83",
X"e08c08f8",
X"05087083",
X"e0800c54",
X"893d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"800b83e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"80259938",
X"83e08c08",
X"88050830",
X"83e08c08",
X"88050c81",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"8c050880",
X"25903883",
X"e08c088c",
X"05083083",
X"e08c088c",
X"050c8153",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"bd3f83e0",
X"80087083",
X"e08c08f8",
X"050c5483",
X"e08c08fc",
X"0508802e",
X"903883e0",
X"8c08f805",
X"083083e0",
X"8c08f805",
X"0c83e08c",
X"08f80508",
X"7083e080",
X"0c54873d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cfd",
X"3d0d810b",
X"83e08c08",
X"fc050c80",
X"0b83e08c",
X"08f8050c",
X"83e08c08",
X"8c050883",
X"e08c0888",
X"050827b9",
X"3883e08c",
X"08fc0508",
X"802eae38",
X"800b83e0",
X"8c088c05",
X"0824a238",
X"83e08c08",
X"8c050810",
X"83e08c08",
X"8c050c83",
X"e08c08fc",
X"05081083",
X"e08c08fc",
X"050cffb8",
X"3983e08c",
X"08fc0508",
X"802e80e1",
X"3883e08c",
X"088c0508",
X"83e08c08",
X"88050826",
X"ad3883e0",
X"8c088805",
X"0883e08c",
X"088c0508",
X"3183e08c",
X"0888050c",
X"83e08c08",
X"f8050883",
X"e08c08fc",
X"05080783",
X"e08c08f8",
X"050c83e0",
X"8c08fc05",
X"08812a83",
X"e08c08fc",
X"050c83e0",
X"8c088c05",
X"08812a83",
X"e08c088c",
X"050cff95",
X"3983e08c",
X"08900508",
X"802e9338",
X"83e08c08",
X"88050870",
X"83e08c08",
X"f4050c51",
X"913983e0",
X"8c08f805",
X"087083e0",
X"8c08f405",
X"0c5183e0",
X"8c08f405",
X"0883e080",
X"0c853d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cff3d",
X"0d800b83",
X"e08c08fc",
X"050c83e0",
X"8c088805",
X"088106ff",
X"11700970",
X"83e08c08",
X"8c050806",
X"83e08c08",
X"fc050811",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"0508812a",
X"83e08c08",
X"88050c83",
X"e08c088c",
X"05081083",
X"e08c088c",
X"050c5151",
X"515183e0",
X"8c088805",
X"08802e84",
X"38ffab39",
X"83e08c08",
X"fc050870",
X"83e0800c",
X"51833d0d",
X"83e08c0c",
X"04fc3d0d",
X"7670797b",
X"55555555",
X"8f72278c",
X"38727507",
X"83065170",
X"802ea938",
X"ff125271",
X"ff2e9838",
X"72708105",
X"54337470",
X"81055634",
X"ff125271",
X"ff2e0981",
X"06ea3874",
X"83e0800c",
X"863d0d04",
X"74517270",
X"84055408",
X"71708405",
X"530c7270",
X"84055408",
X"71708405",
X"530c7270",
X"84055408",
X"71708405",
X"530c7270",
X"84055408",
X"71708405",
X"530cf012",
X"52718f26",
X"c9388372",
X"27953872",
X"70840554",
X"08717084",
X"05530cfc",
X"12527183",
X"26ed3870",
X"54ff8139",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"000009a7",
X"000009e8",
X"00000a0a",
X"00000a28",
X"00000a28",
X"00000a28",
X"00000a28",
X"00000a97",
X"00000ac7",
X"70704740",
X"9c704268",
X"9c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"43617274",
X"72696467",
X"6520386b",
X"2073696d",
X"706c6500",
X"45786974",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"25732025",
X"73000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"524f4d00",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"6e616d65",
X"20000000",
X"25303278",
X"00000000",
X"00000000",
X"00000000",
X"00003c9c",
X"00003ca0",
X"00003ca8",
X"00003cb4",
X"00003cc0",
X"00003ccc",
X"00003cd8",
X"00003cdc",
X"0001d20f",
X"0001d400",
X"0001d401",
X"0001d409",
X"0001d010",
X"0001d301",
X"0001d300",
X"0001d20a",
X"0001d01b",
X"0001d016",
X"0001d019",
X"0001d018",
X"0001d017",
X"0001d01a",
X"0001d403",
X"0001d402",
X"0001d40e",
X"0004007c",
X"00040078",
X"00040074",
X"00040068",
X"00040060",
X"0004005c",
X"00040058",
X"00040054",
X"00040050",
X"0004004c",
X"00040048",
X"00040044",
X"00040040",
X"00040034",
X"00040030",
X"0004002c",
X"00040028",
X"00040024",
X"00040020",
X"0004001c",
X"00040018",
X"00040014",
X"00040010",
X"0004000c",
X"00040008",
X"00040004",
X"00040000",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"69383030",
X"00000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
