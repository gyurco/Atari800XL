
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80dd",
X"98738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80e0",
X"b80c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580d7",
X"c62d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580d5da",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80cf9904",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"775193ae",
X"3f83e080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3380e0c0",
X"0b80e0c0",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"52775192",
X"dd3f83e0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583e0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"55b3903f",
X"83e08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"811451b2",
X"a83f83e0",
X"80083070",
X"83e08008",
X"07802583",
X"e0800c53",
X"863d0d04",
X"fc3d0d76",
X"70525599",
X"c93f83e0",
X"80085481",
X"5383e080",
X"0880c738",
X"7451998c",
X"3f83e080",
X"080b0b80",
X"def85383",
X"e0800852",
X"53ff8f3f",
X"83e08008",
X"a5380b0b",
X"80defc52",
X"7251fefe",
X"3f83e080",
X"0894380b",
X"0b80df80",
X"527251fe",
X"ed3f83e0",
X"8008802e",
X"83388154",
X"73537283",
X"e0800c86",
X"3d0d04fd",
X"3d0d7570",
X"525498e2",
X"3f815383",
X"e0800898",
X"38735198",
X"ab3f83e0",
X"a0085283",
X"e0800851",
X"feb43f83",
X"e0800853",
X"7283e080",
X"0c853d0d",
X"04e03d0d",
X"a33d0870",
X"525e8ed1",
X"3f83e080",
X"0833943d",
X"56547394",
X"3880e1c4",
X"52745184",
X"c6397d52",
X"785191d4",
X"3f84d039",
X"7d518eb9",
X"3f83e080",
X"08527451",
X"8de93f83",
X"e0a80852",
X"933d7052",
X"5d94c43f",
X"83e08008",
X"59800b83",
X"e0800855",
X"5b83e080",
X"087b2e94",
X"38811b74",
X"525b97c5",
X"3f83e080",
X"085483e0",
X"8008ee38",
X"805aff7a",
X"437a427a",
X"415f7909",
X"709f2c7b",
X"065b547a",
X"7a248438",
X"ff1b5af6",
X"1a700970",
X"9f2c7206",
X"7bff125a",
X"5a525555",
X"80752595",
X"38765197",
X"843f83e0",
X"800876ff",
X"18585557",
X"738024ed",
X"38747f2e",
X"8638b8a2",
X"3f745f78",
X"ff1b7058",
X"5d58807a",
X"25953877",
X"5196da3f",
X"83e08008",
X"76ff1858",
X"55587380",
X"24ed3880",
X"0b83e3a8",
X"0c800b83",
X"e3c80c0b",
X"0b80df84",
X"518bad3f",
X"81800b83",
X"e3c80c0b",
X"0b80df8c",
X"518b9d3f",
X"a80b83e3",
X"a80c7680",
X"2e80e838",
X"83e3a808",
X"77793270",
X"30707207",
X"80257087",
X"2b83e3c8",
X"0c515678",
X"53565696",
X"8d3f83e0",
X"8008802e",
X"8a380b0b",
X"80df9451",
X"8ae23f76",
X"5195cd3f",
X"83e08008",
X"520b0b80",
X"dfc8518a",
X"cf3f7651",
X"95d33f83",
X"e0800883",
X"e3a80855",
X"57757425",
X"8638a816",
X"56f73975",
X"83e3a80c",
X"86f07624",
X"ff943887",
X"980b83e3",
X"a80c7780",
X"2eb73877",
X"5195893f",
X"83e08008",
X"78525595",
X"a93f0b0b",
X"80df9c54",
X"83e08008",
X"8f388739",
X"807634fd",
X"96390b0b",
X"80df9854",
X"74537352",
X"0b0b80de",
X"e85189e8",
X"3f80540b",
X"0b80def0",
X"5189dd3f",
X"81145473",
X"a82e0981",
X"06ed3886",
X"8da051b4",
X"a53f8052",
X"903d7052",
X"5480c2a6",
X"3f835273",
X"5180c29e",
X"3f61802e",
X"80ff387b",
X"5473ff2e",
X"96387880",
X"2e818038",
X"785194a9",
X"3f83e080",
X"08ff1555",
X"59e73978",
X"802e80eb",
X"38785194",
X"a53f83e0",
X"8008802e",
X"fc843878",
X"5193ed3f",
X"83e08008",
X"520b0b80",
X"def451ab",
X"cb3f83e0",
X"8008a438",
X"7c51ad83",
X"3f83e080",
X"085574ff",
X"16565480",
X"7425fbef",
X"38741d70",
X"33555673",
X"af2efec8",
X"38e83978",
X"5193ab3f",
X"83e08008",
X"527c51ac",
X"ba3ffbcf",
X"397f8829",
X"6010057a",
X"0561055a",
X"fc8039a2",
X"3d0d0480",
X"3d0d9080",
X"f8337081",
X"ff067084",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d38a8",
X"0b9080f8",
X"34b80b90",
X"80f83470",
X"83e0800c",
X"823d0d04",
X"803d0d90",
X"80f83370",
X"81ff0670",
X"852a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"980b9080",
X"f834b80b",
X"9080f834",
X"7083e080",
X"0c823d0d",
X"04930b90",
X"80fc34ff",
X"0b9080e8",
X"3404ff3d",
X"0d028f05",
X"3352800b",
X"9080fc34",
X"8a51b1fa",
X"3fdf3f80",
X"f80b9080",
X"e034800b",
X"9080c834",
X"fa125271",
X"9080c034",
X"800b9080",
X"d8347190",
X"80d03490",
X"80f85280",
X"7234b872",
X"34833d0d",
X"04803d0d",
X"028b0533",
X"51709080",
X"f434febf",
X"3f83e080",
X"08802ef6",
X"38823d0d",
X"04803d0d",
X"8439bae9",
X"3ffed93f",
X"83e08008",
X"802ef338",
X"9080f433",
X"7081ff06",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"a30b9080",
X"fc34ff0b",
X"9080e834",
X"9080f851",
X"a87134b8",
X"7134823d",
X"0d04803d",
X"0d9080fc",
X"337081c0",
X"06703070",
X"802583e0",
X"800c5151",
X"51823d0d",
X"04803d0d",
X"9080f833",
X"7081ff06",
X"70832a81",
X"32708106",
X"51515151",
X"70802ee8",
X"38b00b90",
X"80f834b8",
X"0b9080f8",
X"34823d0d",
X"04803d0d",
X"9080ac08",
X"810683e0",
X"800c823d",
X"0d04fd3d",
X"0d757754",
X"54807325",
X"94387370",
X"81055533",
X"5280dfa0",
X"5185a13f",
X"ff1353e9",
X"39853d0d",
X"04f63d0d",
X"7c7e6062",
X"5a5d5b56",
X"80598155",
X"8539747a",
X"29557452",
X"755180c0",
X"bf3f83e0",
X"80087a27",
X"ed387480",
X"2e80e038",
X"74527551",
X"80c0a93f",
X"83e08008",
X"75537652",
X"5480c0cf",
X"3f83e080",
X"087a5375",
X"525680c0",
X"8f3f83e0",
X"80087930",
X"707b079f",
X"2a707780",
X"24075151",
X"54557287",
X"3883e080",
X"08c23876",
X"8118b016",
X"55585889",
X"74258b38",
X"b714537a",
X"853880d7",
X"14537278",
X"34811959",
X"ff9c3980",
X"77348c3d",
X"0d04f73d",
X"0d7b7d7f",
X"62029005",
X"bb053357",
X"59565a5a",
X"b0587283",
X"38a05875",
X"70708105",
X"52337159",
X"54559039",
X"8074258e",
X"38ff1477",
X"70810559",
X"33545472",
X"ef3873ff",
X"15555380",
X"73258938",
X"77527951",
X"782def39",
X"75337557",
X"5372802e",
X"90387252",
X"7951782d",
X"75708105",
X"573353ed",
X"398b3d0d",
X"04ee3d0d",
X"64666969",
X"70708105",
X"52335b4a",
X"5c5e5e76",
X"802e82f9",
X"3876a52e",
X"09810682",
X"e0388070",
X"41677070",
X"81055233",
X"714a5957",
X"5f76b02e",
X"0981068c",
X"38757081",
X"05573376",
X"4857815f",
X"d0175675",
X"892680da",
X"3876675c",
X"59805c93",
X"39778a24",
X"80c3387b",
X"8a29187b",
X"7081055d",
X"335a5cd0",
X"197081ff",
X"06585889",
X"7727a438",
X"ff9f1970",
X"81ff06ff",
X"a91b5a51",
X"56857627",
X"9238ffbf",
X"197081ff",
X"06515675",
X"85268a38",
X"c9195877",
X"8025ffb9",
X"387a477b",
X"407881ff",
X"06577680",
X"e42e80e5",
X"387680e4",
X"24a73876",
X"80d82e81",
X"86387680",
X"d8249038",
X"76802e81",
X"cc3876a5",
X"2e81b638",
X"81b93976",
X"80e32e81",
X"8c3881af",
X"397680f5",
X"2e9b3876",
X"80f5248b",
X"387680f3",
X"2e818138",
X"81993976",
X"80f82e80",
X"ca38818f",
X"39913d70",
X"55578053",
X"8a527984",
X"1b710853",
X"5b56fbfd",
X"3f7655ab",
X"3979841b",
X"7108943d",
X"705b5b52",
X"5b567580",
X"258c3875",
X"3056ad78",
X"340280c1",
X"05577654",
X"80538a52",
X"7551fbd1",
X"3f77557e",
X"54b83991",
X"3d705577",
X"80d83270",
X"30708025",
X"56515856",
X"90527984",
X"1b710853",
X"5b57fbad",
X"3f7555db",
X"3979841b",
X"83123354",
X"5b569839",
X"79841b71",
X"08575b56",
X"80547f53",
X"7c527d51",
X"fc9c3f87",
X"3976527d",
X"517c2d66",
X"70335881",
X"0547fd83",
X"39943d0d",
X"047283e0",
X"900c7183",
X"e0940c04",
X"fb3d0d88",
X"3d707084",
X"05520857",
X"54755383",
X"e0900852",
X"83e09408",
X"51fcc63f",
X"873d0d04",
X"ff3d0d73",
X"70085351",
X"02930533",
X"72347008",
X"8105710c",
X"833d0d04",
X"fc3d0d87",
X"3d881155",
X"785499d0",
X"5351fc99",
X"3f805287",
X"3d51d13f",
X"863d0d04",
X"fd3d0d75",
X"705254a3",
X"c23f83e0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83e0",
X"8008732e",
X"a13883e0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183e0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83e2d408",
X"248a38b9",
X"a93fff0b",
X"83e2d40c",
X"800b83e0",
X"800c04ff",
X"3d0d7352",
X"83e0b008",
X"722e8d38",
X"d93f7151",
X"96973f71",
X"83e0b00c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"558154bc",
X"15088191",
X"387451cf",
X"3f795880",
X"7a2580f7",
X"3883e384",
X"0870892a",
X"5783ff06",
X"78848072",
X"31565657",
X"73782583",
X"38735575",
X"83e2d408",
X"2e8438ff",
X"893f83e2",
X"d4088025",
X"a6387589",
X"2b5198da",
X"3f83e384",
X"088f3dfc",
X"11555c54",
X"8152f81b",
X"5196c43f",
X"761483e3",
X"840c7583",
X"e2d40c74",
X"53765278",
X"51b7bc3f",
X"83e08008",
X"83e38408",
X"1683e384",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8b3861",
X"7a710c54",
X"75547580",
X"2e833881",
X"547383e0",
X"800c8e3d",
X"0d04fc3d",
X"0dfe9b3f",
X"7651feaf",
X"3f863dfc",
X"05537852",
X"775195e7",
X"3f797571",
X"0c5483e0",
X"80085483",
X"e0800880",
X"2e833881",
X"547383e0",
X"800c863d",
X"0d04fe3d",
X"0d7583e2",
X"d4085353",
X"80722489",
X"3871732e",
X"8438fdd6",
X"3f7451fd",
X"ea3f7251",
X"97ac3f83",
X"e0800852",
X"83e08008",
X"802e8338",
X"81527183",
X"e0800c84",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"e0800c51",
X"823d0d04",
X"80c40b83",
X"e0800c04",
X"fd3d0d75",
X"77715470",
X"5355539f",
X"9a3f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfceb3f",
X"735193a9",
X"3f7383e0",
X"b00c83e0",
X"80085383",
X"e0800880",
X"2e833881",
X"537283e0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcbf3f",
X"72802ea5",
X"38bc1308",
X"5273519e",
X"a43f83e0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"e0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83e0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83e2d4",
X"0c7483e0",
X"b40c7583",
X"e2d00cb4",
X"803f83e0",
X"800881ff",
X"06528153",
X"71993883",
X"e2ec518e",
X"933f83e0",
X"80085283",
X"e0800880",
X"2e833872",
X"52715372",
X"83e0800c",
X"843d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"519c953f",
X"83e08008",
X"557483e0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"e0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283e2d0",
X"0851b3c8",
X"3f83e080",
X"0857f9e2",
X"3f795283",
X"e2d85195",
X"b43f83e0",
X"80085480",
X"5383e080",
X"08732e09",
X"81068283",
X"3883e0b4",
X"080b0b80",
X"def45370",
X"52569bd3",
X"3f0b0b80",
X"def45280",
X"c016519b",
X"c63f75bc",
X"170c7382",
X"c0170c81",
X"0b82c417",
X"0c810b82",
X"c8170c73",
X"82cc170c",
X"ff1782d0",
X"17555781",
X"913983e0",
X"c0337082",
X"2a708106",
X"51545572",
X"81803874",
X"812a8106",
X"587780f6",
X"3874842a",
X"810682c4",
X"150c83e0",
X"c0338106",
X"82c8150c",
X"79527351",
X"9aed3f73",
X"519b843f",
X"83e08008",
X"1453af73",
X"70810555",
X"3472bc15",
X"0c83e0c1",
X"5272519a",
X"ce3f83e0",
X"b80882c0",
X"150c83e0",
X"ce5280c0",
X"14519abb",
X"3f78802e",
X"8d387351",
X"782d83e0",
X"8008802e",
X"99387782",
X"cc150c75",
X"802e8638",
X"7382cc17",
X"0c7382d0",
X"15ff1959",
X"55567680",
X"2e9b3883",
X"e0b85283",
X"e2d85194",
X"aa3f83e0",
X"80088a38",
X"83e0c133",
X"5372fed2",
X"3878802e",
X"893883e0",
X"b40851fc",
X"b93f83e0",
X"b4085372",
X"83e0800c",
X"8b3d0d04",
X"ff3d0d80",
X"527351fd",
X"b63f833d",
X"0d04f03d",
X"0d627052",
X"54f6913f",
X"83e08008",
X"7453873d",
X"70535555",
X"f6b13ff7",
X"913f7351",
X"d33f6353",
X"745283e0",
X"800851fa",
X"b93f923d",
X"0d047183",
X"e0800c04",
X"80c01283",
X"e0800c04",
X"803d0d72",
X"82c01108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"7282cc11",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282c4",
X"110883e0",
X"800c5182",
X"3d0d04f9",
X"3d0d7983",
X"e0980857",
X"57817727",
X"81963876",
X"88170827",
X"818e3875",
X"33557482",
X"2e893874",
X"832eb338",
X"80fe3974",
X"54761083",
X"fe065376",
X"882a8c17",
X"08055289",
X"3dfc0551",
X"ae9c3f83",
X"e0800880",
X"df38029d",
X"0533893d",
X"3371882b",
X"07565680",
X"d1398454",
X"76822b83",
X"fc065376",
X"872a8c17",
X"08055289",
X"3dfc0551",
X"adec3f83",
X"e08008b0",
X"38029f05",
X"33028405",
X"9e053371",
X"982b7190",
X"2b07028c",
X"059d0533",
X"70882b72",
X"078d3d33",
X"7180ffff",
X"fe800607",
X"51525357",
X"58568339",
X"81557483",
X"e0800c89",
X"3d0d04fb",
X"3d0d83e0",
X"9808fe19",
X"881208fe",
X"05555654",
X"80567473",
X"278d3882",
X"14337571",
X"29941608",
X"05575375",
X"83e0800c",
X"873d0d04",
X"fc3d0d76",
X"52800b83",
X"e0980870",
X"33515253",
X"70832e09",
X"81069138",
X"95123394",
X"13337198",
X"2b71902b",
X"07555551",
X"9b12339a",
X"13337188",
X"2b077407",
X"83e0800c",
X"55863d0d",
X"04fc3d0d",
X"7683e098",
X"08555580",
X"75238815",
X"08537281",
X"2e883888",
X"14087326",
X"85388152",
X"b2397290",
X"38733352",
X"71832e09",
X"81068538",
X"90140853",
X"728c160c",
X"72802e8d",
X"387251fe",
X"d63f83e0",
X"80085285",
X"39901408",
X"52719016",
X"0c805271",
X"83e0800c",
X"863d0d04",
X"fa3d0d78",
X"83e09808",
X"71228105",
X"7083ffff",
X"06575457",
X"5573802e",
X"88389015",
X"08537286",
X"38835280",
X"e739738f",
X"06527180",
X"da388113",
X"90160c8c",
X"15085372",
X"9038830b",
X"84172257",
X"52737627",
X"80c638bf",
X"39821633",
X"ff057484",
X"2a065271",
X"b2387251",
X"fcb13f81",
X"527183e0",
X"800827a8",
X"38835283",
X"e0800888",
X"1708279c",
X"3883e080",
X"088c160c",
X"83e08008",
X"51fdbc3f",
X"83e08008",
X"90160c73",
X"75238052",
X"7183e080",
X"0c883d0d",
X"04f23d0d",
X"60626458",
X"5e5b7533",
X"5574a02e",
X"09810688",
X"38811670",
X"4456ef39",
X"62703356",
X"5674af2e",
X"09810684",
X"38811643",
X"800b881c",
X"0c627033",
X"5155749f",
X"2691387a",
X"51fdd23f",
X"83e08008",
X"56807d34",
X"83813993",
X"3d841c08",
X"7058595f",
X"8a55a076",
X"70810558",
X"34ff1555",
X"74ff2e09",
X"8106ef38",
X"80705a5c",
X"887f085f",
X"5a7b811d",
X"7081ff06",
X"60137033",
X"70af3270",
X"30a07327",
X"71802507",
X"5151525b",
X"535e5755",
X"7480e738",
X"76ae2e09",
X"81068338",
X"8155787a",
X"27750755",
X"74802e9f",
X"38798832",
X"703078ae",
X"32703070",
X"73079f2a",
X"53515751",
X"5675bb38",
X"88598b5a",
X"ffab3976",
X"982b5574",
X"80258738",
X"80dca817",
X"3357ff9f",
X"17557499",
X"268938e0",
X"177081ff",
X"06585578",
X"811a7081",
X"ff06721b",
X"535b5755",
X"767534fe",
X"f8397b1e",
X"7f0c8055",
X"76a02683",
X"38815574",
X"8b19347a",
X"51fc823f",
X"83e08008",
X"80f538a0",
X"547a2270",
X"852b83e0",
X"06545590",
X"1b08527c",
X"51a8a73f",
X"83e08008",
X"5783e080",
X"08818138",
X"7c335574",
X"802e80f4",
X"388b1d33",
X"70832a70",
X"81065156",
X"5674b438",
X"8b7d841d",
X"0883e080",
X"08595b5b",
X"58ff1858",
X"77ff2e9a",
X"38797081",
X"055b3379",
X"7081055b",
X"33717131",
X"52565675",
X"802ee238",
X"86397580",
X"2e96387a",
X"51fbe53f",
X"ff863983",
X"e0800856",
X"83e08008",
X"b6388339",
X"7656841b",
X"088b1133",
X"515574a7",
X"388b1d33",
X"70842a70",
X"81065156",
X"56748938",
X"83569439",
X"81569039",
X"7c51fa94",
X"3f83e080",
X"08881c0c",
X"fd813975",
X"83e0800c",
X"903d0d04",
X"f83d0d7a",
X"7c595782",
X"5483fe53",
X"77527651",
X"a6ec3f83",
X"5683e080",
X"0880ec38",
X"81173377",
X"3371882b",
X"07565682",
X"567482d4",
X"d52e0981",
X"0680d438",
X"7554b653",
X"77527651",
X"a6c03f83",
X"e0800898",
X"38811733",
X"77337188",
X"2b0783e0",
X"80085256",
X"56748182",
X"c62eac38",
X"825480d2",
X"53775276",
X"51a6973f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62e83",
X"38815675",
X"83e0800c",
X"8a3d0d04",
X"eb3d0d67",
X"5a800b83",
X"e0980ca5",
X"cc3f83e0",
X"80088106",
X"55825674",
X"83ee3874",
X"75538f3d",
X"70535759",
X"feca3f83",
X"e0800881",
X"ff065776",
X"812e0981",
X"0680d438",
X"905483be",
X"53745275",
X"51a5ab3f",
X"83e08008",
X"80c9388f",
X"3d335574",
X"802e80c9",
X"3802bf05",
X"33028405",
X"be053371",
X"982b7190",
X"2b07028c",
X"05bd0533",
X"70882b72",
X"07953d33",
X"71077058",
X"7b575e52",
X"5e575957",
X"fdee3f83",
X"e0800881",
X"ff065776",
X"832e0981",
X"06863881",
X"5682f139",
X"76802e86",
X"38865682",
X"e739a454",
X"8d537852",
X"7551a4c2",
X"3f815683",
X"e0800882",
X"d33802be",
X"05330284",
X"05bd0533",
X"71882b07",
X"595d77ab",
X"380280ce",
X"05330284",
X"0580cd05",
X"3371982b",
X"71902b07",
X"973d3370",
X"882b7207",
X"02940580",
X"cb053371",
X"0754525e",
X"57595602",
X"b7053378",
X"71290288",
X"05b60533",
X"028c05b5",
X"05337188",
X"2b07701d",
X"707f8c05",
X"0c5f5957",
X"595d8e3d",
X"33821b34",
X"02b90533",
X"903d3371",
X"882b075a",
X"5c78841b",
X"2302bb05",
X"33028405",
X"ba053371",
X"882b0756",
X"5c74ab38",
X"0280ca05",
X"33028405",
X"80c90533",
X"71982b71",
X"902b0796",
X"3d337088",
X"2b720702",
X"940580c7",
X"05337107",
X"51525357",
X"5e5c7476",
X"31783179",
X"842a903d",
X"33547171",
X"31535656",
X"a4ae3f83",
X"e0800882",
X"0570881c",
X"0c83e080",
X"08e08a05",
X"56567483",
X"dffe2683",
X"38825783",
X"fff67627",
X"85388357",
X"89398656",
X"76802e80",
X"db38767a",
X"3476832e",
X"098106b0",
X"380280d6",
X"05330284",
X"0580d505",
X"3371982b",
X"71902b07",
X"993d3370",
X"882b7207",
X"02940580",
X"d3053371",
X"077f9005",
X"0c525e57",
X"58568639",
X"771b901b",
X"0c841a22",
X"8c1b0819",
X"71842a05",
X"941c0c5d",
X"800b811b",
X"347983e0",
X"980c8056",
X"7583e080",
X"0c973d0d",
X"04e93d0d",
X"83e09808",
X"56855475",
X"802e8182",
X"38800b81",
X"1734993d",
X"e011466a",
X"548a3d70",
X"5458ec05",
X"51f6e63f",
X"83e08008",
X"5483e080",
X"0880df38",
X"893d3354",
X"73802e91",
X"3802ab05",
X"3370842a",
X"81065155",
X"74802e86",
X"38835480",
X"c1397651",
X"f48a3f83",
X"e08008a0",
X"170c02bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"3371079c",
X"1c0c5278",
X"981b0c53",
X"56595781",
X"0b811734",
X"74547383",
X"e0800c99",
X"3d0d04f5",
X"3d0d7d7f",
X"617283e0",
X"98085a5d",
X"5d595c80",
X"7b0c8557",
X"75802e81",
X"e0388116",
X"33810655",
X"84577480",
X"2e81d238",
X"91397481",
X"17348639",
X"800b8117",
X"34815781",
X"c0399c16",
X"08981708",
X"31557478",
X"27833874",
X"5877802e",
X"81a93898",
X"16087083",
X"ff065657",
X"7480cf38",
X"821633ff",
X"0577892a",
X"067081ff",
X"065a5578",
X"a0387687",
X"38a01608",
X"558d39a4",
X"160851f0",
X"ea3f83e0",
X"80085581",
X"7527ffa8",
X"3874a417",
X"0ca41608",
X"51f2843f",
X"83e08008",
X"5583e080",
X"08802eff",
X"893883e0",
X"800819a8",
X"170c9816",
X"0883ff06",
X"84807131",
X"51557775",
X"27833877",
X"557483ff",
X"ff065498",
X"160883ff",
X"0653a816",
X"08527957",
X"7b83387b",
X"5776519e",
X"e93f83e0",
X"8008fed0",
X"38981608",
X"1598170c",
X"741a7876",
X"317c0817",
X"7d0c595a",
X"fed33980",
X"577683e0",
X"800c8d3d",
X"0d04fa3d",
X"0d7883e0",
X"98085556",
X"85557380",
X"2e81e138",
X"81143381",
X"06538455",
X"72802e81",
X"d3389c14",
X"08537276",
X"27833872",
X"56981408",
X"57800b98",
X"150c7580",
X"2e81b738",
X"82143370",
X"892b5653",
X"76802eb5",
X"387452ff",
X"16519fb0",
X"3f83e080",
X"08ff1876",
X"54705358",
X"539fa13f",
X"83e08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed93f83",
X"e0800853",
X"810b83e0",
X"8008278b",
X"38881408",
X"83e08008",
X"26883880",
X"0b811534",
X"b03983e0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc83f",
X"83e08008",
X"8c3883e0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683e0",
X"800805a8",
X"150c8055",
X"7483e080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83e09808",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1d23f",
X"83e08008",
X"5583e080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef8",
X"3f83e080",
X"0888170c",
X"7551efa9",
X"3f83e080",
X"08557483",
X"e0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683e0",
X"9808802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f83f83e0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"9af43f83",
X"e0800841",
X"83e08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"ede23f83",
X"e0800841",
X"83e08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"83a53f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f33f83e0",
X"80088332",
X"70307072",
X"079f2c83",
X"e0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"81b13f75",
X"83e0800c",
X"9e3d0d04",
X"fd3d0d75",
X"77535473",
X"33517089",
X"38713351",
X"70802ea1",
X"38733372",
X"33525372",
X"71278538",
X"ff519439",
X"70732785",
X"3881518b",
X"39811481",
X"135354d3",
X"39805170",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"77545472",
X"337081ff",
X"06525270",
X"802ea338",
X"7181ff06",
X"8114ffbf",
X"12535452",
X"70992689",
X"38a01270",
X"81ff0653",
X"51717470",
X"81055634",
X"d2398074",
X"34853d0d",
X"04ffbd3d",
X"0d80c63d",
X"0852a53d",
X"705254ff",
X"b33f80c7",
X"3d085285",
X"3d705253",
X"ffa63f72",
X"527351fe",
X"df3f80c5",
X"3d0d04fe",
X"3d0d7476",
X"53537170",
X"81055333",
X"51707370",
X"81055534",
X"70f03884",
X"3d0d04fe",
X"3d0d7452",
X"80723352",
X"5370732e",
X"8d388112",
X"81147133",
X"53545270",
X"f5387283",
X"e0800c84",
X"3d0d0471",
X"83e39c0c",
X"8880800b",
X"83e3980c",
X"8480800b",
X"83e3a00c",
X"04f03d0d",
X"83808056",
X"83e39c08",
X"1683e398",
X"08175654",
X"74337434",
X"83e3a008",
X"16548074",
X"34811656",
X"758380a0",
X"2e098106",
X"db3883d0",
X"805683e3",
X"9c081683",
X"e3980817",
X"56547433",
X"743483e3",
X"a0081654",
X"80743481",
X"16567583",
X"d0a02e09",
X"8106db38",
X"83a88056",
X"83e39c08",
X"1683e398",
X"08175654",
X"74337434",
X"83e3a008",
X"16548074",
X"34811656",
X"7583a890",
X"2e098106",
X"db388056",
X"83e39c08",
X"1683e3a0",
X"08175555",
X"73337534",
X"81165675",
X"8180802e",
X"098106e4",
X"3886c33f",
X"893d58a2",
X"5380dea8",
X"5277519c",
X"c23f8057",
X"8c805683",
X"e3a00816",
X"77195555",
X"73337534",
X"81168118",
X"585676a2",
X"2e098106",
X"e638860b",
X"87a88334",
X"800b87a8",
X"8234800b",
X"87809a34",
X"af0b8780",
X"9634bf0b",
X"87809734",
X"800b8780",
X"98349f0b",
X"87809934",
X"800b8780",
X"9b34f80b",
X"87a88934",
X"7687a880",
X"34820b87",
X"d08f3482",
X"0b87a881",
X"34923d0d",
X"04fe3d0d",
X"805383e3",
X"a0081383",
X"e39c0814",
X"52527033",
X"72348113",
X"53728180",
X"802e0981",
X"06e43883",
X"80805383",
X"e3a00813",
X"83e39c08",
X"14525270",
X"33723481",
X"13537283",
X"80a02e09",
X"8106e438",
X"83d08053",
X"83e3a008",
X"1383e39c",
X"08145252",
X"70337234",
X"81135372",
X"83d0a02e",
X"098106e4",
X"3883a880",
X"5383e3a0",
X"081383e3",
X"9c081452",
X"52703372",
X"34811353",
X"7283a890",
X"2e098106",
X"e438843d",
X"0d04803d",
X"0d908090",
X"08810683",
X"e0800c82",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe067607",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"812c8106",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fd06",
X"76100772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087082",
X"2cbf0683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fe8306",
X"76822b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"882c8706",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f1ff",
X"0676882b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"708b2cbf",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870f8",
X"8fff0676",
X"8b2b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087091",
X"2cbf0683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fc87ff",
X"ff067691",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908080",
X"0870882c",
X"810683e0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"80087089",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8a2c8106",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708b2c81",
X"0683e080",
X"0c51823d",
X"0d04fe3d",
X"0d7481e6",
X"29872a90",
X"80a00c84",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70810554",
X"34ff1151",
X"f039843d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"8405540c",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"81808053",
X"80528880",
X"0a51ffb3",
X"3fa08053",
X"80528280",
X"0a51c73f",
X"843d0d04",
X"803d0d81",
X"51fcc03f",
X"72802e83",
X"38d33f81",
X"51fcde3f",
X"8051fcd9",
X"3f8051fc",
X"aa3f823d",
X"0d04fd3d",
X"0d755280",
X"5480ff72",
X"25883881",
X"0bff8013",
X"5354ffbf",
X"12517099",
X"268638e0",
X"12529e39",
X"ff9f1251",
X"99712795",
X"38d012e0",
X"13705454",
X"51897127",
X"88388f73",
X"27833880",
X"5273802e",
X"85388180",
X"12527181",
X"ff0683e0",
X"800c853d",
X"0d04803d",
X"0d84d8c0",
X"51807170",
X"81055334",
X"7084e0c0",
X"2e098106",
X"f038823d",
X"0d04fe3d",
X"0d029705",
X"3351ff86",
X"3f83e080",
X"0881ff06",
X"83e3a808",
X"54528073",
X"249b3883",
X"e3c40813",
X"7283e3c8",
X"08075353",
X"71733483",
X"e3a80881",
X"0583e3a8",
X"0c843d0d",
X"04fa3d0d",
X"82800a1b",
X"55805788",
X"3dfc0554",
X"79537452",
X"7851d69a",
X"3f883d0d",
X"04fe3d0d",
X"83e3c008",
X"527451dc",
X"fd3f83e0",
X"80088c38",
X"76537552",
X"83e3c008",
X"51c73f84",
X"3d0d04fe",
X"3d0d83e3",
X"c0085375",
X"527451d7",
X"bd3f83e0",
X"80088d38",
X"77537652",
X"83e3c008",
X"51ffa23f",
X"843d0d04",
X"fd3d0d83",
X"e3c00851",
X"d6b13f83",
X"e0800890",
X"802e0981",
X"06ad3880",
X"5483c180",
X"805383e0",
X"80085283",
X"e3c00851",
X"fef33f87",
X"c1808014",
X"3387c190",
X"80153481",
X"14547390",
X"802e0981",
X"06e93885",
X"3d0d0480",
X"dfa80b83",
X"e0800c04",
X"f73d0d80",
X"5a805980",
X"58807057",
X"57fde73f",
X"800b83e3",
X"a80c800b",
X"83e3c80c",
X"80dfac51",
X"d1963f81",
X"800b83e3",
X"c80c80df",
X"b051d188",
X"3f80d00b",
X"83e3a80c",
X"75307077",
X"07802570",
X"872b83e3",
X"c80c5154",
X"f9bd3f83",
X"e0800852",
X"80dfb851",
X"d0e23f80",
X"f80b83e3",
X"a80c7581",
X"32703070",
X"72078025",
X"70872b83",
X"e3c80c51",
X"5555ff83",
X"3f83e080",
X"085280df",
X"c451d0b8",
X"3f81a00b",
X"83e3a80c",
X"75823270",
X"30707207",
X"80257087",
X"2b83e3c8",
X"0c515583",
X"e3c00852",
X"55d1d23f",
X"83e08008",
X"5280dfcc",
X"51d0893f",
X"81c80b83",
X"e3a80c75",
X"83327030",
X"70720780",
X"2570872b",
X"83e3c80c",
X"515580df",
X"d45255cf",
X"e73f81f0",
X"0b83e3a8",
X"0c758432",
X"70307072",
X"07802570",
X"872b83e3",
X"c80c5155",
X"80dfe452",
X"55cfc53f",
X"82980b83",
X"e3a80c75",
X"85327030",
X"70720780",
X"2570872b",
X"83e3c80c",
X"515580df",
X"fc5255cf",
X"a33f82c0",
X"0b83e3a8",
X"0c758632",
X"70307072",
X"07802570",
X"872b83e3",
X"c80c5155",
X"80e09452",
X"55cf813f",
X"868da051",
X"f9d43f80",
X"52883d70",
X"525487d6",
X"3f835273",
X"5187cf3f",
X"78165675",
X"80258538",
X"80569039",
X"86762585",
X"38865687",
X"39758626",
X"82da3875",
X"842980de",
X"cc055473",
X"0804f78f",
X"3f83e080",
X"08785654",
X"74812e09",
X"81068938",
X"83e08008",
X"10549039",
X"74ff2e09",
X"81068838",
X"83e08008",
X"812c5490",
X"74258538",
X"90548839",
X"73802483",
X"38815473",
X"51f6e93f",
X"828e39f6",
X"fb3f83e0",
X"80081854",
X"73802585",
X"38805488",
X"39877425",
X"83388754",
X"7351f6f5",
X"3f81ed39",
X"77873879",
X"802e81e4",
X"3883e0a4",
X"0883e0a0",
X"0c8bdf0b",
X"83e0a80c",
X"83e3c008",
X"51c0a23f",
X"fbb63f81",
X"c7397980",
X"2e81c138",
X"83e09c08",
X"83e0a00c",
X"8bdf0b83",
X"e0a80c83",
X"e3bc0851",
X"ffbffe3f",
X"75832e09",
X"81069438",
X"81808053",
X"82808052",
X"83e3bc08",
X"51fa9a3f",
X"81873975",
X"842e0981",
X"06af3882",
X"80805381",
X"80805283",
X"e3bc0851",
X"f9ff3f80",
X"54848280",
X"80143384",
X"81808015",
X"34811454",
X"73818080",
X"2e098106",
X"e83880d1",
X"3975852e",
X"09810680",
X"c8388054",
X"81808053",
X"80c08052",
X"83e3bc08",
X"51f9c63f",
X"82808053",
X"80c08052",
X"83e3bc08",
X"51f9b63f",
X"84818080",
X"14338481",
X"c0801534",
X"84828080",
X"14338482",
X"c0801534",
X"81145473",
X"80c0802e",
X"098106dc",
X"3881548c",
X"39798738",
X"76802efa",
X"c4388054",
X"7383e080",
X"0c8b3d0d",
X"04ff3d0d",
X"f5e43f83",
X"e0800880",
X"2e863880",
X"5180dd39",
X"f5e93f83",
X"e0800880",
X"d138f689",
X"3f83e080",
X"08802eaa",
X"388151f3",
X"c63ff08d",
X"3f800b83",
X"e3a80cf9",
X"f33f83e0",
X"800852ff",
X"0b83e3a8",
X"0cf2923f",
X"71a43871",
X"51f3a43f",
X"a239f5c0",
X"3f83e080",
X"08802e97",
X"388151f3",
X"923fefd9",
X"3fff0b83",
X"e3a80cf1",
X"ec3f8151",
X"f6ba3f83",
X"3d0d04fc",
X"3d0d9080",
X"80528684",
X"808051d0",
X"bb3f83e0",
X"8008b838",
X"80e1b451",
X"d4fe3f83",
X"e0800883",
X"e3c00854",
X"80e0a053",
X"83e08008",
X"5255cfda",
X"3f83e080",
X"088438f8",
X"ab3f8180",
X"80548280",
X"805380e0",
X"9c527451",
X"f7f53f81",
X"51f5e53f",
X"feb73ffc",
X"3983e08c",
X"080283e0",
X"8c0cfb3d",
X"0d0280e0",
X"ac0b83e0",
X"a40c80e0",
X"b00b83e0",
X"9c0c80e0",
X"b40b83e0",
X"ac0c83e0",
X"8c08fc05",
X"0c800b83",
X"e3ac0b83",
X"e08c08f8",
X"050c83e0",
X"8c08f405",
X"0ccea93f",
X"83e08008",
X"8605fc06",
X"83e08c08",
X"f0050c02",
X"83e08c08",
X"f0050831",
X"0d833d70",
X"83e08c08",
X"f8050870",
X"840583e0",
X"8c08f805",
X"0c0c51ca",
X"f23f83e0",
X"8c08f405",
X"08810583",
X"e08c08f4",
X"050c83e0",
X"8c08f405",
X"08862e09",
X"8106ffad",
X"38869480",
X"8051edbf",
X"3fff0b83",
X"e3a80c80",
X"0b83e3c8",
X"0c84d8c0",
X"0b83e3c4",
X"0c8151f0",
X"f23f8151",
X"f1973f80",
X"51f1923f",
X"8151f1b8",
X"3f8151f2",
X"8d3f8251",
X"f1db3f80",
X"51f2b13f",
X"80c68a52",
X"8051c8b1",
X"3ffdcc3f",
X"83e08c08",
X"fc05080d",
X"800b83e0",
X"800c873d",
X"0d83e08c",
X"0c04fd3d",
X"0d755480",
X"740c800b",
X"84150c80",
X"0b88150c",
X"87d08933",
X"87d08f33",
X"70822a70",
X"81067030",
X"70720770",
X"09709f2c",
X"77069e06",
X"54515155",
X"51515353",
X"80729806",
X"52537088",
X"2e098106",
X"83388153",
X"70983270",
X"30708025",
X"75713184",
X"180c5151",
X"51807286",
X"06525370",
X"822e0981",
X"06833881",
X"53708632",
X"70307080",
X"25757131",
X"770c5151",
X"51719432",
X"70307080",
X"2588170c",
X"5151853d",
X"0d04fe3d",
X"0d747654",
X"527151fe",
X"ed3f7281",
X"2ea23881",
X"73268d38",
X"72822eab",
X"3872832e",
X"9f38e639",
X"7108e238",
X"841208dd",
X"38881208",
X"d838a039",
X"88120881",
X"2e098106",
X"cc389439",
X"88120881",
X"2e8d3871",
X"08893884",
X"1208802e",
X"ffb73884",
X"3d0d04ff",
X"3d0d7352",
X"7183e3d0",
X"082ea638",
X"71a00a07",
X"90809c0c",
X"90808c08",
X"5170802e",
X"f738800b",
X"90809c0c",
X"90808c08",
X"5170f938",
X"7183e3d0",
X"0c833d0d",
X"04ff0b83",
X"e3d00c81",
X"80800b83",
X"e3cc0c80",
X"0b83e080",
X"0c04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"9e3f7280",
X"2ea33883",
X"e3cc0814",
X"52713375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552da",
X"39800b83",
X"e0800c86",
X"3d0d04f7",
X"3d0d7b7d",
X"7f115855",
X"59805573",
X"762eb138",
X"83e3cc08",
X"8b3d5957",
X"74197033",
X"75fc0619",
X"70085d76",
X"83067b07",
X"53545451",
X"72713479",
X"720c8114",
X"81165654",
X"73762e09",
X"8106d938",
X"800b83e0",
X"800c8b3d",
X"0d04803d",
X"0d83e3d0",
X"08900a07",
X"90809c0c",
X"90808c08",
X"5170802e",
X"f738800b",
X"90809c0c",
X"90808c08",
X"5170f938",
X"823d0d04",
X"83e08c08",
X"0283e08c",
X"0cfd3d0d",
X"805383e0",
X"8c088c05",
X"085283e0",
X"8c088805",
X"085183d4",
X"3f83e080",
X"087083e0",
X"800c5485",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"fd3d0d81",
X"5383e08c",
X"088c0508",
X"5283e08c",
X"08880508",
X"5183a13f",
X"83e08008",
X"7083e080",
X"0c54853d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cf9",
X"3d0d800b",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"05088025",
X"b93883e0",
X"8c088805",
X"083083e0",
X"8c088805",
X"0c800b83",
X"e08c08f4",
X"050c83e0",
X"8c08fc05",
X"088a3881",
X"0b83e08c",
X"08f4050c",
X"83e08c08",
X"f4050883",
X"e08c08fc",
X"050c83e0",
X"8c088c05",
X"088025b9",
X"3883e08c",
X"088c0508",
X"3083e08c",
X"088c050c",
X"800b83e0",
X"8c08f005",
X"0c83e08c",
X"08fc0508",
X"8a38810b",
X"83e08c08",
X"f0050c83",
X"e08c08f0",
X"050883e0",
X"8c08fc05",
X"0c805383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"05085181",
X"df3f83e0",
X"80087083",
X"e08c08f8",
X"050c5483",
X"e08c08fc",
X"0508802e",
X"903883e0",
X"8c08f805",
X"083083e0",
X"8c08f805",
X"0c83e08c",
X"08f80508",
X"7083e080",
X"0c54893d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cfb",
X"3d0d800b",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"05088025",
X"993883e0",
X"8c088805",
X"083083e0",
X"8c088805",
X"0c810b83",
X"e08c08fc",
X"050c83e0",
X"8c088c05",
X"08802590",
X"3883e08c",
X"088c0508",
X"3083e08c",
X"088c050c",
X"815383e0",
X"8c088c05",
X"085283e0",
X"8c088805",
X"0851bd3f",
X"83e08008",
X"7083e08c",
X"08f8050c",
X"5483e08c",
X"08fc0508",
X"802e9038",
X"83e08c08",
X"f8050830",
X"83e08c08",
X"f8050c83",
X"e08c08f8",
X"05087083",
X"e0800c54",
X"873d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cfd3d0d",
X"810b83e0",
X"8c08fc05",
X"0c800b83",
X"e08c08f8",
X"050c83e0",
X"8c088c05",
X"0883e08c",
X"08880508",
X"27b93883",
X"e08c08fc",
X"0508802e",
X"ae38800b",
X"83e08c08",
X"8c050824",
X"a23883e0",
X"8c088c05",
X"081083e0",
X"8c088c05",
X"0c83e08c",
X"08fc0508",
X"1083e08c",
X"08fc050c",
X"ffb83983",
X"e08c08fc",
X"0508802e",
X"80e13883",
X"e08c088c",
X"050883e0",
X"8c088805",
X"0826ad38",
X"83e08c08",
X"88050883",
X"e08c088c",
X"05083183",
X"e08c0888",
X"050c83e0",
X"8c08f805",
X"0883e08c",
X"08fc0508",
X"0783e08c",
X"08f8050c",
X"83e08c08",
X"fc050881",
X"2a83e08c",
X"08fc050c",
X"83e08c08",
X"8c050881",
X"2a83e08c",
X"088c050c",
X"ff953983",
X"e08c0890",
X"0508802e",
X"933883e0",
X"8c088805",
X"087083e0",
X"8c08f405",
X"0c519139",
X"83e08c08",
X"f8050870",
X"83e08c08",
X"f4050c51",
X"83e08c08",
X"f4050883",
X"e0800c85",
X"3d0d83e0",
X"8c0c0483",
X"e08c0802",
X"83e08c0c",
X"ff3d0d80",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"88050881",
X"06ff1170",
X"097083e0",
X"8c088c05",
X"080683e0",
X"8c08fc05",
X"081183e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"812a83e0",
X"8c088805",
X"0c83e08c",
X"088c0508",
X"1083e08c",
X"088c050c",
X"51515151",
X"83e08c08",
X"88050880",
X"2e8438ff",
X"ab3983e0",
X"8c08fc05",
X"087083e0",
X"800c5183",
X"3d0d83e0",
X"8c0c04fc",
X"3d0d7670",
X"797b5555",
X"55558f72",
X"278c3872",
X"75078306",
X"5170802e",
X"a938ff12",
X"5271ff2e",
X"98387270",
X"81055433",
X"74708105",
X"5634ff12",
X"5271ff2e",
X"098106ea",
X"387483e0",
X"800c863d",
X"0d047451",
X"72708405",
X"54087170",
X"8405530c",
X"72708405",
X"54087170",
X"8405530c",
X"72708405",
X"54087170",
X"8405530c",
X"72708405",
X"54087170",
X"8405530c",
X"f0125271",
X"8f26c938",
X"83722795",
X"38727084",
X"05540871",
X"70840553",
X"0cfc1252",
X"718326ed",
X"387054ff",
X"81390000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"0000256e",
X"000025af",
X"000025d0",
X"000025f6",
X"000025f6",
X"000025f6",
X"000026b9",
X"25732025",
X"73000000",
X"20000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"31364b00",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"43617274",
X"72696467",
X"65203332",
X"6b000000",
X"43617274",
X"72696467",
X"65203136",
X"6b206f6e",
X"65206368",
X"69700000",
X"43617274",
X"72696467",
X"65203136",
X"6b207477",
X"6f206368",
X"69700000",
X"45786974",
X"00000000",
X"61636964",
X"35323030",
X"2e726f6d",
X"00000000",
X"524f4d00",
X"42494e00",
X"43415200",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
