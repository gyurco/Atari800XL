
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81e0",
X"8c738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81e9",
X"980c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757581da",
X"bb2d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7581d8cf",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80e89804",
X"fd3d0d75",
X"705254ae",
X"c33f83c0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"c0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83c0",
X"8008732e",
X"a13883c0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183c0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83c2d808",
X"248a38b5",
X"983fff0b",
X"83c2d80c",
X"800b83c0",
X"800c04ff",
X"3d0d7352",
X"83c0b408",
X"722e9b38",
X"d93f8183",
X"0b9088a0",
X"0c715196",
X"c93f8193",
X"0b9088a0",
X"0c7183c0",
X"b40c833d",
X"0d04f43d",
X"0d7e6062",
X"5c5a5580",
X"568154bc",
X"1508762e",
X"09810681",
X"92387451",
X"ffb93f79",
X"58757a25",
X"80f73883",
X"c3880870",
X"892a5783",
X"ff067884",
X"80723156",
X"56577378",
X"25833873",
X"557583c2",
X"d8082e84",
X"38fef33f",
X"83c2d808",
X"8025a638",
X"75892b51",
X"98fd3f83",
X"c388088f",
X"3dfc1155",
X"5c548152",
X"f81b5196",
X"e73f7614",
X"83c3880c",
X"7583c2d8",
X"0c745376",
X"527851b3",
X"b33f83c0",
X"800883c3",
X"88081683",
X"c3880c78",
X"7631761b",
X"5b595677",
X"8024ff8b",
X"38617a71",
X"0c547554",
X"75802e83",
X"38815473",
X"83c0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"853f7651",
X"fe993f86",
X"3dfc0553",
X"78527751",
X"968a3f79",
X"75710c54",
X"83c08008",
X"5483c080",
X"08802e83",
X"38815473",
X"83c0800c",
X"863d0d04",
X"fe3d0d75",
X"83c2d808",
X"53538072",
X"24953871",
X"732e9038",
X"80c30b90",
X"88a00c71",
X"9088a40c",
X"fdb43f80",
X"d30b9088",
X"a00c7451",
X"fdc13f80",
X"e30b9088",
X"a00c7251",
X"97b53f80",
X"f30b9088",
X"a00c83c0",
X"80085283",
X"c0800880",
X"2e833881",
X"527183c0",
X"800c843d",
X"0d04803d",
X"0d7280c0",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"3d0d72bc",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"c40b83c0",
X"800c04fd",
X"3d0d7577",
X"71547053",
X"5553a9e4",
X"3f82c813",
X"08bc150c",
X"82c01308",
X"80c0150c",
X"fcb43f73",
X"5193ab3f",
X"7383c0b4",
X"0c83c080",
X"085383c0",
X"8008802e",
X"83388153",
X"7283c080",
X"0c853d0d",
X"04fd3d0d",
X"75775553",
X"fc883f72",
X"802ea538",
X"bc130852",
X"7351a8ee",
X"3f83c080",
X"088f3877",
X"527251ff",
X"9a3f83c0",
X"8008538a",
X"3982cc13",
X"0853d839",
X"81537283",
X"c0800c85",
X"3d0d04fe",
X"3d0dff0b",
X"83c2d80c",
X"7483c0b8",
X"0c7583c2",
X"d40cafc6",
X"3f83c080",
X"0881ff06",
X"52815371",
X"993883c2",
X"f0518e94",
X"3f83c080",
X"085283c0",
X"8008802e",
X"83387252",
X"71537283",
X"c0800c84",
X"3d0d04fa",
X"3d0d787a",
X"82c41208",
X"82c41208",
X"70722459",
X"56565757",
X"73732e09",
X"81069138",
X"80c01652",
X"80c01751",
X"a6df3f83",
X"c0800855",
X"7483c080",
X"0c883d0d",
X"04f63d0d",
X"7c5b807b",
X"715c5457",
X"7a772e8c",
X"38811a82",
X"cc140854",
X"5a72f638",
X"805980d9",
X"397a5481",
X"5780707b",
X"7b315a57",
X"55ff1853",
X"74732580",
X"c13882cc",
X"14085273",
X"51ff8c3f",
X"800b83c0",
X"800825a1",
X"3882cc14",
X"0882cc11",
X"0882cc16",
X"0c7482cc",
X"120c5375",
X"802e8638",
X"7282cc17",
X"0c725480",
X"577382cc",
X"15088117",
X"575556ff",
X"b8398119",
X"59800bff",
X"1b545478",
X"73258338",
X"81547681",
X"32707506",
X"515372ff",
X"90388c3d",
X"0d04f73d",
X"0d7b7d5a",
X"5a82d052",
X"83c2d408",
X"5181c6d5",
X"3f83c080",
X"0857f9aa",
X"3f795283",
X"c2dc5195",
X"b73f83c0",
X"80085480",
X"5383c080",
X"08732e09",
X"81068283",
X"3883c0b8",
X"080b0b81",
X"e5e05370",
X"5256a69c",
X"3f0b0b81",
X"e5e05280",
X"c01651a6",
X"8f3f75bc",
X"170c7382",
X"c0170c81",
X"0b82c417",
X"0c810b82",
X"c8170c73",
X"82cc170c",
X"ff1782d0",
X"17555781",
X"913983c0",
X"c4337082",
X"2a708106",
X"51545572",
X"81803874",
X"812a8106",
X"587780f6",
X"3874842a",
X"810682c4",
X"150c83c0",
X"c4338106",
X"82c8150c",
X"79527351",
X"a5b63f73",
X"51a5cd3f",
X"83c08008",
X"1453af73",
X"70810555",
X"3472bc15",
X"0c83c0c5",
X"527251a5",
X"973f83c0",
X"bc0882c0",
X"150c83c0",
X"d25280c0",
X"1451a584",
X"3f78802e",
X"8d387351",
X"782d83c0",
X"8008802e",
X"99387782",
X"cc150c75",
X"802e8638",
X"7382cc17",
X"0c7382d0",
X"15ff1959",
X"55567680",
X"2e9b3883",
X"c0bc5283",
X"c2dc5194",
X"ad3f83c0",
X"80088a38",
X"83c0c533",
X"5372fed2",
X"3878802e",
X"893883c0",
X"b80851fc",
X"b83f83c0",
X"b8085372",
X"83c0800c",
X"8b3d0d04",
X"ff3d0d80",
X"527351fd",
X"b53f833d",
X"0d04f03d",
X"0d627052",
X"54f5d93f",
X"83c08008",
X"7453873d",
X"70535555",
X"f5f93ff6",
X"d93f7351",
X"d33f6353",
X"745283c0",
X"800851fa",
X"b83f923d",
X"0d047183",
X"c0800c04",
X"80c01283",
X"c0800c04",
X"803d0d72",
X"82c01108",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"7282cc11",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d7282c4",
X"110883c0",
X"800c5182",
X"3d0d04f9",
X"3d0d7983",
X"c0900857",
X"57817727",
X"81963876",
X"88170827",
X"818e3875",
X"33557482",
X"2e893874",
X"832eb338",
X"80fe3974",
X"54761083",
X"fe065376",
X"882a8c17",
X"08055289",
X"3dfc0551",
X"a9f43f83",
X"c0800880",
X"df38029d",
X"0533893d",
X"3371882b",
X"07565680",
X"d1398454",
X"76822b83",
X"fc065376",
X"872a8c17",
X"08055289",
X"3dfc0551",
X"a9c43f83",
X"c08008b0",
X"38029f05",
X"33028405",
X"9e053371",
X"982b7190",
X"2b07028c",
X"059d0533",
X"70882b72",
X"078d3d33",
X"7180ffff",
X"fe800607",
X"51525357",
X"58568339",
X"81557483",
X"c0800c89",
X"3d0d04fb",
X"3d0d83c0",
X"9008fe19",
X"881208fe",
X"05555654",
X"80567473",
X"278d3882",
X"14337571",
X"29941608",
X"05575375",
X"83c0800c",
X"873d0d04",
X"fc3d0d76",
X"52800b83",
X"c0900870",
X"33515253",
X"70832e09",
X"81069138",
X"95123394",
X"13337198",
X"2b71902b",
X"07555551",
X"9b12339a",
X"13337188",
X"2b077407",
X"83c0800c",
X"55863d0d",
X"04fc3d0d",
X"7683c090",
X"08555580",
X"75238815",
X"08537281",
X"2e883888",
X"14087326",
X"85388152",
X"b2397290",
X"38733352",
X"71832e09",
X"81068538",
X"90140853",
X"728c160c",
X"72802e8d",
X"387251fe",
X"d63f83c0",
X"80085285",
X"39901408",
X"52719016",
X"0c805271",
X"83c0800c",
X"863d0d04",
X"fa3d0d78",
X"83c09008",
X"71228105",
X"7083ffff",
X"06575457",
X"5573802e",
X"88389015",
X"08537286",
X"38835280",
X"e739738f",
X"06527180",
X"da388113",
X"90160c8c",
X"15085372",
X"9038830b",
X"84172257",
X"52737627",
X"80c638bf",
X"39821633",
X"ff057484",
X"2a065271",
X"b2387251",
X"fcb13f81",
X"527183c0",
X"800827a8",
X"38835283",
X"c0800888",
X"1708279c",
X"3883c080",
X"088c160c",
X"83c08008",
X"51fdbc3f",
X"83c08008",
X"90160c73",
X"75238052",
X"7183c080",
X"0c883d0d",
X"04f23d0d",
X"60626458",
X"5e5b7533",
X"5574a02e",
X"09810688",
X"38811670",
X"4456ef39",
X"62703356",
X"5674af2e",
X"09810684",
X"38811643",
X"800b881c",
X"0c627033",
X"5155749f",
X"2691387a",
X"51fdd23f",
X"83c08008",
X"56807d34",
X"83813993",
X"3d841c08",
X"7058595f",
X"8a55a076",
X"70810558",
X"34ff1555",
X"74ff2e09",
X"8106ef38",
X"80705a5c",
X"887f085f",
X"5a7b811d",
X"7081ff06",
X"60137033",
X"70af3270",
X"30a07327",
X"71802507",
X"5151525b",
X"535e5755",
X"7480e738",
X"76ae2e09",
X"81068338",
X"8155787a",
X"27750755",
X"74802e9f",
X"38798832",
X"703078ae",
X"32703070",
X"73079f2a",
X"53515751",
X"5675bb38",
X"88598b5a",
X"ffab3976",
X"982b5574",
X"80258738",
X"81df9c17",
X"3357ff9f",
X"17557499",
X"268938e0",
X"177081ff",
X"06585578",
X"811a7081",
X"ff06721b",
X"535b5755",
X"767534fe",
X"f8397b1e",
X"7f0c8055",
X"76a02683",
X"38815574",
X"8b19347a",
X"51fc823f",
X"83c08008",
X"80f538a0",
X"547a2270",
X"852b83e0",
X"06545590",
X"1b08527c",
X"51a3ff3f",
X"83c08008",
X"5783c080",
X"08818138",
X"7c335574",
X"802e80f4",
X"388b1d33",
X"70832a70",
X"81065156",
X"5674b438",
X"8b7d841d",
X"0883c080",
X"08595b5b",
X"58ff1858",
X"77ff2e9a",
X"38797081",
X"055b3379",
X"7081055b",
X"33717131",
X"52565675",
X"802ee238",
X"86397580",
X"2e96387a",
X"51fbe53f",
X"ff863983",
X"c0800856",
X"83c08008",
X"b6388339",
X"7656841b",
X"088b1133",
X"515574a7",
X"388b1d33",
X"70842a70",
X"81065156",
X"56748938",
X"83569439",
X"81569039",
X"7c51fa94",
X"3f83c080",
X"08881c0c",
X"fd813975",
X"83c0800c",
X"903d0d04",
X"f83d0d7a",
X"7c595782",
X"5483fe53",
X"77527651",
X"a2c43f83",
X"5683c080",
X"0880ec38",
X"81173377",
X"3371882b",
X"07565682",
X"567482d4",
X"d52e0981",
X"0680d438",
X"7554b653",
X"77527651",
X"a2983f83",
X"c0800898",
X"38811733",
X"77337188",
X"2b0783c0",
X"80085256",
X"56748182",
X"c62eac38",
X"825480d2",
X"53775276",
X"51a1ef3f",
X"83c08008",
X"98388117",
X"33773371",
X"882b0783",
X"c0800852",
X"56567481",
X"82c62e83",
X"38815675",
X"83c0800c",
X"8a3d0d04",
X"eb3d0d67",
X"5a800b83",
X"c0900ca1",
X"913f83c0",
X"80088106",
X"55825674",
X"83ef3874",
X"75538f3d",
X"70535759",
X"feca3f83",
X"c0800881",
X"ff065776",
X"812e0981",
X"0680d438",
X"905483be",
X"53745275",
X"51a1833f",
X"83c08008",
X"80c9388f",
X"3d335574",
X"802e80c9",
X"3802bf05",
X"33028405",
X"be053371",
X"982b7190",
X"2b07028c",
X"05bd0533",
X"70882b72",
X"07953d33",
X"71077058",
X"7b575e52",
X"5e575957",
X"fdee3f83",
X"c0800881",
X"ff065776",
X"832e0981",
X"06863881",
X"5682f239",
X"76802e86",
X"38865682",
X"e839a454",
X"8d537852",
X"7551a09a",
X"3f815683",
X"c0800882",
X"d43802be",
X"05330284",
X"05bd0533",
X"71882b07",
X"595d77ab",
X"380280ce",
X"05330284",
X"0580cd05",
X"3371982b",
X"71902b07",
X"973d3370",
X"882b7207",
X"02940580",
X"cb053371",
X"0754525e",
X"57595602",
X"b7053378",
X"71290288",
X"05b60533",
X"028c05b5",
X"05337188",
X"2b07701d",
X"707f8c05",
X"0c5f5957",
X"595d8e3d",
X"33821b34",
X"02b90533",
X"903d3371",
X"882b075a",
X"5c78841b",
X"2302bb05",
X"33028405",
X"ba053371",
X"882b0756",
X"5c74ab38",
X"0280ca05",
X"33028405",
X"80c90533",
X"71982b71",
X"902b0796",
X"3d337088",
X"2b720702",
X"940580c7",
X"05337107",
X"51525357",
X"5e5c7476",
X"31783179",
X"842a903d",
X"33547171",
X"31535656",
X"81b7ba3f",
X"83c08008",
X"82057088",
X"1c0c83c0",
X"8008e08a",
X"05565674",
X"83dffe26",
X"83388257",
X"83fff676",
X"27853883",
X"57893986",
X"5676802e",
X"80db3876",
X"7a347683",
X"2e098106",
X"b0380280",
X"d6053302",
X"840580d5",
X"05337198",
X"2b71902b",
X"07993d33",
X"70882b72",
X"07029405",
X"80d30533",
X"71077f90",
X"050c525e",
X"57585686",
X"39771b90",
X"1b0c841a",
X"228c1b08",
X"1971842a",
X"05941c0c",
X"5d800b81",
X"1b347983",
X"c0900c80",
X"567583c0",
X"800c973d",
X"0d04e93d",
X"0d83c090",
X"08568554",
X"75802e81",
X"8238800b",
X"81173499",
X"3de01146",
X"6a548a3d",
X"705458ec",
X"0551f6e5",
X"3f83c080",
X"085483c0",
X"800880df",
X"38893d33",
X"5473802e",
X"913802ab",
X"05337084",
X"2a810651",
X"5574802e",
X"86388354",
X"80c13976",
X"51f4893f",
X"83c08008",
X"a0170c02",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"9c1c0c52",
X"78981b0c",
X"53565957",
X"810b8117",
X"34745473",
X"83c0800c",
X"993d0d04",
X"f53d0d7d",
X"7f617283",
X"c090085a",
X"5d5d595c",
X"807b0c85",
X"5775802e",
X"81e03881",
X"16338106",
X"55845774",
X"802e81d2",
X"38913974",
X"81173486",
X"39800b81",
X"17348157",
X"81c0399c",
X"16089817",
X"08315574",
X"78278338",
X"74587780",
X"2e81a938",
X"98160870",
X"83ff0656",
X"577480cf",
X"38821633",
X"ff057789",
X"2a067081",
X"ff065a55",
X"78a03876",
X"8738a016",
X"08558d39",
X"a4160851",
X"f0e93f83",
X"c0800855",
X"817527ff",
X"a83874a4",
X"170ca416",
X"0851f283",
X"3f83c080",
X"085583c0",
X"8008802e",
X"ff893883",
X"c0800819",
X"a8170c98",
X"160883ff",
X"06848071",
X"31515577",
X"75278338",
X"77557483",
X"ffff0654",
X"98160883",
X"ff0653a8",
X"16085279",
X"577b8338",
X"7b577651",
X"9ac03f83",
X"c08008fe",
X"d0389816",
X"08159817",
X"0c741a78",
X"76317c08",
X"177d0c59",
X"5afed339",
X"80577683",
X"c0800c8d",
X"3d0d04fa",
X"3d0d7883",
X"c0900855",
X"56855573",
X"802e81e3",
X"38811433",
X"81065384",
X"5572802e",
X"81d5389c",
X"14085372",
X"76278338",
X"72569814",
X"0857800b",
X"98150c75",
X"802e81b9",
X"38821433",
X"70892b56",
X"5376802e",
X"b7387452",
X"ff165181",
X"b2bb3f83",
X"c08008ff",
X"18765470",
X"53585381",
X"b2ab3f83",
X"c0800873",
X"26963874",
X"30707806",
X"7098170c",
X"777131a4",
X"17085258",
X"51538939",
X"a0140870",
X"a4160c53",
X"747627b9",
X"387251ee",
X"d63f83c0",
X"80085381",
X"0b83c080",
X"08278b38",
X"88140883",
X"c0800826",
X"8838800b",
X"811534b0",
X"3983c080",
X"08a4150c",
X"98140815",
X"98150c75",
X"753156c4",
X"39981408",
X"16709816",
X"0c735256",
X"efc53f83",
X"c080088c",
X"3883c080",
X"08811534",
X"81559439",
X"821433ff",
X"0576892a",
X"0683c080",
X"0805a815",
X"0c805574",
X"83c0800c",
X"883d0d04",
X"ef3d0d63",
X"56855583",
X"c0900880",
X"2e80d238",
X"933df405",
X"84170c64",
X"53883d70",
X"53765257",
X"f1cf3f83",
X"c0800855",
X"83c08008",
X"b438883d",
X"33547380",
X"2ea13802",
X"a7053370",
X"842a7081",
X"06515555",
X"83557380",
X"2e973876",
X"51eef53f",
X"83c08008",
X"88170c75",
X"51efa63f",
X"83c08008",
X"557483c0",
X"800c933d",
X"0d04e43d",
X"0d6ea13d",
X"08405e85",
X"5683c090",
X"08802e84",
X"85389e3d",
X"f405841f",
X"0c7e9838",
X"7d51eef5",
X"3f83c080",
X"085683ee",
X"39814181",
X"f6398341",
X"81f13993",
X"3d7f9605",
X"4159807f",
X"8295055e",
X"56756081",
X"ff053483",
X"41901e08",
X"762e81d3",
X"38a0547d",
X"2270852b",
X"83e00654",
X"58901e08",
X"52785196",
X"c93f83c0",
X"80084183",
X"c08008ff",
X"b8387833",
X"5c7b802e",
X"ffb4388b",
X"193370bf",
X"06718106",
X"52435574",
X"802e80de",
X"387b81bf",
X"0655748f",
X"2480d338",
X"9a193355",
X"7480cb38",
X"f31d7058",
X"5d815675",
X"8b2e0981",
X"0685388e",
X"568b3975",
X"9a2e0981",
X"0683389c",
X"56751970",
X"70810552",
X"33713381",
X"1a821a5f",
X"5b525b55",
X"74863879",
X"77348539",
X"80df7734",
X"777b5757",
X"7aa02e09",
X"8106c038",
X"81567b81",
X"e5327030",
X"709f2a51",
X"51557bae",
X"2e933874",
X"802e8e38",
X"61832a70",
X"81065155",
X"74802e97",
X"387d51ed",
X"df3f83c0",
X"80084183",
X"c0800887",
X"38901e08",
X"feaf3880",
X"60347580",
X"2e88387c",
X"527f518d",
X"eb3f6080",
X"2e863880",
X"0b901f0c",
X"60566083",
X"2e853860",
X"81d03889",
X"1f57901e",
X"08802e81",
X"a8388056",
X"75197033",
X"515574a0",
X"2ea03874",
X"852e0981",
X"06843881",
X"e5557477",
X"70810559",
X"34811670",
X"81ff0657",
X"55877627",
X"d7388819",
X"335574a0",
X"2ea938ae",
X"77708105",
X"59348856",
X"75197033",
X"515574a0",
X"2e953874",
X"77708105",
X"59348116",
X"7081ff06",
X"57558a76",
X"27e2388b",
X"19337f88",
X"05349f19",
X"339e1a33",
X"71982b71",
X"902b079d",
X"1c337088",
X"2b72079c",
X"1e337107",
X"640c5299",
X"1d33981e",
X"3371882b",
X"07535153",
X"57595674",
X"7f840523",
X"97193396",
X"1a337188",
X"2b075656",
X"747f8605",
X"23807734",
X"7d51ebf0",
X"3f83c080",
X"08833270",
X"30707207",
X"9f2c83c0",
X"80080652",
X"5656961f",
X"3355748a",
X"38891f52",
X"961f518b",
X"f73f7583",
X"c0800c9e",
X"3d0d04f4",
X"3d0d7e8f",
X"3dec1156",
X"56589053",
X"f0155277",
X"51e0b13f",
X"83c08008",
X"80d63878",
X"902e0981",
X"0680cd38",
X"02ab0533",
X"81e9a00b",
X"81e9a033",
X"5758568c",
X"3974762e",
X"8a388417",
X"70335657",
X"74f33876",
X"33705755",
X"74802eac",
X"38821722",
X"708a2b90",
X"3dec0556",
X"70555656",
X"96800a52",
X"7751dfe0",
X"3f83c080",
X"08863878",
X"752e8538",
X"80568539",
X"81173356",
X"7583c080",
X"0c8e3d0d",
X"04fc3d0d",
X"76705255",
X"8afe3f83",
X"c0800815",
X"ff055473",
X"752e8e38",
X"73335372",
X"ae2e8638",
X"ff1454ef",
X"39775281",
X"14518a96",
X"3f83c080",
X"08307083",
X"c0800807",
X"802583c0",
X"800c5386",
X"3d0d04fa",
X"3d0d7857",
X"80775256",
X"e6c23f83",
X"c0800883",
X"c0800833",
X"53547176",
X"2e80c738",
X"733383c0",
X"94173356",
X"53749138",
X"765183c3",
X"ac085271",
X"2d83c080",
X"0852ad39",
X"ff9f1352",
X"71992689",
X"38e01370",
X"81ff0654",
X"52747332",
X"70307072",
X"07802578",
X"05811770",
X"33545758",
X"545271ff",
X"bb388052",
X"7183c080",
X"0c883d0d",
X"04fc3d0d",
X"76705255",
X"e6803f83",
X"c0800854",
X"815383c0",
X"800880d0",
X"387451e5",
X"c33f83c0",
X"800881e5",
X"f05383c0",
X"80085253",
X"fea33f83",
X"c08008b0",
X"3881e5f4",
X"527251fe",
X"943f83c0",
X"8008a138",
X"81e5f852",
X"7251fe85",
X"3f83c080",
X"08923881",
X"e5fc5272",
X"51fdf63f",
X"83c08008",
X"802e8338",
X"81547353",
X"7283c080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"e5903f81",
X"5383c080",
X"08983873",
X"51e4d93f",
X"83c3a008",
X"5283c080",
X"0851fdbd",
X"3f83c080",
X"08537283",
X"c0800c85",
X"3d0d04dd",
X"3d0da63d",
X"085f800b",
X"83c7e033",
X"555b737b",
X"2e85cc38",
X"86537a52",
X"83c09451",
X"a1c73f7e",
X"51daae3f",
X"83c08008",
X"33973d56",
X"54737b2e",
X"09810696",
X"3881eae0",
X"52745187",
X"db3f9a39",
X"7e527851",
X"dde13f85",
X"96397e51",
X"da8f3f83",
X"c0800852",
X"7451d9bf",
X"3f804480",
X"43804280",
X"41adbb52",
X"963d7052",
X"5ee0cb3f",
X"83c08008",
X"59800b83",
X"c0800855",
X"5c83c080",
X"087c2e94",
X"38811c74",
X"525ce3cd",
X"3f83c080",
X"085483c0",
X"8008ee38",
X"805aff40",
X"7909709f",
X"2c7b065b",
X"547b7a24",
X"8438ff1c",
X"5af61a70",
X"09709f2c",
X"72067bff",
X"125a5a52",
X"55558075",
X"25953876",
X"51e3923f",
X"83c08008",
X"76ff1858",
X"55577380",
X"24ed3874",
X"602e8638",
X"a2823f74",
X"4078ff1b",
X"70585e58",
X"807a2595",
X"387751e2",
X"e83f83c0",
X"800876ff",
X"18585558",
X"738024ed",
X"38800b83",
X"c7dc0c81",
X"800b83c8",
X"a80c81e6",
X"80518bdf",
X"3f800b83",
X"c8a80c83",
X"c0945281",
X"e688518b",
X"ce3fa80b",
X"83c7dc0c",
X"76802e80",
X"e43883c7",
X"dc087779",
X"32703070",
X"72078025",
X"70872b83",
X"c8a80c51",
X"56785356",
X"56e29b3f",
X"83c08008",
X"802e8838",
X"81e69451",
X"8b953f76",
X"51e1dd3f",
X"83c08008",
X"5281e8c0",
X"518b843f",
X"7651e1e5",
X"3f83c080",
X"0883c7dc",
X"08555775",
X"74258638",
X"a81656f7",
X"397583c7",
X"dc0c86f0",
X"7624ff98",
X"3887980b",
X"83c7dc0c",
X"77802ea9",
X"387751e1",
X"9b3f83c0",
X"80087852",
X"55e1bb3f",
X"81e69c54",
X"83c08008",
X"853881e6",
X"98547453",
X"735281e5",
X"e4518aab",
X"3f805481",
X"e5ec518a",
X"a23f8114",
X"5473a82e",
X"098106ef",
X"38868da0",
X"519e803f",
X"8052913d",
X"705257ba",
X"ad3f8352",
X"7651baa6",
X"3f645473",
X"ff2e0981",
X"069738ff",
X"1b700970",
X"9f2c7206",
X"52555b80",
X"0b83c094",
X"1c3481c2",
X"39807425",
X"ab387a85",
X"2e098106",
X"91388653",
X"805283c0",
X"94519dbd",
X"3f805b81",
X"a5397383",
X"c0941c34",
X"811b5b81",
X"99398076",
X"34819339",
X"63818f38",
X"62802e80",
X"fb387c54",
X"73ff2e96",
X"3878802e",
X"81893878",
X"51dffa3f",
X"83c08008",
X"ff155559",
X"e7397880",
X"2e80f438",
X"7851dff6",
X"3f83c080",
X"08802efb",
X"c7387851",
X"dfbe3f83",
X"c0800852",
X"81e5e051",
X"81e73f83",
X"c08008a3",
X"387d5183",
X"9f3f83c0",
X"80085574",
X"ff165654",
X"807425ae",
X"38741e70",
X"33555673",
X"af2eff8a",
X"38e93978",
X"51deff3f",
X"83c08008",
X"527d5182",
X"d73f8f39",
X"60882961",
X"10057a05",
X"62055afb",
X"c7396380",
X"2efb8a38",
X"80527651",
X"b8b83fa5",
X"3d0d04ff",
X"3d0d028f",
X"05337010",
X"81059088",
X"900c5283",
X"3d0d04ff",
X"3d0d028f",
X"05335290",
X"88840870",
X"892a7081",
X"06515151",
X"70802e86",
X"38afca3f",
X"ea397190",
X"88800c83",
X"3d0d0480",
X"3d0d9088",
X"8c087088",
X"2a708106",
X"51515170",
X"802e8638",
X"afa73fea",
X"39908888",
X"0883c080",
X"0c823d0d",
X"04908894",
X"0883c080",
X"0c04fd3d",
X"0d757754",
X"54807325",
X"94387370",
X"81055533",
X"5281e6a0",
X"5187883f",
X"ff1353e9",
X"39853d0d",
X"04fd3d0d",
X"75775354",
X"73335170",
X"89387133",
X"5170802e",
X"a1387333",
X"72335253",
X"72712785",
X"38ff5194",
X"39707327",
X"85388151",
X"8b398114",
X"81135354",
X"d3398051",
X"7083c080",
X"0c853d0d",
X"04fd3d0d",
X"75775454",
X"72337081",
X"ff065252",
X"70802ea3",
X"387181ff",
X"068114ff",
X"bf125354",
X"52709926",
X"8938a012",
X"7081ff06",
X"53517174",
X"70810556",
X"34d23980",
X"7434853d",
X"0d04ffbd",
X"3d0d80c6",
X"3d0852a5",
X"3d705254",
X"ffb33f80",
X"c73d0852",
X"853d7052",
X"53ffa63f",
X"72527351",
X"fedf3f80",
X"c53d0d04",
X"fe3d0d74",
X"76535371",
X"70810553",
X"33517073",
X"70810555",
X"3470f038",
X"843d0d04",
X"fe3d0d74",
X"52807233",
X"52537073",
X"2e8d3881",
X"12811471",
X"33535452",
X"70f53872",
X"83c0800c",
X"843d0d04",
X"f63d0d7c",
X"7e60625a",
X"5d5b5680",
X"59815585",
X"39747a29",
X"55745275",
X"51819fa9",
X"3f83c080",
X"087a27ed",
X"3874802e",
X"80e03874",
X"52755181",
X"9f933f83",
X"c0800875",
X"53765254",
X"819fb93f",
X"83c08008",
X"7a537552",
X"56819ef9",
X"3f83c080",
X"08793070",
X"7b079f2a",
X"70778024",
X"07515154",
X"55728738",
X"83c08008",
X"c2387681",
X"18b01655",
X"58588974",
X"258b38b7",
X"14537a85",
X"3880d714",
X"53727834",
X"811959ff",
X"9c398077",
X"348c3d0d",
X"04f73d0d",
X"7b7d7f62",
X"029005bb",
X"05335759",
X"565a5ab0",
X"58728338",
X"a0587570",
X"70810552",
X"33715954",
X"55903980",
X"74258e38",
X"ff147770",
X"81055933",
X"545472ef",
X"3873ff15",
X"55538073",
X"25893877",
X"52795178",
X"2def3975",
X"33755753",
X"72802e90",
X"38725279",
X"51782d75",
X"70810557",
X"3353ed39",
X"8b3d0d04",
X"ee3d0d64",
X"66696970",
X"70810552",
X"335b4a5c",
X"5e5e7680",
X"2e82f938",
X"76a52e09",
X"810682e0",
X"38807041",
X"67707081",
X"05523371",
X"4a59575f",
X"76b02e09",
X"81068c38",
X"75708105",
X"57337648",
X"57815fd0",
X"17567589",
X"2680da38",
X"76675c59",
X"805c9339",
X"778a2480",
X"c3387b8a",
X"29187b70",
X"81055d33",
X"5a5cd019",
X"7081ff06",
X"58588977",
X"27a438ff",
X"9f197081",
X"ff06ffa9",
X"1b5a5156",
X"85762792",
X"38ffbf19",
X"7081ff06",
X"51567585",
X"268a38c9",
X"19587780",
X"25ffb938",
X"7a477b40",
X"7881ff06",
X"577680e4",
X"2e80e538",
X"7680e424",
X"a7387680",
X"d82e8186",
X"387680d8",
X"24903876",
X"802e81cc",
X"3876a52e",
X"81b63881",
X"b9397680",
X"e32e818c",
X"3881af39",
X"7680f52e",
X"9b387680",
X"f5248b38",
X"7680f32e",
X"81813881",
X"99397680",
X"f82e80ca",
X"38818f39",
X"913d7055",
X"5780538a",
X"5279841b",
X"7108535b",
X"56fbfd3f",
X"7655ab39",
X"79841b71",
X"08943d70",
X"5b5b525b",
X"56758025",
X"8c387530",
X"56ad7834",
X"0280c105",
X"57765480",
X"538a5275",
X"51fbd13f",
X"77557e54",
X"b839913d",
X"70557780",
X"d8327030",
X"70802556",
X"51585690",
X"5279841b",
X"7108535b",
X"57fbad3f",
X"7555db39",
X"79841b83",
X"1233545b",
X"56983979",
X"841b7108",
X"575b5680",
X"547f537c",
X"527d51fc",
X"9c3f8739",
X"76527d51",
X"7c2d6670",
X"33588105",
X"47fd8339",
X"943d0d04",
X"7283c09c",
X"0c7183c0",
X"a00c04fb",
X"3d0d883d",
X"70708405",
X"52085754",
X"755383c0",
X"9c085283",
X"c0a00851",
X"fcc63f87",
X"3d0d04ff",
X"3d0d7370",
X"08535102",
X"93053372",
X"34700881",
X"05710c83",
X"3d0d04fc",
X"3d0d873d",
X"88115578",
X"54bddb53",
X"51fc993f",
X"8052873d",
X"51d13f86",
X"3d0d04fc",
X"3d0d7655",
X"7483c3b8",
X"082eaf38",
X"80537451",
X"87cc3f83",
X"c0800881",
X"ff06ff14",
X"7081ff06",
X"7230709f",
X"2a515255",
X"53547280",
X"2e843871",
X"dd3873fe",
X"387483c3",
X"b80c863d",
X"0d04ff3d",
X"0dff0b83",
X"c3b80c84",
X"b43f8151",
X"87903f83",
X"c0800881",
X"ff065271",
X"ee3881d4",
X"3f7183c0",
X"800c833d",
X"0d04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"823f7280",
X"2ea03883",
X"c3cc1433",
X"75708105",
X"57348114",
X"7083ffff",
X"06ff1570",
X"83ffff06",
X"56525552",
X"dd39800b",
X"83c0800c",
X"863d0d04",
X"fc3d0d76",
X"787a1156",
X"53558053",
X"71742e93",
X"38721551",
X"703383c3",
X"cc133481",
X"12811454",
X"52ea3980",
X"0b83c080",
X"0c863d0d",
X"04fd3d0d",
X"905483c3",
X"b8085186",
X"fd3f83c0",
X"800881ff",
X"06ff1571",
X"30713070",
X"73079f2a",
X"729f2a06",
X"52555255",
X"5372db38",
X"853d0d04",
X"803d0d83",
X"c3c40883",
X"2b83c3c0",
X"08079080",
X"a80c823d",
X"0d04800b",
X"83c3c40c",
X"e33f0481",
X"0b83c3c4",
X"0cda3f04",
X"ed3f0471",
X"83c3bc0c",
X"04803d0d",
X"8051f43f",
X"810b83c3",
X"c40c860b",
X"83c3c00c",
X"ffba3f82",
X"3d0d0484",
X"0b83c3c0",
X"0cffad3f",
X"04860b83",
X"c3c00cff",
X"a33f0483",
X"0b83c3c0",
X"0cff993f",
X"04870b83",
X"c3c00cff",
X"8f3f0480",
X"3d0d028b",
X"05339080",
X"a40c9080",
X"a8087081",
X"06515170",
X"f5389080",
X"a4087081",
X"ff0683c0",
X"800c5182",
X"3d0d0480",
X"3d0d81ff",
X"51d13f83",
X"c0800881",
X"ff0683c0",
X"800c823d",
X"0d04803d",
X"0d73902b",
X"73079080",
X"b40c823d",
X"0d0404fb",
X"3d0d7802",
X"84059f05",
X"3370982b",
X"55575572",
X"80259b38",
X"7580ff06",
X"56805280",
X"f751e03f",
X"83c08008",
X"81ff0654",
X"73812680",
X"fb38fee1",
X"3fffa43f",
X"fed13fff",
X"9e3f7551",
X"fef13f74",
X"982a51fe",
X"ea3f7490",
X"2a7081ff",
X"065253fe",
X"de3f7488",
X"2a7081ff",
X"065253fe",
X"d23f7481",
X"ff0651fe",
X"ca3f8155",
X"7580c02e",
X"09810686",
X"38819555",
X"8d397580",
X"c82e0981",
X"06843881",
X"87557451",
X"fea93f8a",
X"55fecc3f",
X"83c08008",
X"81ff0670",
X"982b5454",
X"7280258c",
X"38ff1570",
X"81ff0656",
X"5374e238",
X"7383c080",
X"0c873d0d",
X"04fa3d0d",
X"fdb73ffd",
X"d83f8a54",
X"fe993fff",
X"147081ff",
X"06555373",
X"f3387374",
X"535580c0",
X"51feac3f",
X"83c08008",
X"81ff0654",
X"73812e09",
X"8106829f",
X"3883aa52",
X"80c851fe",
X"923f83c0",
X"800881ff",
X"06537281",
X"2e098106",
X"81a83874",
X"54873d74",
X"115456fd",
X"ce3f83c0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e5",
X"38029a05",
X"33537281",
X"2e098106",
X"81d93802",
X"9b053353",
X"80ce9054",
X"7281aa2e",
X"8d3881c7",
X"3980e451",
X"8d8d3fff",
X"14547380",
X"2e81b838",
X"820a5281",
X"e951fdab",
X"3f83c080",
X"0881ff06",
X"5372de38",
X"725280fa",
X"51fd983f",
X"83c08008",
X"81ff0653",
X"72819038",
X"72547316",
X"53fcdc3f",
X"83c08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e83887",
X"3d337086",
X"2a708106",
X"5154548c",
X"557280e3",
X"38845580",
X"de397452",
X"81e951fc",
X"d23f83c0",
X"800881ff",
X"06538255",
X"81e95681",
X"73278638",
X"735580c1",
X"5680ce90",
X"548a3980",
X"e4518bff",
X"3fff1454",
X"73802ea9",
X"38805275",
X"51fca03f",
X"83c08008",
X"81ff0653",
X"72e13884",
X"805280d0",
X"51fc8c3f",
X"83c08008",
X"81ff0653",
X"72802e83",
X"38805574",
X"83c3c834",
X"fb873ffb",
X"ca3f883d",
X"0d04fb3d",
X"0d775480",
X"0b83c3c8",
X"3370832a",
X"70810651",
X"55575572",
X"752e0981",
X"06853873",
X"892b5473",
X"5280d151",
X"fbc53f83",
X"c0800881",
X"ff065372",
X"bd3882b8",
X"c054fb8b",
X"3f83c080",
X"0881ff06",
X"537281ff",
X"2e098106",
X"8938ff14",
X"5473e738",
X"9f397281",
X"fe2e0981",
X"06963883",
X"c7cc5283",
X"c3cc51fa",
X"f53ffadb",
X"3ffad83f",
X"83398155",
X"fa8b3ffa",
X"ce3f7481",
X"ff0683c0",
X"800c873d",
X"0d04fb3d",
X"0d7783c3",
X"cc5654f9",
X"e63f83c3",
X"c8337083",
X"2a708106",
X"51545672",
X"85387389",
X"2b547352",
X"80d851fa",
X"c23f83c0",
X"800881ff",
X"06537280",
X"e73881ff",
X"51f9e03f",
X"81fe51f9",
X"da3f8480",
X"53747081",
X"05563351",
X"f9cd3fff",
X"137083ff",
X"ff065153",
X"72eb3872",
X"51f9bc3f",
X"7251f9b7",
X"3ff9dc3f",
X"83c08008",
X"9f0653a7",
X"88547285",
X"2e8c389e",
X"3980e451",
X"89bd3fff",
X"1454f9bf",
X"3f83c080",
X"0881ff06",
X"537281ff",
X"2e843873",
X"e438f8e5",
X"3ff9a83f",
X"800b83c0",
X"800c873d",
X"0d047183",
X"c7d00c88",
X"80800b83",
X"c7cc0c84",
X"80800b83",
X"c7d40c04",
X"f03d0d83",
X"80805683",
X"c7d00816",
X"83c7cc08",
X"17565474",
X"33743483",
X"c7d40816",
X"54807434",
X"81165675",
X"8380a02e",
X"098106db",
X"3883d080",
X"5683c7d0",
X"081683c7",
X"cc081756",
X"54743374",
X"3483c7d4",
X"08165480",
X"74348116",
X"567583d0",
X"902e0981",
X"06db3883",
X"a8805683",
X"c7d00816",
X"83c7cc08",
X"17565474",
X"33743483",
X"c7d40816",
X"54807434",
X"81165675",
X"83a8902e",
X"098106db",
X"38805683",
X"c7d00816",
X"83c7d408",
X"17555573",
X"33753481",
X"16567581",
X"80802e09",
X"8106e438",
X"89da3f89",
X"3d58a253",
X"81e19c52",
X"77518195",
X"933f8057",
X"8c805683",
X"c7d40816",
X"77195555",
X"73337534",
X"81168118",
X"585676a2",
X"2e098106",
X"e638860b",
X"87a88334",
X"800b87a8",
X"8234800b",
X"87809a34",
X"af0b8780",
X"9634bf0b",
X"87809734",
X"800b8780",
X"98349f0b",
X"87809934",
X"800b8780",
X"9b34f80b",
X"87a88934",
X"7687a880",
X"34820b87",
X"d08f3482",
X"0b87a881",
X"34840b87",
X"809f34ff",
X"0b87d08b",
X"34923d0d",
X"04fe3d0d",
X"805383c7",
X"d4081383",
X"c7d00814",
X"52527033",
X"72348113",
X"53728180",
X"802e0981",
X"06e43883",
X"80805383",
X"c7d40813",
X"83c7d008",
X"14525270",
X"33723481",
X"13537283",
X"80a02e09",
X"8106e438",
X"83d08053",
X"83c7d408",
X"1383c7d0",
X"08145252",
X"70337234",
X"81135372",
X"83d0902e",
X"098106e4",
X"3883a880",
X"5383c7d4",
X"081383c7",
X"d0081452",
X"52703372",
X"34811353",
X"7283a890",
X"2e098106",
X"e438843d",
X"0d04803d",
X"0d908090",
X"08810683",
X"c0800c82",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe067607",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"812c8106",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fd06",
X"76100772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087082",
X"2cbf0683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fe8306",
X"76822b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"882c8706",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f1ff",
X"0676882b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"708b2c81",
X"0683c080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870ef",
X"ff06768b",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870912c",
X"bf0683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fc87ffff",
X"0676912b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70992c81",
X"0683c080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870ff",
X"bf0a0676",
X"992b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"9008709a",
X"2c830683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70cf0a06",
X"769a2b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"9c2c8706",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f10a",
X"06769c2b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"9080bc08",
X"870683c0",
X"800c823d",
X"0d04ff3d",
X"0d9080bc",
X"700870f8",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"bc087084",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80bc7008",
X"70ef0676",
X"842b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"bc087085",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80bc7008",
X"70df0676",
X"852b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"bc087086",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80bc7008",
X"70ffbf06",
X"76862b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80800870",
X"882c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"70892c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708a2c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708b",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8c2cbf06",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"70922c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"0870932c",
X"810683c0",
X"800c5182",
X"3d0d0471",
X"9080a00c",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727081",
X"055434ff",
X"1151f039",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708405",
X"540cff11",
X"51f03984",
X"3d0d04fe",
X"3d0d8880",
X"53805288",
X"800a51ff",
X"b43f8280",
X"53805282",
X"800a51c8",
X"3f800b87",
X"aa803484",
X"3d0d0480",
X"3d0d8151",
X"f9d53f72",
X"802e9038",
X"8051fbd6",
X"3fc93f81",
X"ea943351",
X"fbcc3f81",
X"51f9e63f",
X"8051f9e1",
X"3f8051f9",
X"b23f823d",
X"0d04fd3d",
X"0d755280",
X"5480ff72",
X"25883881",
X"0bff8013",
X"5354ffbf",
X"12517099",
X"268638e0",
X"1252b039",
X"ff9f1251",
X"997127a7",
X"38d012e0",
X"13545170",
X"89268538",
X"72529839",
X"728f2685",
X"3872528f",
X"3971ba2e",
X"09810685",
X"389a5283",
X"39805273",
X"802e8538",
X"81801252",
X"7181ff06",
X"83c0800c",
X"853d0d04",
X"803d0d84",
X"98c05180",
X"71708105",
X"53347084",
X"a0c02e09",
X"8106f038",
X"823d0d04",
X"fe3d0d02",
X"97053351",
X"fef43f83",
X"c0800881",
X"ff0683c7",
X"dc085452",
X"8073249b",
X"3883c8a4",
X"08137283",
X"c8a80807",
X"53537173",
X"3483c7dc",
X"08810583",
X"c7dc0c84",
X"3d0d04fb",
X"3d0d8056",
X"873dfc05",
X"54785379",
X"527751ff",
X"b8aa3f87",
X"3d0d04fe",
X"3d0d83c7",
X"f8085274",
X"51ffbfae",
X"3f83c080",
X"088c3876",
X"53755283",
X"c7f80851",
X"ca3f843d",
X"0d04fe3d",
X"0d83c7f8",
X"08537552",
X"7451ffb9",
X"ec3f83c0",
X"80088d38",
X"77537652",
X"83c7f808",
X"51ffa43f",
X"843d0d04",
X"f73d0d9c",
X"ec3f83c0",
X"800881ff",
X"06ff0557",
X"76833881",
X"5780e9c8",
X"3f83c080",
X"0883c080",
X"08565a87",
X"15335473",
X"802e80df",
X"38740881",
X"e1d82e09",
X"810680d3",
X"38800b91",
X"16335559",
X"73792e80",
X"c6387456",
X"9a163354",
X"73832e09",
X"8106a438",
X"a4167033",
X"55588052",
X"73519ad6",
X"3f805380",
X"5273519a",
X"f63f8114",
X"54767425",
X"83388054",
X"73783481",
X"1980d817",
X"91173356",
X"57597874",
X"2e098106",
X"ffbe3881",
X"c4158ca0",
X"1b555574",
X"742e0981",
X"06ff8838",
X"8b3d0d04",
X"f63d0d80",
X"e8ba3f83",
X"c080087d",
X"83c08008",
X"58595b77",
X"83c7dc0c",
X"87163355",
X"74802e81",
X"a7387508",
X"547381e5",
X"b82e0981",
X"06933890",
X"16335387",
X"16335281",
X"e6a851e6",
X"fe3f8188",
X"397381e1",
X"d82e0981",
X"0680fd38",
X"745281e6",
X"bc51e6e7",
X"3f807091",
X"1833565b",
X"5973792e",
X"80e638a4",
X"1657f617",
X"33557980",
X"2e9138ff",
X"15547382",
X"268938a8",
X"187083c7",
X"dc0c5874",
X"812e0981",
X"06873881",
X"e6c4518d",
X"3974822e",
X"0981068a",
X"3881e6cc",
X"51e6a03f",
X"95397483",
X"2e098106",
X"8f387633",
X"81055281",
X"e6d851e6",
X"8a3f815a",
X"811980d8",
X"18911833",
X"56585978",
X"742e0981",
X"06ff9f38",
X"a81881c4",
X"178ca01d",
X"56575875",
X"742e0981",
X"06feb838",
X"8c3d0d04",
X"803d0d72",
X"842981ea",
X"98057008",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"72842981",
X"eab40570",
X"0883c080",
X"0c51823d",
X"0d04f73d",
X"0d81eac8",
X"51ffbbb0",
X"3f908090",
X"08599080",
X"bc085a78",
X"57795883",
X"c7e03355",
X"74802e80",
X"ca3883c7",
X"fc085381",
X"e7a85283",
X"c0800851",
X"ffb5f63f",
X"83c08008",
X"b23883c0",
X"8008568b",
X"3dec1155",
X"558853f8",
X"155283c7",
X"fc0851ff",
X"b3de3f76",
X"93f88083",
X"0679ec87",
X"fffc0607",
X"705a9080",
X"900c7990",
X"80bc0c8b",
X"3d0d04f9",
X"3d0d81ea",
X"c851ffba",
X"bf3f9080",
X"90085790",
X"80bc0858",
X"83c7e033",
X"5574802e",
X"80c63883",
X"c7fc0853",
X"81e7a852",
X"83c08008",
X"51ffb589",
X"3f83c080",
X"085583c0",
X"8008a938",
X"83c08008",
X"5283c7fc",
X"0851ffb3",
X"ab3f7456",
X"893df411",
X"55558853",
X"f8155283",
X"c7fc0851",
X"ffb1af3f",
X"ffb0e73f",
X"893d0d04",
X"fd3d0d83",
X"c7f80851",
X"ffb3db3f",
X"83c08008",
X"90802e09",
X"8106ad38",
X"805487c1",
X"80805383",
X"c0800852",
X"83c7f808",
X"51f9f03f",
X"87c18080",
X"143387c1",
X"90801534",
X"81145473",
X"90802e09",
X"8106e938",
X"853d0d04",
X"fd3d0d90",
X"80805286",
X"84808051",
X"ffb4b83f",
X"805483c0",
X"8008742e",
X"098106b4",
X"3883c880",
X"085180fa",
X"d33f81ea",
X"c851ffb8",
X"eb3f83c7",
X"f8085381",
X"e7b45283",
X"c0800851",
X"ffb3ca3f",
X"83c08008",
X"742e0981",
X"068438fe",
X"eb3f8154",
X"7383c080",
X"0c853d0d",
X"0481e7c0",
X"0b83c080",
X"0c04fc3d",
X"0d765473",
X"902e8182",
X"38739024",
X"8e387384",
X"2e983873",
X"862ea738",
X"82bf3973",
X"932e8199",
X"3873942e",
X"81d43882",
X"b0398481",
X"80805382",
X"80805283",
X"c7f40851",
X"f8b53f82",
X"ba398054",
X"84818080",
X"5380c080",
X"5283c7f4",
X"0851f89f",
X"3f848280",
X"805380c0",
X"805283c7",
X"f40851f8",
X"8e3f8481",
X"80801433",
X"8481c080",
X"15348482",
X"80801433",
X"8482c080",
X"15348114",
X"547380c0",
X"802e0981",
X"06dc3881",
X"ee398482",
X"80805381",
X"80805283",
X"c7f40851",
X"f7d53f80",
X"54848280",
X"80143384",
X"81808015",
X"34811454",
X"73818080",
X"2e098106",
X"e83881bf",
X"39848180",
X"805380c0",
X"805283c7",
X"f40851f7",
X"a63f8055",
X"84818080",
X"15547333",
X"8481c080",
X"16347333",
X"84828080",
X"16347333",
X"8482c080",
X"16348115",
X"557480c0",
X"802e0981",
X"06d63880",
X"fe398481",
X"808053a0",
X"805283c7",
X"f40851f6",
X"e63f8055",
X"84818080",
X"15547333",
X"8481a080",
X"16347333",
X"8481c080",
X"16347333",
X"8481e080",
X"16347333",
X"84828080",
X"16347333",
X"8482a080",
X"16347333",
X"8482c080",
X"16347333",
X"8482e080",
X"16348115",
X"5574a080",
X"2e098106",
X"ffb6389f",
X"39f5bd3f",
X"800b83c7",
X"dc0c800b",
X"83c8a80c",
X"81e7c451",
X"dfbd3f81",
X"b78dc051",
X"f3a53f86",
X"3d0d04fc",
X"3d0d7670",
X"5255ffb6",
X"9d3f83c0",
X"80085481",
X"5383c080",
X"0880c238",
X"7451ffb5",
X"df3f83c0",
X"800881e7",
X"e05383c0",
X"80085253",
X"cebf3f83",
X"c08008a1",
X"3881e7e4",
X"527251ce",
X"b03f83c0",
X"80089238",
X"81e7e852",
X"7251cea1",
X"3f83c080",
X"08802e83",
X"38815473",
X"537283c0",
X"800c863d",
X"0d04f03d",
X"0d80de8b",
X"0b83c3ac",
X"0c83c7f4",
X"0851d0cb",
X"3f83c7f4",
X"0851ffab",
X"943fff0b",
X"81e7e453",
X"83c08008",
X"5256cde1",
X"3f83c080",
X"08802e9f",
X"38805892",
X"3dd81155",
X"559053f0",
X"155283c7",
X"f40851ff",
X"ad863f02",
X"bb053356",
X"81a53983",
X"c7f40851",
X"ffae833f",
X"83c08008",
X"5783c080",
X"08828080",
X"2e098106",
X"83388456",
X"83c08008",
X"8180802e",
X"09810680",
X"e138805c",
X"805b805a",
X"8059f3b4",
X"3f800b83",
X"c7dc0c80",
X"0b83c8a8",
X"0c81e7ec",
X"51ddb43f",
X"80d00b83",
X"c7dc0c81",
X"e7fc51dd",
X"a63f80f8",
X"0b83c7dc",
X"0c81e890",
X"51dd983f",
X"758025a2",
X"38805289",
X"3d705255",
X"8db03f83",
X"5274518d",
X"a93f7855",
X"74802583",
X"38905680",
X"7525dd38",
X"86567680",
X"c0802e09",
X"81068538",
X"93568c39",
X"76a0802e",
X"09810683",
X"38945675",
X"51faa73f",
X"923d0d04",
X"f63d0d80",
X"5a805980",
X"58805780",
X"705656f2",
X"ab3f800b",
X"83c7dc0c",
X"800b83c8",
X"a80c81e8",
X"a451dcab",
X"3f81800b",
X"83c8a80c",
X"81e8a851",
X"dc9d3f80",
X"d00b83c7",
X"dc0c7430",
X"70760780",
X"2570872b",
X"83c8a80c",
X"5153eaf7",
X"3f83c080",
X"085281e8",
X"b051dbf7",
X"3f80f80b",
X"83c7dc0c",
X"74813270",
X"30707207",
X"80257087",
X"2b83c8a8",
X"0c515454",
X"f9a33f83",
X"c0800852",
X"81e8bc51",
X"dbcd3f81",
X"a00b83c7",
X"dc0c7482",
X"32703070",
X"72078025",
X"70872b83",
X"c8a80c51",
X"5483c7f8",
X"085254ff",
X"a88b3f83",
X"c0800852",
X"81e8c451",
X"db9d3f81",
X"c80b83c7",
X"dc0c7483",
X"32703070",
X"72078025",
X"70872b83",
X"c8a80c51",
X"5483c7f4",
X"085254ff",
X"a7db3f81",
X"e8cc5383",
X"c0800880",
X"2e8f3883",
X"c7f40851",
X"ffa7c63f",
X"83c08008",
X"53725281",
X"e8d451da",
X"d63f81f0",
X"0b83c7dc",
X"0c748432",
X"70307072",
X"07802570",
X"872b83c8",
X"a80c5154",
X"81e8dc52",
X"54dab43f",
X"82c00b83",
X"c7dc0c74",
X"85327030",
X"70720780",
X"2570872b",
X"83c8a80c",
X"515481e8",
X"f45254da",
X"923f800b",
X"83c8a80c",
X"839051f2",
X"cb3f868d",
X"a051edef",
X"3f805287",
X"3d705253",
X"8a9c3f83",
X"5272518a",
X"953f7953",
X"7281cb38",
X"77155574",
X"80258538",
X"72559039",
X"85752585",
X"38855587",
X"39748526",
X"81aa3874",
X"842981e1",
X"c0055372",
X"0804e8b3",
X"3f83c080",
X"08775553",
X"73812e09",
X"81068938",
X"83c08008",
X"10539039",
X"73ff2e09",
X"81068838",
X"83c08008",
X"812c5390",
X"73258538",
X"90538839",
X"72802483",
X"38815372",
X"51e88d3f",
X"80de39e8",
X"9f3f83c0",
X"80081753",
X"72802585",
X"38805388",
X"39877325",
X"83388753",
X"7251e899",
X"3fbe3976",
X"86387880",
X"2eb63883",
X"c3a40883",
X"c3a00caf",
X"990b83c3",
X"ac0c83c7",
X"f80851ca",
X"d23ff4e8",
X"3f9a3978",
X"802e9538",
X"f9e83f81",
X"53963978",
X"802e8938",
X"efce3f84",
X"39788738",
X"75802efb",
X"de388053",
X"7283c080",
X"0c8c3d0d",
X"04fd3d0d",
X"83c89451",
X"80e8dc3f",
X"83c88451",
X"80e8d43f",
X"8053ebc1",
X"3f83c080",
X"08732e09",
X"81068338",
X"8153800b",
X"83c7e033",
X"53547174",
X"2e098106",
X"83388154",
X"72812e09",
X"81069838",
X"73730652",
X"71802e8f",
X"38f4b93f",
X"83c08008",
X"863883c0",
X"80085380",
X"0b83c7e0",
X"33535471",
X"812e0981",
X"06833871",
X"5472a638",
X"73810652",
X"71802e9d",
X"387283c7",
X"e4555273",
X"70840555",
X"0851ffa4",
X"823f8112",
X"5271882e",
X"098106eb",
X"387283c7",
X"e034e9d8",
X"3f83c080",
X"08802e86",
X"38805180",
X"da39e9dd",
X"3f83c080",
X"0880ce38",
X"e9e83f83",
X"c0800880",
X"2eaa3881",
X"51e5883f",
X"e1c23f80",
X"0b83c7dc",
X"0cf9f93f",
X"83c08008",
X"52ff0b83",
X"c7dc0ce3",
X"d43f71a1",
X"387151e4",
X"e63f9f39",
X"e9c93f83",
X"c0800880",
X"2e943881",
X"51e4d43f",
X"e18e3ff7",
X"cd3fe3b1",
X"3f8151ea",
X"ea3f853d",
X"0d04fd3d",
X"0d805283",
X"c8945180",
X"d78f3f81",
X"5283c884",
X"5180d785",
X"3f828080",
X"53805281",
X"81808051",
X"e9df3f80",
X"c0805380",
X"52848180",
X"8051e9f0",
X"3f8054e9",
X"9c3f83c0",
X"80088338",
X"81547383",
X"c7e03473",
X"81ff0654",
X"73802e92",
X"38f2ad3f",
X"83c08008",
X"893883c0",
X"800883c7",
X"e0348151",
X"ea813ffd",
X"943ffc39",
X"83c08c08",
X"0283c08c",
X"0cfb3d0d",
X"0280d3c4",
X"5383c08c",
X"08fc050c",
X"8051d4fc",
X"3f81e8fc",
X"0b83c3a4",
X"0c81e7e8",
X"0b83c39c",
X"0c81e7e4",
X"0b83c3b4",
X"0c81e980",
X"0b83c3b0",
X"0c81e984",
X"0b83c3a8",
X"0c800b83",
X"c7e40b83",
X"c08c08f8",
X"050c83c0",
X"8c08f405",
X"0cffa4f7",
X"3f83c080",
X"088605fc",
X"0683c08c",
X"08f0050c",
X"0283c08c",
X"08f00508",
X"310d833d",
X"7083c08c",
X"08f80508",
X"70840583",
X"c08c08f8",
X"050c0c51",
X"ffa1883f",
X"83c08c08",
X"f4050881",
X"0583c08c",
X"08f4050c",
X"83c08c08",
X"f4050888",
X"2e098106",
X"ffab3886",
X"94808051",
X"dec83fff",
X"0b83c7dc",
X"0c800b83",
X"c8a80c84",
X"98c00b83",
X"c8a40c81",
X"51e2883f",
X"8151e2ad",
X"3f8051e2",
X"a83f8151",
X"e2ce3f82",
X"51e2f63f",
X"8051e3cb",
X"3f8051e3",
X"f53f8051",
X"e49e3f80",
X"51e4c63f",
X"8051e38a",
X"3fc80b87",
X"809a34fd",
X"913f83c0",
X"8c08fc05",
X"080d800b",
X"83c0800c",
X"873d0d83",
X"c08c0c04",
X"fa3d0d78",
X"5580750c",
X"800b8416",
X"0c800b88",
X"160c800b",
X"8c160c80",
X"0b90160c",
X"83c89451",
X"80e3b83f",
X"83c88451",
X"80e3b03f",
X"e68a3f83",
X"c0800887",
X"d0883370",
X"81ff0651",
X"535671a7",
X"3887d080",
X"3383c8b8",
X"3487d081",
X"3383c8b4",
X"3487d082",
X"3383c8ac",
X"3487d083",
X"3383c8b0",
X"34ff0b87",
X"d08b3487",
X"d0893387",
X"d08f3370",
X"822a7081",
X"06703070",
X"72077009",
X"709f2c77",
X"069e0657",
X"51515651",
X"51545480",
X"74980653",
X"5371882e",
X"09810683",
X"38815371",
X"98327030",
X"70802575",
X"71318419",
X"0c515152",
X"80748606",
X"53537182",
X"2e098106",
X"83388153",
X"71863270",
X"30708025",
X"75713178",
X"0c515152",
X"83c8b833",
X"5281aa72",
X"27843881",
X"750c83c8",
X"b8335271",
X"bb268438",
X"ff750c83",
X"c8b43352",
X"81aa7227",
X"8638810b",
X"84160c83",
X"c8b43352",
X"71bb2686",
X"38ff0b84",
X"160c83c8",
X"ac335281",
X"aa722784",
X"3881750c",
X"83c8ac33",
X"5271bb26",
X"8438ff75",
X"0c83c8b0",
X"335281aa",
X"72278638",
X"810b8416",
X"0c83c8b0",
X"335271bb",
X"268638ff",
X"0b84160c",
X"80577394",
X"2eaa3887",
X"80903387",
X"80913387",
X"80923370",
X"81ff0672",
X"74060687",
X"80933371",
X"06810651",
X"52545454",
X"72772e09",
X"81068338",
X"81577688",
X"160c7580",
X"2eb03875",
X"812a7081",
X"06778106",
X"3184170c",
X"5275832a",
X"76822a71",
X"81067181",
X"0631770c",
X"53537584",
X"2a810688",
X"160c7585",
X"2a81068c",
X"160c883d",
X"0d04fe3d",
X"0d747654",
X"527151fc",
X"c73f7281",
X"2ea23881",
X"73268d38",
X"72822ea8",
X"3872832e",
X"9c38e639",
X"7108e238",
X"841208dd",
X"38881208",
X"d838a539",
X"88120881",
X"2e9e3891",
X"39881208",
X"812e9538",
X"71089138",
X"8412088c",
X"388c1208",
X"812e0981",
X"06ffb238",
X"843d0d04",
X"fb3d0d78",
X"0284059f",
X"05335556",
X"800b81e3",
X"c4565381",
X"732b7406",
X"5271802e",
X"83388152",
X"74708205",
X"56227073",
X"902b0790",
X"809c0c51",
X"81135372",
X"882e0981",
X"06d93880",
X"5383c8c0",
X"13335170",
X"81ff2eb8",
X"38701081",
X"e1e40570",
X"22535171",
X"81ff2ea8",
X"38807317",
X"70337010",
X"81e1e405",
X"70225151",
X"51525471",
X"712e9138",
X"81145473",
X"862e0981",
X"06f13871",
X"90809c0c",
X"81135372",
X"862e0981",
X"06ffb238",
X"80537216",
X"70335151",
X"7081ff2e",
X"9a387010",
X"81e1e405",
X"70225151",
X"7081ff2e",
X"8a387084",
X"80800790",
X"809c0c81",
X"13537286",
X"2e098106",
X"d1388053",
X"72165170",
X"3383c8c0",
X"14348113",
X"5372862e",
X"098106ec",
X"38873d0d",
X"0404fe3d",
X"0d750284",
X"05930533",
X"81065252",
X"70883871",
X"9080940c",
X"8e397081",
X"2e098106",
X"86387190",
X"80980c84",
X"3d0d04fb",
X"3d0d7898",
X"2b70982c",
X"7b982b70",
X"982c0290",
X"059f0533",
X"810683c8",
X"dc117033",
X"70982b70",
X"982c5158",
X"5c5a5651",
X"55515470",
X"742e0981",
X"06943883",
X"c8bc1233",
X"70982b70",
X"982c5152",
X"5670732e",
X"b1387375",
X"347283c8",
X"bc133483",
X"c8bd3383",
X"c8dd3371",
X"982b7190",
X"2b0783c8",
X"bc337088",
X"2b720783",
X"c8dc3371",
X"079080b8",
X"0c525953",
X"5452873d",
X"0d04fe3d",
X"0d748111",
X"33713371",
X"882b0783",
X"c0800c53",
X"51843d0d",
X"0483c8c8",
X"3383c080",
X"0c0483c0",
X"8c080283",
X"c08c0cf5",
X"3d0d83c0",
X"8c088805",
X"0883c08c",
X"088f0533",
X"83c08c08",
X"92052202",
X"8c057390",
X"0583c08c",
X"08e8050c",
X"83c08c08",
X"f8050c83",
X"c08c08f0",
X"050c83c0",
X"8c08ec05",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08f005",
X"0883c08c",
X"08e0050c",
X"83c08c08",
X"fc050c83",
X"c08c08f0",
X"05088927",
X"8a38890b",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"05088605",
X"87fffc06",
X"83c08c08",
X"e0050c02",
X"83c08c08",
X"e0050831",
X"0d853d70",
X"5583c08c",
X"08ec0508",
X"5483c08c",
X"08f00508",
X"5383c08c",
X"08f40508",
X"5283c08c",
X"08e4050c",
X"80e1b73f",
X"83c08008",
X"81ff0683",
X"c08c08e4",
X"050883c0",
X"8c08ec05",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"e0050880",
X"2e8c3883",
X"c08c08f8",
X"05080d89",
X"c83983c0",
X"8c08f005",
X"08802e89",
X"a63883c0",
X"8c08ec05",
X"08810533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508842e",
X"a938840b",
X"83c08c08",
X"e0050825",
X"88c73883",
X"c08c08e0",
X"0508852e",
X"859b3883",
X"c08c08e0",
X"0508a12e",
X"87ad3888",
X"ac39800b",
X"83c08c08",
X"ec050885",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08fc050c",
X"83c08c08",
X"e0050883",
X"2e098106",
X"88833883",
X"c08c08e8",
X"05088105",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e0050881",
X"2687e638",
X"810b83c0",
X"8c08e005",
X"0880d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08fc",
X"050c83c0",
X"8c08ec05",
X"08820533",
X"83c08c08",
X"e0050887",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088b",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"e005088c",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088d",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"e005088e",
X"052383c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088a",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"70940508",
X"fcffff06",
X"7194050c",
X"83c08c08",
X"e0050c83",
X"c08c08ec",
X"05088605",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"f4050c83",
X"c08c08e0",
X"050883c0",
X"8c08fc05",
X"082e0981",
X"06b63883",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c83",
X"c08c08fc",
X"050883c0",
X"8c08e005",
X"088b0534",
X"83c08c08",
X"ec050887",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"812e8f38",
X"83c08c08",
X"e0050882",
X"2eb73884",
X"8c3983c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c820b",
X"83c08c08",
X"e005088a",
X"053483d9",
X"3983c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08fc0508",
X"83c08c08",
X"e005088a",
X"053483a1",
X"3983c08c",
X"08fc0508",
X"802e8395",
X"3883c08c",
X"08ec0508",
X"83053383",
X"0683c08c",
X"08e0050c",
X"83c08c08",
X"e0050883",
X"2e098106",
X"82f33883",
X"c08c08ec",
X"05088205",
X"3370982b",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c83c0",
X"8c08e005",
X"08802582",
X"cc3883c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c83c0",
X"8c08ec05",
X"08860533",
X"83c08c08",
X"e0050880",
X"d6053483",
X"c08c08e0",
X"05088405",
X"83c08c08",
X"ec050882",
X"05338f06",
X"83c08c08",
X"e4050c83",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0883c08c",
X"08e00508",
X"3483c08c",
X"08ec0508",
X"84053383",
X"c08c08e0",
X"05088105",
X"34800b83",
X"c08c08e0",
X"05088205",
X"3483c08c",
X"08e00508",
X"08ff83ff",
X"06828007",
X"83c08c08",
X"e005080c",
X"83c08c08",
X"e8050881",
X"05338105",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"050883c0",
X"8c08e805",
X"08810534",
X"81833983",
X"c08c08fc",
X"0508802e",
X"80f73883",
X"c08c08ec",
X"05088605",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e00508a2",
X"2e098106",
X"80d73883",
X"c08c08ec",
X"05088805",
X"3383c08c",
X"08ec0508",
X"87053371",
X"82802905",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c5283c0",
X"8c08e405",
X"0c83c08c",
X"08f4050c",
X"83c08c08",
X"e4050883",
X"c08c08e0",
X"05088805",
X"2383c08c",
X"08ec0508",
X"3383c08c",
X"08f00508",
X"71317083",
X"ffff0683",
X"c08c08f0",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08ec0508",
X"0583c08c",
X"08ec050c",
X"f6d03983",
X"c08c08f8",
X"05080d83",
X"c08c08f0",
X"050883c0",
X"8c08e005",
X"0c83c08c",
X"08f80508",
X"0d83c08c",
X"08e00508",
X"83c0800c",
X"8d3d0d83",
X"c08c0c04",
X"83c08c08",
X"0283c08c",
X"0ce73d0d",
X"83c08c08",
X"88050802",
X"840583c0",
X"8c08e805",
X"0c83c08c",
X"08d4050c",
X"800b83c8",
X"e43483c0",
X"8c08d405",
X"08900583",
X"c08c08c4",
X"050c800b",
X"83c08c08",
X"c4050834",
X"800b83c0",
X"8c08c405",
X"08810534",
X"800b83c0",
X"8c08c805",
X"0c83c08c",
X"08c80508",
X"80d82983",
X"c08c08c4",
X"05080583",
X"c08c08ff",
X"b8050c80",
X"0b83c08c",
X"08ffb805",
X"0880d805",
X"0c83c08c",
X"08ffb805",
X"08840583",
X"c08c08ff",
X"b8050c83",
X"c08c08c8",
X"050883c0",
X"8c08ffb8",
X"05083488",
X"0b83c08c",
X"08ffb805",
X"08810534",
X"800b83c0",
X"8c08ffb8",
X"05088205",
X"3483c08c",
X"08ffb805",
X"0808ffa1",
X"ff06a080",
X"0783c08c",
X"08ffb805",
X"080c83c0",
X"8c08c805",
X"08810570",
X"81ff0683",
X"c08c08c8",
X"050c83c0",
X"8c08ffb8",
X"050c810b",
X"83c08c08",
X"c8050827",
X"fedb3883",
X"c08c08ec",
X"05705483",
X"c08c08cc",
X"050c9252",
X"83c08c08",
X"d4050851",
X"80d4de3f",
X"83c08008",
X"81ff0670",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffbc0508",
X"90c93883",
X"c08c08f4",
X"0551f1ca",
X"3f83c080",
X"0883ffff",
X"0683c08c",
X"08f60552",
X"83c08c08",
X"dc050cf1",
X"b13f83c0",
X"800883ff",
X"ff0683c0",
X"8c08fd05",
X"3383c08c",
X"08ffbc05",
X"0883c08c",
X"08c8050c",
X"83c08c08",
X"c0050c83",
X"c08c08d8",
X"050c83c0",
X"8c08c805",
X"0883c08c",
X"08c00508",
X"2780fe38",
X"83c08c08",
X"cc050854",
X"83c08c08",
X"c8050853",
X"895283c0",
X"8c08d405",
X"085180d3",
X"e53f83c0",
X"800881ff",
X"0683c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffbc05",
X"0883eb38",
X"83c08c08",
X"ee0551f0",
X"b13f83c0",
X"800883ff",
X"ff065383",
X"c08c08c8",
X"05085283",
X"c08c08d4",
X"050851f0",
X"b53f83c0",
X"8c08c805",
X"08810570",
X"81ff0683",
X"c08c08c8",
X"050c83c0",
X"8c08ffb8",
X"050cfef2",
X"3983c08c",
X"08c40508",
X"81053383",
X"c08c08c0",
X"050c83c0",
X"8c08c005",
X"08839e38",
X"83c08c08",
X"c0050883",
X"c08c08ff",
X"b8050c83",
X"c08c08dc",
X"050888de",
X"2e098106",
X"8b38810b",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"d8050885",
X"8e2e0981",
X"0682c538",
X"817083c0",
X"8c08ffb8",
X"05080683",
X"c08c08ff",
X"b8050c83",
X"c08c08c8",
X"050c83c0",
X"8c08ffb8",
X"0508802e",
X"829e3883",
X"c08c08c8",
X"050883c0",
X"8c08c405",
X"08810534",
X"83c08c08",
X"c0050883",
X"c08c08c4",
X"05088705",
X"3483c08c",
X"08c00508",
X"83c08c08",
X"c405088b",
X"053483c0",
X"8c08c005",
X"0883c08c",
X"08c40508",
X"8c053483",
X"0b83c08c",
X"08c40508",
X"8d053483",
X"c08c08c0",
X"050883c0",
X"8c08c405",
X"088e0523",
X"830b83c0",
X"8c08c405",
X"088a0534",
X"83c08c08",
X"c4050894",
X"05088380",
X"800783c0",
X"8c08c405",
X"0894050c",
X"83c8c833",
X"7083c08c",
X"08c80508",
X"0583c08c",
X"08ffb805",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffb805",
X"0883c8c8",
X"3483c08c",
X"08ffbc05",
X"0883c08c",
X"08c40508",
X"94053483",
X"c08c08c8",
X"050883c0",
X"8c08c405",
X"0880d605",
X"3483c08c",
X"08c80508",
X"83c08c08",
X"c4050884",
X"05348e0b",
X"83c08c08",
X"c4050885",
X"053483c0",
X"8c08c005",
X"0883c08c",
X"08c40508",
X"86053483",
X"c08c08c4",
X"05088405",
X"08ff83ff",
X"06828007",
X"83c08c08",
X"c4050884",
X"050ca239",
X"81db0b83",
X"c08c08ff",
X"b8050c8b",
X"c63983c0",
X"8c08ffbc",
X"050883c0",
X"8c08ffb8",
X"050c8bb3",
X"3983c08c",
X"08f10533",
X"5283c08c",
X"08d40508",
X"5180cfea",
X"3f800b83",
X"c08c08c4",
X"05088105",
X"3383c08c",
X"08ffb805",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"c8050883",
X"c08c08ff",
X"b8050827",
X"89ba3883",
X"c08c08c8",
X"050880d8",
X"297083c0",
X"8c08c405",
X"08057088",
X"05708305",
X"3383c08c",
X"08ffb805",
X"0c83c08c",
X"08cc050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"b8050886",
X"fd3883c0",
X"8c08ffbc",
X"05088d05",
X"3383c08c",
X"08d0050c",
X"83c08c08",
X"d0050886",
X"e13883c0",
X"8c08cc05",
X"08220284",
X"05718605",
X"87fffc06",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"e0050c83",
X"c08c08c0",
X"050c0283",
X"c08c08ff",
X"b8050831",
X"0d893d70",
X"5983c08c",
X"08c00508",
X"5883c08c",
X"08ffbc05",
X"08870533",
X"5783c08c",
X"08ffb805",
X"0ca25583",
X"c08c08d0",
X"05085486",
X"53818152",
X"83c08c08",
X"d4050851",
X"80c29d3f",
X"83c08008",
X"81ff0683",
X"c08c08d0",
X"050c83c0",
X"8c08d005",
X"0881c038",
X"83c08c08",
X"ffbc0508",
X"96055383",
X"c08c08c0",
X"05085283",
X"c08c08ff",
X"b8050851",
X"a5d53f83",
X"c0800881",
X"ff0683c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"0508802e",
X"81853883",
X"c08c08ff",
X"bc050894",
X"0583c08c",
X"08ffbc05",
X"08960533",
X"70862a83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08c0",
X"050c83c0",
X"8c08ffb8",
X"0508832e",
X"09810680",
X"c63883c0",
X"8c08ffb8",
X"050883c0",
X"8c08cc05",
X"08820534",
X"83c8c833",
X"70810583",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"b8050883",
X"c8c83483",
X"c08c08ff",
X"bc050883",
X"c08c08c0",
X"05083483",
X"c08c08e0",
X"05080d83",
X"c08c08d0",
X"050881ff",
X"0683c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffbc05",
X"08fbe338",
X"83c08c08",
X"c8050883",
X"ed3883c0",
X"8c08c805",
X"0883c08c",
X"08ffb805",
X"0c83c08c",
X"08dc0508",
X"80f92e09",
X"81068b38",
X"810b83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08d805",
X"08912e09",
X"81068181",
X"3883c08c",
X"08ffb805",
X"08810683",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b8050880",
X"2e80e238",
X"850b83c0",
X"8c08c405",
X"08a60534",
X"a00b83c0",
X"8c08c405",
X"08a70534",
X"850b83c0",
X"8c08c405",
X"08a80534",
X"80c00b83",
X"c08c08c4",
X"0508a905",
X"34860b83",
X"c08c08c4",
X"0508aa05",
X"34900b83",
X"c08c08c4",
X"0508ab05",
X"34860b83",
X"c08c08c4",
X"0508ac05",
X"34a00b83",
X"c08c08c4",
X"0508ad05",
X"3483c08c",
X"08dc0508",
X"89d83270",
X"30708025",
X"515183c0",
X"8c08ffb8",
X"050c83c0",
X"8c08d805",
X"0883edec",
X"2e098106",
X"80ec3881",
X"7083c08c",
X"08ffb805",
X"080683c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb8",
X"0508802e",
X"80c43884",
X"0b83c08c",
X"08c40508",
X"aa053480",
X"c00b83c0",
X"8c08c405",
X"08ab0534",
X"840b83c0",
X"8c08c405",
X"08ac0534",
X"900b83c0",
X"8c08c405",
X"08ad0534",
X"83c08c08",
X"ffbc0508",
X"83c08c08",
X"c405088c",
X"053483c0",
X"8c08dc05",
X"0880f932",
X"70307080",
X"25515183",
X"c08c08ff",
X"b8050c83",
X"c08c08d8",
X"0508862e",
X"098106ba",
X"38817083",
X"c08c08ff",
X"b8050806",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb80508",
X"802e9338",
X"83c08c08",
X"ffbc0508",
X"83c08c08",
X"c405088d",
X"053483c0",
X"8c08dc05",
X"08b4b432",
X"70307080",
X"25515183",
X"c08c08ff",
X"b8050c83",
X"c08c08d8",
X"05089089",
X"2e098106",
X"993883c0",
X"8c08ffb8",
X"0508802e",
X"8d38820b",
X"83c08c08",
X"c405088d",
X"053483c0",
X"8c08e405",
X"0883c08c",
X"08c40508",
X"05708405",
X"70830533",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"cc050c83",
X"c08c08c0",
X"050c8058",
X"805783c0",
X"8c08ffb8",
X"05085680",
X"5580548a",
X"53a15283",
X"c08c08d4",
X"050851bb",
X"df3f83c0",
X"800881ff",
X"06703070",
X"9f2a5183",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"bc0508a0",
X"2e8c3883",
X"c08c08ff",
X"b80508f6",
X"ed3883c0",
X"8c08c005",
X"088b0533",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"802eb338",
X"83c08c08",
X"cc050883",
X"053383c0",
X"8c08ffb8",
X"050c8058",
X"805783c0",
X"8c08ffb8",
X"05085680",
X"5580548b",
X"53a15283",
X"c08c08d4",
X"050851ba",
X"db3f83c0",
X"8c08c805",
X"08810570",
X"81ff0683",
X"c08c08c4",
X"05088105",
X"335283c0",
X"8c08c805",
X"0c83c08c",
X"08ffb805",
X"0cf6b539",
X"800b83c0",
X"8c08c805",
X"0c83c08c",
X"08c80508",
X"80d82983",
X"c08c08d4",
X"05080570",
X"9a053383",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050882",
X"2e098106",
X"bd3883c0",
X"8c08ffb8",
X"05089705",
X"3383c8e4",
X"5983c08c",
X"08ffb805",
X"0c815783",
X"c08c08ff",
X"b8050856",
X"83c08c08",
X"ffbc0508",
X"55805489",
X"53a15283",
X"c08c08d4",
X"050851b9",
X"b73f83c0",
X"8c08c805",
X"08810570",
X"81ff0683",
X"c08c08c8",
X"050c83c0",
X"8c08ffb8",
X"050c810b",
X"83c08c08",
X"c8050827",
X"fee73881",
X"0b83c08c",
X"08c40508",
X"34800b83",
X"c08c08ff",
X"b8050c83",
X"c08c08e8",
X"05080d83",
X"c08c08ff",
X"b8050883",
X"c0800c9b",
X"3d0d83c0",
X"8c0c04f4",
X"3d0d901f",
X"59800b81",
X"1a33555b",
X"7a742781",
X"ad387a80",
X"d829198a",
X"11335555",
X"73832e09",
X"81068188",
X"38941533",
X"57805276",
X"51df9b3f",
X"80538052",
X"7651dfbb",
X"3fadb93f",
X"83c08008",
X"5c805877",
X"81c4291c",
X"87113355",
X"5573802e",
X"80c03874",
X"0881e1d8",
X"2e098106",
X"b5388075",
X"5b567580",
X"d8291a9a",
X"11335555",
X"73832e09",
X"81069238",
X"a4157033",
X"55557674",
X"278738ff",
X"14547375",
X"34811670",
X"81ff0657",
X"54817627",
X"d1388118",
X"7081ff06",
X"59548778",
X"27ffa438",
X"83c8c833",
X"ff055473",
X"83c8c834",
X"811b7081",
X"ff06811b",
X"335f5c54",
X"7c7b26fe",
X"d538800b",
X"83c0800c",
X"8e3d0d04",
X"83c08c08",
X"0283c08c",
X"0cda3d0d",
X"83c08c08",
X"88050802",
X"84057190",
X"05703370",
X"83c08c08",
X"fef8050c",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"ff9c050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"fef40508",
X"802e9a96",
X"38800b83",
X"c08c08ff",
X"9c050881",
X"053383c0",
X"8c08fef4",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08fef4",
X"05082599",
X"db3883c0",
X"8c08ffa4",
X"050880d8",
X"2983c08c",
X"08ff9c05",
X"08058405",
X"70860533",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"ff88050c",
X"83c08c08",
X"fef40508",
X"802e98e1",
X"38aadd3f",
X"83c08c08",
X"ff880508",
X"80d40508",
X"83c08008",
X"2698ca38",
X"0283c08c",
X"08ff8805",
X"08810533",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"fef40508",
X"83c08c08",
X"fc052383",
X"c08c08fe",
X"f4050886",
X"0583fc06",
X"83c08c08",
X"fef4050c",
X"0283c08c",
X"08fef405",
X"08310d85",
X"3d705583",
X"c08c08fc",
X"055483c0",
X"8c08ff88",
X"05085383",
X"c08c08ff",
X"b0050852",
X"83c08c08",
X"ff90050c",
X"b2ae3f83",
X"c0800881",
X"ff0683c0",
X"8c08fef4",
X"050c83c0",
X"8c08fef4",
X"0508978f",
X"3883c08c",
X"08ff8805",
X"08870533",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"fef40508",
X"802e80d7",
X"3883c08c",
X"08ff8805",
X"08860533",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"fef40508",
X"822e0981",
X"06b53883",
X"c08c08fc",
X"052283c0",
X"8c08fef4",
X"050c870b",
X"83c08c08",
X"fef40508",
X"27993883",
X"c08c08ff",
X"90050882",
X"055283c0",
X"8c08ff90",
X"05083351",
X"d8d63f83",
X"c08c08ff",
X"88050886",
X"053383c0",
X"8c08fef4",
X"050c83c0",
X"8c08fef4",
X"0508832e",
X"09810695",
X"f63883c0",
X"8c08ff88",
X"05089205",
X"83c08c08",
X"ff880508",
X"89053383",
X"c08c08fe",
X"f4050c83",
X"c08c08ff",
X"94050c83",
X"c08c08fe",
X"f4050883",
X"2eb73883",
X"c08c08ff",
X"94050882",
X"053383c0",
X"8c08fc05",
X"2283c08c",
X"08fefc05",
X"0c83c08c",
X"08fef805",
X"0c83c08c",
X"08fef805",
X"0883c08c",
X"08fefc05",
X"0826958f",
X"38800b83",
X"c08c08ff",
X"b4050c80",
X"0b83c08c",
X"08ff8c05",
X"0c83c08c",
X"08fef405",
X"08832e09",
X"81068398",
X"3883c08c",
X"08ff9005",
X"083383c0",
X"8c08fef8",
X"050c83c0",
X"8c08fef8",
X"050883c0",
X"8c08ff8c",
X"05082e09",
X"810682d9",
X"3883c08c",
X"08ff9005",
X"08810533",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"fef40508",
X"942e0981",
X"0682b638",
X"b05381e4",
X"cc5283c0",
X"8c08c805",
X"5180c780",
X"3f83c08c",
X"08fef805",
X"0883c08c",
X"08ff8c05",
X"0c83c08c",
X"08ff8c05",
X"081083c0",
X"8c08ff8c",
X"05080583",
X"c08c0805",
X"c8057033",
X"83c08c08",
X"ff900508",
X"05703372",
X"81053371",
X"06515183",
X"c08c08fe",
X"f4050c83",
X"c08c08fe",
X"f8050c83",
X"c08c08fe",
X"f4050880",
X"2ea83883",
X"c08c08fe",
X"f8050882",
X"05338171",
X"2b83c08c",
X"08ffb405",
X"080783c0",
X"8c08ffb4",
X"050c83c0",
X"8c08fef8",
X"050c83c0",
X"8c08ff8c",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ff8c050c",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"ff8c0508",
X"902e0981",
X"06fee238",
X"83c08c08",
X"ff900508",
X"87053370",
X"982b83c0",
X"8c08ff90",
X"05088905",
X"3370982b",
X"70982c73",
X"982c8180",
X"05545153",
X"83c08c08",
X"fefc050c",
X"83c08c08",
X"fef8050c",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"fef80508",
X"83c08c08",
X"f8052380",
X"ff0b83c0",
X"8c08fef4",
X"05083183",
X"c08c08fe",
X"f4050c83",
X"c08c08fe",
X"f4050883",
X"c08c08fa",
X"052384d7",
X"3981800b",
X"83c08c08",
X"f8052381",
X"800b83c0",
X"8c08fa05",
X"2384c039",
X"83c08c08",
X"ff8c0508",
X"1083c08c",
X"0805f805",
X"83c08c08",
X"ff8c0508",
X"842983c0",
X"8c08ff8c",
X"05081005",
X"83c08c08",
X"ff940508",
X"05708405",
X"703383c0",
X"8c08ff90",
X"05080570",
X"3383c08c",
X"08ff8005",
X"0c83c08c",
X"08fef405",
X"0c83c08c",
X"08fef805",
X"0c83c08c",
X"08fefc05",
X"0c83c08c",
X"08ff8405",
X"0c83c08c",
X"08ff8005",
X"0883c08c",
X"08ff8405",
X"082383c0",
X"8c08fef8",
X"05088105",
X"3383c08c",
X"08fef405",
X"0c83c08c",
X"08fef405",
X"08902e09",
X"8106bf38",
X"83c08c08",
X"fef80508",
X"3383c08c",
X"08ff9005",
X"08058105",
X"70337082",
X"802983c0",
X"8c08ff80",
X"05080551",
X"5183c08c",
X"08fef405",
X"0c83c08c",
X"08fef405",
X"0883c08c",
X"08ff8405",
X"082383c0",
X"8c08fefc",
X"05088605",
X"2283c08c",
X"08fef805",
X"0c83c08c",
X"08fef805",
X"08a23883",
X"c08c08fe",
X"fc050888",
X"052283c0",
X"8c08fef4",
X"050c83c0",
X"8c08fef4",
X"050881ff",
X"2e80e538",
X"83c08c08",
X"ff840508",
X"227083c0",
X"8c08fef8",
X"05083170",
X"82802971",
X"3183c08c",
X"08fefc05",
X"08880522",
X"7083c08c",
X"08fef805",
X"08317073",
X"355383c0",
X"8c08fef8",
X"050c83c0",
X"8c08fefc",
X"050c5183",
X"c08c08fe",
X"f4050c83",
X"c08c08ff",
X"80050c83",
X"c08c08fe",
X"f4050883",
X"c08c08ff",
X"84050823",
X"83c08c08",
X"ff8c0508",
X"81057081",
X"ff0683c0",
X"8c08ff8c",
X"050c83c0",
X"8c08fef4",
X"050c810b",
X"83c08c08",
X"ff8c0508",
X"27fcdd38",
X"800b83c0",
X"8c08ff8c",
X"050c83c0",
X"8c08ff8c",
X"05081083",
X"c08c08ff",
X"94050805",
X"70900570",
X"3383c08c",
X"08ff9005",
X"08057033",
X"72810533",
X"70720651",
X"535183c0",
X"8c08fef8",
X"050c5183",
X"c08c08fe",
X"f4050c83",
X"c08c08fe",
X"f4050880",
X"2e9d3890",
X"0b83c08c",
X"08ff8c05",
X"082b83c0",
X"8c08ffb4",
X"05080783",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"8c050881",
X"057081ff",
X"0683c08c",
X"08ff8c05",
X"0c83c08c",
X"08fef405",
X"0c970b83",
X"c08c08ff",
X"8c050827",
X"fef03883",
X"c08c08f8",
X"052283c0",
X"8c08fef4",
X"050c83c0",
X"8c08fef4",
X"0508bf26",
X"933883c0",
X"8c08ffb4",
X"05088207",
X"83c08c08",
X"ffb4050c",
X"81c00b83",
X"c08c08fe",
X"f4050827",
X"933883c0",
X"8c08ffb4",
X"05088107",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"fa052283",
X"c08c08fe",
X"f4050c83",
X"c08c08fe",
X"f40508bf",
X"26933883",
X"c08c08ff",
X"b4050888",
X"0783c08c",
X"08ffb405",
X"0c81c00b",
X"83c08c08",
X"fef40508",
X"27933883",
X"c08c08ff",
X"b4050884",
X"0783c08c",
X"08ffb405",
X"0c83c08c",
X"08ff8805",
X"08900533",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"ff94050c",
X"83c08c08",
X"fef40508",
X"83c08c08",
X"ff880508",
X"8c05082e",
X"85e93883",
X"c08c08fe",
X"f4050883",
X"c08c08ff",
X"8805088c",
X"050c83c0",
X"8c08ff88",
X"05088905",
X"3383c08c",
X"08fef805",
X"0c83c08c",
X"08fef805",
X"08802e85",
X"a13883c0",
X"8c08ffb4",
X"0583c08c",
X"08fef405",
X"0883c08c",
X"08fef405",
X"088f0683",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"80050c83",
X"c08c08ff",
X"a0050c83",
X"c08c08fe",
X"f8050882",
X"2e098106",
X"81c23880",
X"0b83c08c",
X"08fef405",
X"08862a70",
X"81065183",
X"c08c08fe",
X"f4050c83",
X"c08c08fe",
X"f8050c83",
X"c08c08fe",
X"f4050883",
X"c08c08fe",
X"f805082e",
X"8c3881c0",
X"0b83c08c",
X"08fef805",
X"0c83c08c",
X"08ff8005",
X"08872a70",
X"81065183",
X"c08c08fe",
X"f4050c83",
X"c08c08fe",
X"f4050880",
X"2e943883",
X"c08c08fe",
X"f8050881",
X"903283c0",
X"8c08fef8",
X"050c83c0",
X"8c08ff80",
X"0508842a",
X"70810651",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"fef40508",
X"802e9438",
X"83c08c08",
X"fef80508",
X"80d03283",
X"c08c08fe",
X"f8050c83",
X"c08c08ff",
X"80050883",
X"c08c08fe",
X"f8050832",
X"83c08c08",
X"ff80050c",
X"800b83c0",
X"8c08c005",
X"0c800b83",
X"c08c08c4",
X"0523800b",
X"81e3d433",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"ff8c050c",
X"83c08c08",
X"fef40508",
X"83c08c08",
X"ff8c0508",
X"2e82d738",
X"83c08c08",
X"c00581e3",
X"d40b83c0",
X"8c08fefc",
X"050c83c0",
X"8c08ff98",
X"050c83c0",
X"8c08fefc",
X"05083383",
X"c08c08fe",
X"fc050881",
X"05338172",
X"2b81722b",
X"077083c0",
X"8c08ff80",
X"05080653",
X"83c08c08",
X"fef8050c",
X"83c08c08",
X"ff84050c",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"fef40508",
X"83c08c08",
X"fef80508",
X"2e098106",
X"81c13883",
X"c08c08ff",
X"8c050885",
X"2680f738",
X"83c08c08",
X"fefc0508",
X"82053370",
X"81ff0683",
X"c08c08fe",
X"f4050c83",
X"c08c08ff",
X"84050c83",
X"c08c08fe",
X"f4050880",
X"2e80cb38",
X"83c08c08",
X"ff8c0508",
X"83c08c08",
X"ff8c0508",
X"81057081",
X"ff0683c0",
X"8c08ff98",
X"05087305",
X"5383c08c",
X"08ff8c05",
X"0c83c08c",
X"08fef805",
X"0c83c08c",
X"08fef405",
X"0c83c08c",
X"08ff8405",
X"0883c08c",
X"08fef405",
X"083483c0",
X"8c08fefc",
X"05088305",
X"3383c08c",
X"08fef405",
X"0c83c08c",
X"08fef405",
X"08802e9f",
X"38810b83",
X"c08c08fe",
X"f405082b",
X"83c08c08",
X"ffa00508",
X"080783c0",
X"8c08ffa0",
X"05080c83",
X"c08c08fe",
X"fc050884",
X"05703383",
X"c08c08fe",
X"f4050c83",
X"c08c08fe",
X"fc050c83",
X"c08c08fe",
X"f40508fd",
X"c53883c0",
X"8c08c005",
X"528051c8",
X"ab3f83c0",
X"8c08ffb4",
X"05085283",
X"c08c08ff",
X"94050851",
X"c9f03f83",
X"c08c08fb",
X"05337081",
X"800a2981",
X"0a057098",
X"2c5583c0",
X"8c08fef4",
X"050c83c0",
X"8c08f905",
X"33708180",
X"0a29810a",
X"0570982c",
X"5583c08c",
X"08fef405",
X"0c83c08c",
X"08ff9405",
X"085383c0",
X"8c08fefc",
X"050c83c0",
X"8c08fef8",
X"050cc9c7",
X"3f83c08c",
X"08ff8805",
X"08880533",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"fef40508",
X"802e84e7",
X"3883c08c",
X"08ff8805",
X"08900533",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"fef40508",
X"812684c7",
X"38807081",
X"e48c0b81",
X"e48c0b81",
X"053383c0",
X"8c08fef4",
X"050c83c0",
X"8c08fef8",
X"050c83c0",
X"8c08fefc",
X"050c83c0",
X"8c08ff84",
X"050c83c0",
X"8c08fef4",
X"050883c0",
X"8c08ff84",
X"05082e81",
X"af3883c0",
X"8c08fefc",
X"05088429",
X"83c08c08",
X"fef80508",
X"05703383",
X"c08c08ff",
X"90050805",
X"70337281",
X"05337072",
X"06515351",
X"83c08c08",
X"fef8050c",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"fef40508",
X"802eaa38",
X"810b83c0",
X"8c08fefc",
X"05082b83",
X"c08c08ff",
X"84050807",
X"7083ffff",
X"0683c08c",
X"08ff8405",
X"0c83c08c",
X"08fef405",
X"0c83c08c",
X"08fefc05",
X"08810570",
X"81ff0681",
X"e48c7184",
X"29710570",
X"81053351",
X"5383c08c",
X"08fef805",
X"0c83c08c",
X"08fefc05",
X"0c83c08c",
X"08fef405",
X"0c83c08c",
X"08fef405",
X"08fed338",
X"83c08c08",
X"ff880508",
X"8a052283",
X"c08c08ff",
X"90050c83",
X"c08c08ff",
X"84050883",
X"c08c08ff",
X"9005082e",
X"82b13880",
X"0b83c08c",
X"08ffb805",
X"0c800b83",
X"c08c08ff",
X"bc052380",
X"7083c08c",
X"08ffb805",
X"83c08c08",
X"ff8c050c",
X"83c08c08",
X"fefc050c",
X"83c08c08",
X"ff80050c",
X"81af3983",
X"c08c08ff",
X"84050883",
X"c08c08fe",
X"fc05082c",
X"70810651",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"fef40508",
X"802e80e7",
X"3883c08c",
X"08ff8005",
X"0883c08c",
X"08ff8005",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"8c050873",
X"0583c08c",
X"08ff8805",
X"08900533",
X"83c08c08",
X"fefc0508",
X"84290553",
X"5383c08c",
X"08ff8005",
X"0c83c08c",
X"08fef805",
X"0c83c08c",
X"08fef405",
X"0c83c08c",
X"08fef805",
X"0881e48e",
X"053383c0",
X"8c08fef4",
X"05083483",
X"c08c08fe",
X"fc050881",
X"057081ff",
X"0683c08c",
X"08fefc05",
X"0c83c08c",
X"08fef405",
X"0c8f0b83",
X"c08c08fe",
X"fc050827",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"ff800508",
X"85268c38",
X"83c08c08",
X"fef40508",
X"fea93883",
X"c08c08ff",
X"b8055280",
X"51c2d13f",
X"83c08c08",
X"ff840508",
X"83c08c08",
X"ff880508",
X"8a052383",
X"c08c08ff",
X"88050880",
X"d2053383",
X"c08c08ff",
X"88050880",
X"d4050805",
X"83c08c08",
X"ff880508",
X"80d4050c",
X"83c08c08",
X"ffa80508",
X"0d83c08c",
X"08ffa405",
X"0881800a",
X"2981800a",
X"0570982c",
X"83c08c08",
X"ff9c0508",
X"81053383",
X"c08c08fe",
X"f8050c51",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"fef80508",
X"83c08c08",
X"ffa40508",
X"24e6a738",
X"800b83c0",
X"8c08fef8",
X"050c83c0",
X"8c08ffac",
X"05080d83",
X"c08c08fe",
X"f8050883",
X"c0800ca8",
X"3d0d83c0",
X"8c0c04e9",
X"3d0d696c",
X"02880580",
X"ea05225c",
X"5a5b8070",
X"71415e58",
X"ff78797a",
X"7b7c7d46",
X"4c4a4540",
X"5d436299",
X"3d346202",
X"840580dd",
X"05347779",
X"2280ffff",
X"06544572",
X"79237978",
X"2e888738",
X"7a708105",
X"5c337084",
X"2a718c06",
X"70822a5a",
X"56568306",
X"ff1b7083",
X"ffff065c",
X"54568054",
X"75742e91",
X"387a7081",
X"055c33ff",
X"1b7083ff",
X"ff065c54",
X"54817627",
X"9b387381",
X"ff067b70",
X"81055d33",
X"55748280",
X"2905ff1b",
X"7083ffff",
X"065c5454",
X"827627aa",
X"387383ff",
X"ff067b70",
X"81055d33",
X"70902b72",
X"077d7081",
X"055f3370",
X"982b7207",
X"fe1f7083",
X"ffff0640",
X"52525252",
X"54547e80",
X"2e80c438",
X"7686f738",
X"748a2e09",
X"81069438",
X"811f7081",
X"ff06811e",
X"7081ff06",
X"5f524053",
X"86dc3974",
X"8c2e0981",
X"0686d338",
X"ff1f7081",
X"ff06ff1e",
X"7081ff06",
X"5f524053",
X"7b632586",
X"bd38ff43",
X"86b83976",
X"812e83bb",
X"38768124",
X"89387680",
X"2e8d3886",
X"a5397682",
X"2e84a638",
X"869c39f8",
X"15537284",
X"26849538",
X"72842981",
X"e4fc0553",
X"72080464",
X"802e80cd",
X"38782283",
X"80800653",
X"72838080",
X"2e098106",
X"bc388056",
X"756427a4",
X"38751e70",
X"83ffff06",
X"77101b90",
X"1172832a",
X"58515751",
X"53737534",
X"72870681",
X"712b5153",
X"72811634",
X"81167081",
X"ff065753",
X"977627cc",
X"387f8407",
X"40800b99",
X"3d435661",
X"16703370",
X"982b7098",
X"2c515151",
X"53807324",
X"80fb3860",
X"73291e70",
X"83ffff06",
X"7a228380",
X"80065258",
X"53728380",
X"802e0981",
X"0680de38",
X"60883270",
X"30707207",
X"80256390",
X"32703070",
X"72078025",
X"73075354",
X"58515553",
X"73802ebd",
X"38768706",
X"5372b638",
X"75842976",
X"10057911",
X"84117983",
X"2a575751",
X"53737534",
X"60811634",
X"65861423",
X"66881423",
X"7587387f",
X"8107408d",
X"3975812e",
X"09810685",
X"387f8207",
X"40811670",
X"81ff0657",
X"53817627",
X"fee53863",
X"61291e70",
X"83ffff06",
X"5f538070",
X"4642ff02",
X"840580dd",
X"0534ff0b",
X"993d3483",
X"f539811c",
X"7081ff06",
X"5d538042",
X"73812e09",
X"81068e38",
X"7781800a",
X"2981800a",
X"055880d3",
X"3973802e",
X"89387382",
X"2e098106",
X"8d387c81",
X"800a2981",
X"800a055d",
X"a439815f",
X"83b839ff",
X"1c7081ff",
X"065d537b",
X"63258338",
X"ff437c80",
X"2e92387c",
X"81800a29",
X"81ff0a05",
X"5d7c982c",
X"5d839339",
X"77802e92",
X"38778180",
X"0a2981ff",
X"0a055877",
X"982c5882",
X"fd397753",
X"839e3974",
X"892680f4",
X"38748429",
X"81e59005",
X"53720804",
X"73872e82",
X"e1387385",
X"2e82db38",
X"73882e82",
X"d538738c",
X"2e82cf38",
X"73892e09",
X"81068638",
X"814582c2",
X"3973812e",
X"09810682",
X"b9386280",
X"2582b338",
X"7b982b70",
X"982c5143",
X"82a83973",
X"83ffff06",
X"46829f39",
X"7383ffff",
X"06478296",
X"397381ff",
X"0641828e",
X"3973811a",
X"34828739",
X"7381ff06",
X"4481ff39",
X"7e5382a0",
X"3974812e",
X"81e33874",
X"81248938",
X"74802e8d",
X"3881e739",
X"74822e81",
X"d83881de",
X"3974567b",
X"83388156",
X"74537386",
X"2e098106",
X"97387581",
X"06537280",
X"2e8e3878",
X"2282ffff",
X"06fe8080",
X"0753b639",
X"7b833881",
X"5373822e",
X"09810697",
X"38728106",
X"5372802e",
X"8e387822",
X"81ffff06",
X"81808007",
X"5393397b",
X"9638fc14",
X"53728126",
X"8e387822",
X"ff808007",
X"53727923",
X"80e53980",
X"5573812e",
X"09810683",
X"38735577",
X"5377802e",
X"89387481",
X"06537280",
X"ca3872d0",
X"15545572",
X"81268338",
X"81557780",
X"2eb93874",
X"81065372",
X"802eb038",
X"78228380",
X"80065372",
X"8380802e",
X"0981069f",
X"3873b02e",
X"09810687",
X"3861993d",
X"34913973",
X"b12e0981",
X"06893861",
X"02840580",
X"dd053461",
X"8105538c",
X"39617431",
X"81055384",
X"39611453",
X"7283ffff",
X"064279f7",
X"fb387d83",
X"2a537282",
X"1a347822",
X"83808006",
X"53728380",
X"802e0981",
X"06883881",
X"537f872e",
X"83388053",
X"7283c080",
X"0c993d0d",
X"04fd3d0d",
X"75831133",
X"82123371",
X"982b7190",
X"2b078114",
X"3370882b",
X"72077533",
X"710783c0",
X"800c5253",
X"54565452",
X"853d0d04",
X"f63d0d02",
X"b7053302",
X"8405bb05",
X"33028805",
X"bf05335b",
X"5b5b8058",
X"80577888",
X"2b7a0756",
X"80557a54",
X"8153a352",
X"7c5192c8",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8c3d0d04",
X"f63d0d02",
X"b7053302",
X"8405bb05",
X"33028805",
X"bf05335b",
X"5b5b8058",
X"80577888",
X"2b7a0756",
X"80557a54",
X"8353a352",
X"7c51928c",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8c3d0d04",
X"f73d0d02",
X"b3053302",
X"8405b605",
X"22605a58",
X"56805580",
X"54805381",
X"a3527b51",
X"91de3f83",
X"c0800881",
X"ff0683c0",
X"800c8b3d",
X"0d04ee3d",
X"0d649011",
X"5c5c807b",
X"34800b84",
X"1c0c800b",
X"881c3481",
X"0b891c34",
X"880b8a1c",
X"34800b8b",
X"1c34881b",
X"08c10681",
X"07881c0c",
X"8f3d7054",
X"5d88527b",
X"519c8e3f",
X"83c08008",
X"81ff0670",
X"5b597881",
X"a938903d",
X"335e81db",
X"5a7d892e",
X"09810681",
X"99387c53",
X"92527b51",
X"9be73f83",
X"c0800881",
X"ff06705b",
X"59788182",
X"387c5888",
X"577856a9",
X"55785486",
X"5381a052",
X"7b5190cc",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"80e03802",
X"ba05337b",
X"347c5478",
X"537d527b",
X"519bcf3f",
X"83c08008",
X"81ff0670",
X"5b597880",
X"c13802bd",
X"0533527b",
X"519be73f",
X"83c08008",
X"81ff0670",
X"5b5978aa",
X"38817b33",
X"5a5a7979",
X"26993880",
X"54795388",
X"527b51fd",
X"bb3f811a",
X"7081ff06",
X"7c33525b",
X"59e43981",
X"0b881c34",
X"805a7983",
X"c0800c94",
X"3d0d0480",
X"0b83c080",
X"0c04f93d",
X"0d790284",
X"05ab0533",
X"8e3d7054",
X"585858ff",
X"b7cc3f8a",
X"3d8a0551",
X"ffb7c33f",
X"7551fc8d",
X"3f83c080",
X"08848681",
X"2ebe3883",
X"c0800884",
X"86812699",
X"3883c080",
X"08848280",
X"2e80e638",
X"83c08008",
X"8482812e",
X"9f3881b4",
X"3983c080",
X"0880c082",
X"832e80f4",
X"3883c080",
X"0880c086",
X"832e80e8",
X"38819939",
X"83c0a433",
X"55805674",
X"762e0981",
X"06818b38",
X"74547653",
X"91527751",
X"fbd63f74",
X"54765390",
X"527751fb",
X"cb3f7454",
X"76538452",
X"7751fbfc",
X"3f810b83",
X"c0a43481",
X"b15680de",
X"39805476",
X"53915277",
X"51fba93f",
X"80547653",
X"90527751",
X"fb9e3f80",
X"0b83c0a4",
X"34765287",
X"18335197",
X"923fb539",
X"80547653",
X"94527751",
X"fb823f80",
X"54765390",
X"527751fa",
X"f73f7551",
X"ffb5f73f",
X"83c08008",
X"892a8106",
X"53765287",
X"18335190",
X"c93f800b",
X"83c0a434",
X"80567583",
X"c0800c89",
X"3d0d04f2",
X"3d0d6090",
X"115a5880",
X"0b881a33",
X"71595656",
X"74762e82",
X"a53882ac",
X"3f841908",
X"83c08008",
X"26829538",
X"78335a81",
X"0b8e3d23",
X"903df811",
X"55f40553",
X"99185277",
X"518ae13f",
X"83c08008",
X"81ff0670",
X"57557477",
X"2e098106",
X"81d93886",
X"39745681",
X"d2398156",
X"82578e3d",
X"33770655",
X"74802ebb",
X"38800b8d",
X"3d34903d",
X"f0055484",
X"53755277",
X"51facd3f",
X"83c08008",
X"81ff0655",
X"749d387b",
X"53755277",
X"51fce73f",
X"83c08008",
X"81ff0655",
X"7481b12e",
X"818b3874",
X"ffb33876",
X"1081fc06",
X"81177081",
X"ff065856",
X"57877627",
X"ffa83881",
X"56757a26",
X"80eb3880",
X"0b8d3d34",
X"8c3d7055",
X"57845375",
X"527751f9",
X"f73f83c0",
X"800881ff",
X"06557480",
X"c1387651",
X"ffb3f33f",
X"83c08008",
X"82870655",
X"7482812e",
X"098106aa",
X"3802ae05",
X"33810755",
X"74028405",
X"ae05347b",
X"53755277",
X"51fbeb3f",
X"83c08008",
X"81ff0655",
X"7481b12e",
X"903874fe",
X"b8388116",
X"7081ff06",
X"5755ff91",
X"39805675",
X"81ff0656",
X"973f83c0",
X"80088fd0",
X"05841a0c",
X"75577683",
X"c0800c90",
X"3d0d0404",
X"803d0d90",
X"80a00870",
X"8a2c83c0",
X"800c5182",
X"3d0d0404",
X"83c8e80b",
X"83c0800c",
X"04fd3d0d",
X"75775454",
X"800b83c8",
X"c834728a",
X"38909080",
X"0b84150c",
X"90397281",
X"2e098106",
X"88389098",
X"800b8415",
X"0c841408",
X"83c8e00c",
X"800b8815",
X"0c800b8c",
X"150c83c8",
X"e0085382",
X"0b878014",
X"3487e851",
X"ff92983f",
X"83c8e008",
X"53800b88",
X"143483c8",
X"e0085381",
X"0b878014",
X"3483c8e0",
X"0853800b",
X"8c143483",
X"c8e00853",
X"800ba414",
X"34917434",
X"800b83c0",
X"a834800b",
X"83c0ac34",
X"800b83c0",
X"b0348054",
X"7381c429",
X"83c8ec05",
X"53800b83",
X"14348114",
X"7081ff06",
X"55538774",
X"27e63885",
X"3d0d04fe",
X"3d0d7476",
X"82113370",
X"bf068171",
X"2bff0556",
X"51515253",
X"90712783",
X"38ff5276",
X"51717123",
X"83c8e008",
X"51871333",
X"90123480",
X"0b83c0ac",
X"34800b83",
X"c0b03488",
X"13338a14",
X"33525271",
X"802eaa38",
X"7081ff06",
X"51845270",
X"83387052",
X"7183c0ac",
X"348a1333",
X"70307080",
X"25842b70",
X"88075151",
X"52537083",
X"c0b03490",
X"397081ff",
X"06517083",
X"38985271",
X"83c0b034",
X"800b83c0",
X"800c843d",
X"0d04f13d",
X"0d616568",
X"028c0580",
X"cb053302",
X"900580ce",
X"05220294",
X"0580d605",
X"22424041",
X"5a4040fd",
X"8f3f83c0",
X"8008a788",
X"055b8070",
X"715b5b52",
X"83943983",
X"c8e00851",
X"7d941234",
X"83c0ac33",
X"81075580",
X"7054567f",
X"862680ea",
X"387f8429",
X"81e5c405",
X"83c8e008",
X"53517008",
X"04800b84",
X"1334a139",
X"77337030",
X"70802583",
X"71315151",
X"52537084",
X"13348d39",
X"810b8413",
X"34b83983",
X"0b841334",
X"81705456",
X"ad39810b",
X"841334a2",
X"39773370",
X"30708025",
X"83713151",
X"51525370",
X"84133480",
X"78335252",
X"70833881",
X"52717834",
X"81537488",
X"075583c0",
X"b03383c8",
X"e0085257",
X"810b81d0",
X"123483c8",
X"e0085181",
X"0b819012",
X"347e802e",
X"ae387280",
X"2ea9387e",
X"ff1e5254",
X"7083ffff",
X"06537283",
X"ffff2e97",
X"38737081",
X"05553383",
X"c8e00853",
X"517081c0",
X"1334ff13",
X"51de3983",
X"c8e008a8",
X"11335351",
X"76881234",
X"83c8e008",
X"51747134",
X"81ff5291",
X"3983c8e0",
X"08a01133",
X"70810651",
X"5253708f",
X"38fb813f",
X"7a83c080",
X"0826e638",
X"81883981",
X"0ba01434",
X"83c8e008",
X"a8113380",
X"ff067078",
X"07525351",
X"70802e80",
X"ed387186",
X"2a708106",
X"51517080",
X"2e913880",
X"78335253",
X"70833881",
X"53727834",
X"80e03971",
X"842a7081",
X"06515170",
X"802e9b38",
X"81197083",
X"ffff067d",
X"30709f2a",
X"51525a51",
X"787c2e09",
X"8106af38",
X"a4397183",
X"2a708106",
X"51517080",
X"2e933881",
X"1a7081ff",
X"065b5179",
X"832e0981",
X"0690388a",
X"3971a306",
X"5170802e",
X"85387151",
X"9239f9e8",
X"3f7a83c0",
X"800826fc",
X"e2387181",
X"bf065170",
X"83c0800c",
X"913d0d04",
X"f63d0d02",
X"b3053302",
X"8405b705",
X"33028805",
X"ba052259",
X"5959800b",
X"8c3d348c",
X"3dfc0556",
X"80558054",
X"76537752",
X"7851fbf2",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8c3d0d04",
X"f33d0d7f",
X"6264028c",
X"0580c205",
X"22722281",
X"1533425f",
X"415e5959",
X"8078237d",
X"53783352",
X"8151ffa0",
X"3f83c080",
X"0881ff06",
X"5675802e",
X"86387554",
X"81ad3983",
X"c8e008a8",
X"1133821b",
X"3370862a",
X"70810673",
X"982b5351",
X"575c5657",
X"79802583",
X"38815673",
X"762e8738",
X"81f05481",
X"8239818c",
X"17337081",
X"ff067922",
X"7d713190",
X"2b70902c",
X"7009709f",
X"2c720670",
X"52525351",
X"53575754",
X"75742483",
X"38755574",
X"84808029",
X"fc808005",
X"70902c51",
X"5574ff2e",
X"943883c8",
X"e0088180",
X"11335154",
X"737c7081",
X"055e34db",
X"39772276",
X"05547378",
X"23790970",
X"9f2a7081",
X"06821c33",
X"81bf0671",
X"862b0751",
X"51515473",
X"821a347c",
X"76268a38",
X"7722547a",
X"7426febb",
X"38805473",
X"83c0800c",
X"8f3d0d04",
X"f93d0d7a",
X"57800b89",
X"3d23893d",
X"fc055376",
X"527951f8",
X"da3f83c0",
X"800881ff",
X"06705755",
X"7496387c",
X"547b5388",
X"3d225276",
X"51fde53f",
X"83c08008",
X"81ff0656",
X"7583c080",
X"0c893d0d",
X"04f03d0d",
X"62660288",
X"0580ce05",
X"22415d5e",
X"80028405",
X"80d20522",
X"7f810533",
X"ff115a5d",
X"5a5d81da",
X"5876bf26",
X"80e93878",
X"802e80e1",
X"387a5878",
X"7b278338",
X"7858821e",
X"3370872a",
X"585a7692",
X"3d34923d",
X"fc055677",
X"557b547e",
X"537d3352",
X"8251f8de",
X"3f83c080",
X"0881ff06",
X"5d800b92",
X"3d33585a",
X"76802e83",
X"38815a82",
X"1e3380ff",
X"067a872b",
X"07577682",
X"1f347c91",
X"38787831",
X"7083ffff",
X"06791e5e",
X"5a57ff9b",
X"397c5877",
X"83c0800c",
X"923d0d04",
X"f83d0d7b",
X"028405b2",
X"05225858",
X"800b8a3d",
X"238a3dfc",
X"05537752",
X"7a51f6f7",
X"3f83c080",
X"0881ff06",
X"70575574",
X"96387d54",
X"7653893d",
X"22527751",
X"feaf3f83",
X"c0800881",
X"ff065675",
X"83c0800c",
X"8a3d0d04",
X"ec3d0d66",
X"6e028805",
X"80df0533",
X"028c0580",
X"e3053302",
X"900580e7",
X"05330294",
X"0580eb05",
X"33029805",
X"80ee0522",
X"4143415f",
X"5c405702",
X"80f20522",
X"963d2396",
X"3df00553",
X"84177053",
X"775259f6",
X"863f83c0",
X"800881ff",
X"06587781",
X"e538777a",
X"81800658",
X"40807725",
X"83388140",
X"79943d34",
X"7b028405",
X"80c90534",
X"7c028405",
X"80ca0534",
X"7d028405",
X"80cb0534",
X"7a953d34",
X"7a882a57",
X"76028405",
X"80cd0534",
X"953d2257",
X"76028405",
X"80ce0534",
X"76882a57",
X"76028405",
X"80cf0534",
X"77923d34",
X"963dec11",
X"57578855",
X"f4175492",
X"3d225377",
X"527751f6",
X"953f83c0",
X"800881ff",
X"06587780",
X"ed387e80",
X"2e80cb38",
X"923d2279",
X"0858587f",
X"802e9c38",
X"76818080",
X"07790c7e",
X"54963dfc",
X"05537783",
X"ffff0652",
X"7851f9fc",
X"3f993976",
X"82808007",
X"790c7e54",
X"953d2253",
X"7783ffff",
X"06527851",
X"fc8f3f83",
X"c0800881",
X"ff065877",
X"9d38923d",
X"22538052",
X"7f307080",
X"25847131",
X"535157f9",
X"873f83c0",
X"800881ff",
X"06587783",
X"c0800c96",
X"3d0d04f6",
X"3d0d7c02",
X"8405b705",
X"335b5b80",
X"58805780",
X"56805579",
X"54855380",
X"527a51fd",
X"a33f83c0",
X"800881ff",
X"06597885",
X"3879871c",
X"347883c0",
X"800c8c3d",
X"0d04f93d",
X"0d02a705",
X"33028405",
X"ab053302",
X"8805af05",
X"33585957",
X"800b83c8",
X"ef335454",
X"72742e9f",
X"38811470",
X"81ff0655",
X"53738726",
X"81b63873",
X"81c42983",
X"c8ec0583",
X"11335153",
X"72e33873",
X"81c42983",
X"c8e80555",
X"800b8716",
X"34768816",
X"34758a16",
X"34778916",
X"3480750c",
X"83c8e008",
X"8c160c80",
X"0b841634",
X"880b8516",
X"34800b86",
X"16348415",
X"08ffa1ff",
X"06a08007",
X"84160c81",
X"147081ff",
X"06535374",
X"51febc3f",
X"83c08008",
X"81ff0670",
X"55537280",
X"cd388a39",
X"7308750c",
X"725480c2",
X"397281ea",
X"bc555681",
X"eabc0880",
X"2eb23875",
X"84291470",
X"08765370",
X"08515454",
X"722d83c0",
X"800881ff",
X"06537280",
X"2ece3881",
X"167081ff",
X"0681eabc",
X"71842911",
X"53565753",
X"7208d038",
X"80547383",
X"c0800c89",
X"3d0d04f9",
X"3d0d7957",
X"800b8418",
X"0883c8e0",
X"0c58f08c",
X"3f881708",
X"83c08008",
X"2783ed38",
X"effe3f83",
X"c0800881",
X"0588180c",
X"83c8e008",
X"b8113370",
X"81ff0651",
X"51547381",
X"2ea43873",
X"81248838",
X"73782e8a",
X"38b83973",
X"822e9538",
X"b1397633",
X"81f00654",
X"73902ea6",
X"38917734",
X"a1397358",
X"763381f0",
X"06547390",
X"2e098106",
X"9138efac",
X"3f83c080",
X"0881c805",
X"8c180ca0",
X"77348056",
X"7581c429",
X"83c8ef11",
X"33555573",
X"802eaa38",
X"83c8e815",
X"70085654",
X"74802e9d",
X"38881508",
X"802e9638",
X"8c140883",
X"c8e0082e",
X"09810689",
X"38735188",
X"15085473",
X"2d811670",
X"81ff0657",
X"54877627",
X"ffba3876",
X"335473b0",
X"2e819938",
X"73b0248f",
X"3873912e",
X"ab3873a0",
X"2e80f538",
X"82a63973",
X"80d02e81",
X"e4387380",
X"d0248b38",
X"7380c02e",
X"81993882",
X"8f397381",
X"802e81fb",
X"38828539",
X"80567581",
X"c42983c8",
X"ec118311",
X"33565955",
X"73802ea8",
X"3883c8e8",
X"15700856",
X"5474802e",
X"9b388c14",
X"0883c8e0",
X"082e0981",
X"068e3873",
X"51841508",
X"54732d80",
X"0b831934",
X"81167081",
X"ff065754",
X"877627ff",
X"b9389277",
X"3481b539",
X"edc63f8c",
X"170883c0",
X"80082781",
X"a738b077",
X"3481a139",
X"83c8e008",
X"54800b8c",
X"153483c8",
X"e0085484",
X"0b881534",
X"80c07734",
X"ed9a3f83",
X"c08008b2",
X"058c180c",
X"80fa39ed",
X"8b3f8c17",
X"0883c080",
X"082780ec",
X"3883c8e0",
X"0854810b",
X"8c153483",
X"c8e00854",
X"800b8815",
X"3483c8e0",
X"0854880b",
X"a01534ec",
X"df3f83c0",
X"80089405",
X"8c180c80",
X"d07734bc",
X"3983c8e0",
X"08a01133",
X"70832a70",
X"81065151",
X"55557380",
X"2ea63888",
X"0ba01634",
X"ecb23f8c",
X"170883c0",
X"80082794",
X"38ff8077",
X"348e3977",
X"53805280",
X"51fa8b3f",
X"ff907734",
X"83c8e008",
X"a0113370",
X"832a7081",
X"06515155",
X"5573802e",
X"8638880b",
X"a0163489",
X"3d0d04f4",
X"3d0d02bb",
X"05330284",
X"05bf0533",
X"5d5d800b",
X"83c8ec0b",
X"83c8e80b",
X"8c117271",
X"8814755c",
X"5a5b5f5c",
X"595b5883",
X"15335372",
X"802e8188",
X"38733353",
X"7c732e09",
X"810680fc",
X"38811433",
X"537b732e",
X"09810680",
X"ef387508",
X"83c8e008",
X"2e098106",
X"80e23880",
X"567581c4",
X"2983c8f0",
X"11703383",
X"1e335b57",
X"55537478",
X"2e098106",
X"973883c8",
X"f4130879",
X"082e0981",
X"068a3881",
X"14335274",
X"51fef83f",
X"81167081",
X"ff065753",
X"877627c5",
X"38807708",
X"54547274",
X"2e913876",
X"51841308",
X"53722d83",
X"c0800881",
X"ff065480",
X"0b831b34",
X"7353a939",
X"811881c4",
X"1681c416",
X"81c41981",
X"c41f81c4",
X"1e81c41d",
X"6081c405",
X"415d5e5f",
X"59565658",
X"877825fe",
X"ca388053",
X"7283c080",
X"0c8e3d0d",
X"04f83d0d",
X"02ae0522",
X"7d595780",
X"56815580",
X"54865381",
X"80527a51",
X"f4ee3f83",
X"c0800881",
X"ff0683c0",
X"800c8a3d",
X"0d04f73d",
X"0d02b205",
X"22028405",
X"b7053360",
X"5a5b5780",
X"56825579",
X"54865381",
X"80527b51",
X"f4be3f83",
X"c0800881",
X"ff0683c0",
X"800c8b3d",
X"0d04f83d",
X"0d02af05",
X"33598058",
X"80578056",
X"80557854",
X"89538052",
X"7a51f494",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8a3d0d04",
X"ffb83d0d",
X"80cb3d08",
X"705381e9",
X"885256fe",
X"be9c3f83",
X"c0800880",
X"f3387551",
X"feb8873f",
X"83ffff0b",
X"83c08008",
X"2580e138",
X"7551feb8",
X"863f83c0",
X"80085583",
X"c0800880",
X"cf388280",
X"5383c080",
X"08528a3d",
X"705257fe",
X"fbbf3f74",
X"527551fe",
X"b6f63f80",
X"5980ca3d",
X"fdfc0554",
X"82805376",
X"527551fe",
X"b4fc3f81",
X"15557488",
X"802e0981",
X"06e13880",
X"527551fe",
X"b6ce3f80",
X"0b83d58c",
X"0c7583d5",
X"880c8739",
X"800b83d5",
X"880c80ca",
X"3d0d04ff",
X"3d0d7370",
X"08535102",
X"93053372",
X"34700881",
X"05710c83",
X"3d0d04ff",
X"b83d0d80",
X"cb3d7070",
X"84055208",
X"585683d5",
X"8808802e",
X"80fa388a",
X"3d705a76",
X"55775481",
X"d6bb5380",
X"cb3dfdfc",
X"055255fe",
X"e39a3f80",
X"5280ca3d",
X"fdfc0551",
X"ffad3f83",
X"d58c0852",
X"83d58808",
X"51feb5d4",
X"3f805874",
X"51fee0dc",
X"3f80ca3d",
X"fdf80554",
X"83c08008",
X"53745283",
X"d5880851",
X"feb3cf3f",
X"83d58c08",
X"1883d58c",
X"0c80ca3d",
X"fdf80554",
X"815381e9",
X"945283d5",
X"880851fe",
X"b3b03f83",
X"d58c0818",
X"83d58c0c",
X"80ca3d0d",
X"0483c08c",
X"080283c0",
X"8c0cfd3d",
X"0d805383",
X"c08c088c",
X"05085283",
X"c08c0888",
X"05085183",
X"d43f83c0",
X"80087083",
X"c0800c54",
X"853d0d83",
X"c08c0c04",
X"83c08c08",
X"0283c08c",
X"0cfd3d0d",
X"815383c0",
X"8c088c05",
X"085283c0",
X"8c088805",
X"085183a1",
X"3f83c080",
X"087083c0",
X"800c5485",
X"3d0d83c0",
X"8c0c0483",
X"c08c0802",
X"83c08c0c",
X"f93d0d80",
X"0b83c08c",
X"08fc050c",
X"83c08c08",
X"88050880",
X"25b93883",
X"c08c0888",
X"05083083",
X"c08c0888",
X"050c800b",
X"83c08c08",
X"f4050c83",
X"c08c08fc",
X"05088a38",
X"810b83c0",
X"8c08f405",
X"0c83c08c",
X"08f40508",
X"83c08c08",
X"fc050c83",
X"c08c088c",
X"05088025",
X"b93883c0",
X"8c088c05",
X"083083c0",
X"8c088c05",
X"0c800b83",
X"c08c08f0",
X"050c83c0",
X"8c08fc05",
X"088a3881",
X"0b83c08c",
X"08f0050c",
X"83c08c08",
X"f0050883",
X"c08c08fc",
X"050c8053",
X"83c08c08",
X"8c050852",
X"83c08c08",
X"88050851",
X"81df3f83",
X"c0800870",
X"83c08c08",
X"f8050c54",
X"83c08c08",
X"fc050880",
X"2e903883",
X"c08c08f8",
X"05083083",
X"c08c08f8",
X"050c83c0",
X"8c08f805",
X"087083c0",
X"800c5489",
X"3d0d83c0",
X"8c0c0483",
X"c08c0802",
X"83c08c0c",
X"fb3d0d80",
X"0b83c08c",
X"08fc050c",
X"83c08c08",
X"88050880",
X"25993883",
X"c08c0888",
X"05083083",
X"c08c0888",
X"050c810b",
X"83c08c08",
X"fc050c83",
X"c08c088c",
X"05088025",
X"903883c0",
X"8c088c05",
X"083083c0",
X"8c088c05",
X"0c815383",
X"c08c088c",
X"05085283",
X"c08c0888",
X"050851bd",
X"3f83c080",
X"087083c0",
X"8c08f805",
X"0c5483c0",
X"8c08fc05",
X"08802e90",
X"3883c08c",
X"08f80508",
X"3083c08c",
X"08f8050c",
X"83c08c08",
X"f8050870",
X"83c0800c",
X"54873d0d",
X"83c08c0c",
X"0483c08c",
X"080283c0",
X"8c0cfd3d",
X"0d810b83",
X"c08c08fc",
X"050c800b",
X"83c08c08",
X"f8050c83",
X"c08c088c",
X"050883c0",
X"8c088805",
X"0827b938",
X"83c08c08",
X"fc050880",
X"2eae3880",
X"0b83c08c",
X"088c0508",
X"24a23883",
X"c08c088c",
X"05081083",
X"c08c088c",
X"050c83c0",
X"8c08fc05",
X"081083c0",
X"8c08fc05",
X"0cffb839",
X"83c08c08",
X"fc050880",
X"2e80e138",
X"83c08c08",
X"8c050883",
X"c08c0888",
X"050826ad",
X"3883c08c",
X"08880508",
X"83c08c08",
X"8c050831",
X"83c08c08",
X"88050c83",
X"c08c08f8",
X"050883c0",
X"8c08fc05",
X"080783c0",
X"8c08f805",
X"0c83c08c",
X"08fc0508",
X"812a83c0",
X"8c08fc05",
X"0c83c08c",
X"088c0508",
X"812a83c0",
X"8c088c05",
X"0cff9539",
X"83c08c08",
X"90050880",
X"2e933883",
X"c08c0888",
X"05087083",
X"c08c08f4",
X"050c5191",
X"3983c08c",
X"08f80508",
X"7083c08c",
X"08f4050c",
X"5183c08c",
X"08f40508",
X"83c0800c",
X"853d0d83",
X"c08c0c04",
X"83c08c08",
X"0283c08c",
X"0cff3d0d",
X"800b83c0",
X"8c08fc05",
X"0c83c08c",
X"08880508",
X"8106ff11",
X"70097083",
X"c08c088c",
X"05080683",
X"c08c08fc",
X"05081183",
X"c08c08fc",
X"050c83c0",
X"8c088805",
X"08812a83",
X"c08c0888",
X"050c83c0",
X"8c088c05",
X"081083c0",
X"8c088c05",
X"0c515151",
X"5183c08c",
X"08880508",
X"802e8438",
X"ffab3983",
X"c08c08fc",
X"05087083",
X"c0800c51",
X"833d0d83",
X"c08c0c04",
X"fc3d0d76",
X"70797b55",
X"5555558f",
X"72278c38",
X"72750783",
X"06517080",
X"2ea938ff",
X"125271ff",
X"2e983872",
X"70810554",
X"33747081",
X"055634ff",
X"125271ff",
X"2e098106",
X"ea387483",
X"c0800c86",
X"3d0d0474",
X"51727084",
X"05540871",
X"70840553",
X"0c727084",
X"05540871",
X"70840553",
X"0c727084",
X"05540871",
X"70840553",
X"0c727084",
X"05540871",
X"70840553",
X"0cf01252",
X"718f26c9",
X"38837227",
X"95387270",
X"84055408",
X"71708405",
X"530cfc12",
X"52718326",
X"ed387054",
X"ff813900",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"70704740",
X"0c704268",
X"0c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"000031fa",
X"0000323b",
X"0000325b",
X"0000327f",
X"0000328b",
X"00003295",
X"00003ea8",
X"0000484b",
X"00004914",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3a00",
X"0c0c3b00",
X"0a0a0005",
X"0b0b0005",
X"06060005",
X"07070004",
X"04044500",
X"05054400",
X"0e0f2900",
X"08080004",
X"09090004",
X"0a0f4300",
X"090f4200",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"02010302",
X"02020204",
X"01020800",
X"03800403",
X"20050310",
X"06034007",
X"03010803",
X"02090480",
X"0a05800b",
X"02200c02",
X"100d0240",
X"0e02800f",
X"000057d3",
X"00005ada",
X"000058e6",
X"00005ada",
X"00005923",
X"00005974",
X"000059b3",
X"000059bc",
X"00005ada",
X"00005ada",
X"00005ada",
X"00005ada",
X"000059c5",
X"000059cd",
X"000059d4",
X"00005bda",
X"00005cd3",
X"00005de7",
X"000060d9",
X"000060f4",
X"000060e0",
X"000060f4",
X"000060fb",
X"00006106",
X"0000610d",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"41545800",
X"63686f6f",
X"73652000",
X"66696c65",
X"20202573",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"25782e48",
X"75622e20",
X"25642070",
X"6f727473",
X"00000000",
X"25782e48",
X"49440000",
X"204d6f75",
X"73650000",
X"204b6579",
X"626f6172",
X"64000000",
X"204a6f79",
X"73746963",
X"6b3a2564",
X"00000000",
X"52474200",
X"5343414e",
X"444f5542",
X"4c450000",
X"53564944",
X"454f0000",
X"48444d49",
X"00000000",
X"44564900",
X"56474100",
X"434f4d50",
X"4f534954",
X"45000000",
X"4e545343",
X"00000000",
X"50414c00",
X"73657474",
X"696e6773",
X"00000000",
X"35323030",
X"2e726f6d",
X"00000000",
X"31364b00",
X"556e6b6e",
X"6f776e20",
X"74797065",
X"206f6620",
X"63617274",
X"72696467",
X"65210000",
X"41353200",
X"43415200",
X"42494e00",
X"31366b20",
X"63617274",
X"20747970",
X"65000000",
X"4c656674",
X"20666f72",
X"206f6e65",
X"20636869",
X"70000000",
X"52696768",
X"7420666f",
X"72207477",
X"6f206368",
X"69700000",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a257300",
X"526f7461",
X"74652055",
X"5342206a",
X"6f797374",
X"69636b73",
X"00000000",
X"45786974",
X"00000000",
X"524f4d00",
X"4d454d00",
X"52504400",
X"2f757362",
X"2e6c6f67",
X"00000000",
X"0a000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"00000000",
X"00007368",
X"0000736c",
X"00007378",
X"00007380",
X"00007388",
X"0000738c",
X"00007390",
X"0000739c",
X"000073a4",
X"000072b8",
X"000070d8",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"35323030",
X"00000000",
X"2f617461",
X"72353230",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
