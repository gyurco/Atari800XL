
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f8",
X"80738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80fb",
X"d80c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f2",
X"b02d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580f0c4",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80daa004",
X"fc3d0d76",
X"705255b3",
X"f73f83e0",
X"800815ff",
X"05547375",
X"2e8e3873",
X"335372ae",
X"2e8638ff",
X"1454ef39",
X"77528114",
X"51b38f3f",
X"83e08008",
X"307083e0",
X"80080780",
X"2583e080",
X"0c53863d",
X"0d04fc3d",
X"0d767052",
X"559ab03f",
X"83e08008",
X"54815383",
X"e0800880",
X"c7387451",
X"99f33f83",
X"e080080b",
X"0b80f9e4",
X"5383e080",
X"085253ff",
X"8f3f83e0",
X"8008a538",
X"0b0b80f9",
X"e8527251",
X"fefe3f83",
X"e0800894",
X"380b0b80",
X"f9ec5272",
X"51feed3f",
X"83e08008",
X"802e8338",
X"81547353",
X"7283e080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"99c93f81",
X"5383e080",
X"08993873",
X"5199923f",
X"0b0b80f9",
X"f05283e0",
X"800851fe",
X"b33f83e0",
X"80085372",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"70525499",
X"963f8153",
X"83e08008",
X"99387351",
X"98df3f0b",
X"0b80f9f4",
X"5283e080",
X"0851fe80",
X"3f83e080",
X"08537283",
X"e0800c85",
X"3d0d04e0",
X"3d0da33d",
X"0870525e",
X"8f893f83",
X"e0800833",
X"943d5654",
X"73943880",
X"fefc5274",
X"5184c739",
X"7d527851",
X"92863f84",
X"d1397d51",
X"8ef13f83",
X"e0800852",
X"74518ea1",
X"3f83e09c",
X"0852933d",
X"70525d94",
X"f63f83e0",
X"80085980",
X"0b83e080",
X"08555b83",
X"e080087b",
X"2e943881",
X"1b74525b",
X"97f83f83",
X"e0800854",
X"83e08008",
X"ee38805a",
X"ff7a437a",
X"427a415f",
X"7909709f",
X"2c7b065b",
X"547a7a24",
X"8438ff1b",
X"5af61a70",
X"09709f2c",
X"72067bff",
X"125a5a52",
X"55558075",
X"25953876",
X"5197b73f",
X"83e08008",
X"76ff1858",
X"55577380",
X"24ed3874",
X"7f2e8738",
X"80c3c93f",
X"745f78ff",
X"1b70585d",
X"58807a25",
X"95387751",
X"978c3f83",
X"e0800876",
X"ff185855",
X"58738024",
X"ed38800b",
X"83e7ac0c",
X"800b83e7",
X"cc0c0b0b",
X"80f9f851",
X"8be43f81",
X"800b83e7",
X"cc0c0b0b",
X"80fa8051",
X"8bd43fa8",
X"0b83e7ac",
X"0c76802e",
X"80e83883",
X"e7ac0877",
X"79327030",
X"70720780",
X"2570872b",
X"83e7cc0c",
X"51567853",
X"565696bf",
X"3f83e080",
X"08802e8a",
X"380b0b80",
X"fa88518b",
X"993f7651",
X"95ff3f83",
X"e0800852",
X"0b0b80fb",
X"94518b86",
X"3f765196",
X"853f83e0",
X"800883e7",
X"ac085557",
X"75742586",
X"38a81656",
X"f7397583",
X"e7ac0c86",
X"f07624ff",
X"94388798",
X"0b83e7ac",
X"0c77802e",
X"b7387751",
X"95bb3f83",
X"e0800878",
X"525595db",
X"3f0b0b80",
X"fa905483",
X"e080088f",
X"38873980",
X"7634fd95",
X"390b0b80",
X"fa8c5474",
X"5373520b",
X"0b80f9d8",
X"518a9f3f",
X"80540b0b",
X"80fbd451",
X"8a943f81",
X"145473a8",
X"2e098106",
X"ed38868d",
X"a051bfc8",
X"3f805290",
X"3d705254",
X"80dfe63f",
X"83527351",
X"80dfde3f",
X"61802e80",
X"ff387b54",
X"73ff2e96",
X"3878802e",
X"81803878",
X"5194db3f",
X"83e08008",
X"ff155559",
X"e7397880",
X"2e80eb38",
X"785194d7",
X"3f83e080",
X"08802efc",
X"83387851",
X"949f3f83",
X"e0800852",
X"0b0b80f9",
X"e051abfd",
X"3f83e080",
X"08a4387c",
X"51adb53f",
X"83e08008",
X"5574ff16",
X"56548074",
X"25fbee38",
X"741d7033",
X"555673af",
X"2efec838",
X"e8397851",
X"93dd3f83",
X"e0800852",
X"7c51acec",
X"3ffbce39",
X"7f882960",
X"10057a05",
X"61055afb",
X"ff39a23d",
X"0d04fe3d",
X"0d80fdfc",
X"08703370",
X"81ff0670",
X"842a8132",
X"81065551",
X"52537180",
X"2e8c38a8",
X"733480fd",
X"fc0851b8",
X"71347183",
X"e0800c84",
X"3d0d04fe",
X"3d0d80fd",
X"fc087033",
X"7081ff06",
X"70852a81",
X"32810655",
X"51525371",
X"802e8c38",
X"98733480",
X"fdfc0851",
X"b8713471",
X"83e0800c",
X"843d0d04",
X"803d0d80",
X"fdf80851",
X"93713480",
X"fe840851",
X"ff713482",
X"3d0d04fe",
X"3d0d0293",
X"053380fd",
X"f8085353",
X"8072348a",
X"51bd913f",
X"d33f80fe",
X"88085280",
X"f8723480",
X"fea00852",
X"807234fa",
X"1380fea8",
X"08535372",
X"723480fe",
X"90085280",
X"723480fe",
X"98085272",
X"723480fd",
X"fc085280",
X"723480fd",
X"fc0852b8",
X"7234843d",
X"0d04ff3d",
X"0d028f05",
X"3380fe80",
X"08525271",
X"7134fe9e",
X"3f83e080",
X"08802ef6",
X"38833d0d",
X"04803d0d",
X"853980c5",
X"f53ffeb7",
X"3f83e080",
X"08802ef2",
X"3880fe80",
X"08703370",
X"81ff0683",
X"e0800c51",
X"51823d0d",
X"04803d0d",
X"80fdf808",
X"51a37134",
X"80fe8408",
X"51ff7134",
X"80fdfc08",
X"51a87134",
X"80fdfc08",
X"51b87134",
X"823d0d04",
X"803d0d80",
X"fdf80870",
X"337081c0",
X"06703070",
X"802583e0",
X"800c5151",
X"5151823d",
X"0d04ff3d",
X"0d80fdfc",
X"08703370",
X"81ff0670",
X"832a8132",
X"70810651",
X"51515252",
X"70802ee5",
X"38b07234",
X"80fdfc08",
X"51b87134",
X"833d0d04",
X"803d0d80",
X"feb40870",
X"08810683",
X"e0800c51",
X"823d0d04",
X"fd3d0d75",
X"77545480",
X"73259438",
X"73708105",
X"55335280",
X"fa945185",
X"a13fff13",
X"53e93985",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"80dbbf3f",
X"83e08008",
X"7a27ed38",
X"74802e80",
X"e0387452",
X"755180db",
X"a93f83e0",
X"80087553",
X"76525480",
X"dbcf3f83",
X"e080087a",
X"53755256",
X"80db8f3f",
X"83e08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"e08008c2",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9c",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fbfd3f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd13f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbad3f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83e0900c",
X"7183e094",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383e090",
X"085283e0",
X"940851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"99ba5351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fd3d",
X"0d757052",
X"54a3bd3f",
X"83e08008",
X"14537274",
X"2e9238ff",
X"13703353",
X"5371af2e",
X"098106ee",
X"38811353",
X"7283e080",
X"0c853d0d",
X"04fd3d0d",
X"75777053",
X"5454c73f",
X"83e08008",
X"732ea138",
X"83e08008",
X"733152ff",
X"125271ff",
X"2e8f3872",
X"70810554",
X"33747081",
X"055634eb",
X"39ff1454",
X"80743485",
X"3d0d0480",
X"3d0d7251",
X"ff903f82",
X"3d0d0471",
X"83e0800c",
X"04803d0d",
X"72518071",
X"34810bbc",
X"120c800b",
X"80c0120c",
X"823d0d04",
X"800b83e2",
X"c408248a",
X"38a4a73f",
X"ff0b83e2",
X"c40c800b",
X"83e0800c",
X"04ff3d0d",
X"735283e0",
X"a008722e",
X"8d38d93f",
X"71519692",
X"3f7183e0",
X"a00c833d",
X"0d04f43d",
X"0d7e6062",
X"5c5a5581",
X"54bc1508",
X"81913874",
X"51cf3f79",
X"58807a25",
X"80f73883",
X"e2f40870",
X"892a5783",
X"ff067884",
X"80723156",
X"56577378",
X"25833873",
X"557583e2",
X"c4082e84",
X"38ff893f",
X"83e2c408",
X"8025a638",
X"75892b51",
X"98d53f83",
X"e2f4088f",
X"3dfc1155",
X"5c548152",
X"f81b5196",
X"bf3f7614",
X"83e2f40c",
X"7583e2c4",
X"0c745376",
X"527851a2",
X"d83f83e0",
X"800883e2",
X"f4081683",
X"e2f40c78",
X"7631761b",
X"5b595677",
X"8024ff8b",
X"38617a71",
X"0c547554",
X"75802e83",
X"38815473",
X"83e0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"9b3f7651",
X"feaf3f86",
X"3dfc0553",
X"78527751",
X"95e23f79",
X"75710c54",
X"83e08008",
X"5483e080",
X"08802e83",
X"38815473",
X"83e0800c",
X"863d0d04",
X"fd3d0d76",
X"83e2c408",
X"53538072",
X"24893871",
X"732e8438",
X"fdd63f75",
X"51fdea3f",
X"725197a7",
X"3f735273",
X"802e8338",
X"81527183",
X"e0800c85",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"e0800c51",
X"823d0d04",
X"80c40b83",
X"e0800c04",
X"fd3d0d75",
X"77715470",
X"5355539f",
X"9b3f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfcf13f",
X"735193aa",
X"3f7383e0",
X"a00c83e0",
X"80085383",
X"e0800880",
X"2e833881",
X"537283e0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcc53f",
X"72802ea5",
X"38bc1308",
X"5273519e",
X"a53f83e0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"e0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83e0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83e2c4",
X"0c7483e0",
X"a40c7583",
X"e2c00c9f",
X"923f83e0",
X"800881ff",
X"06528153",
X"71993883",
X"e2dc518e",
X"943f83e0",
X"80085283",
X"e0800880",
X"2e833872",
X"52715372",
X"83e0800c",
X"843d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"519c963f",
X"83e08008",
X"557483e0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"e0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283e2c0",
X"085180ce",
X"cd3f83e0",
X"800857f9",
X"e73f7952",
X"83e2c851",
X"95b43f83",
X"e0800854",
X"805383e0",
X"8008732e",
X"09810682",
X"833883e0",
X"a4080b0b",
X"80f9e053",
X"7052569b",
X"d33f0b0b",
X"80f9e052",
X"80c01651",
X"9bc63f75",
X"bc170c73",
X"82c0170c",
X"810b82c4",
X"170c810b",
X"82c8170c",
X"7382cc17",
X"0cff1782",
X"d0175557",
X"81913983",
X"e0b03370",
X"822a7081",
X"06515455",
X"72818038",
X"74812a81",
X"06587780",
X"f6387484",
X"2a810682",
X"c4150c83",
X"e0b03381",
X"0682c815",
X"0c795273",
X"519aed3f",
X"73519b84",
X"3f83e080",
X"081453af",
X"73708105",
X"553472bc",
X"150c83e0",
X"b1527251",
X"9ace3f83",
X"e0a80882",
X"c0150c83",
X"e0be5280",
X"c014519a",
X"bb3f7880",
X"2e8d3873",
X"51782d83",
X"e0800880",
X"2e993877",
X"82cc150c",
X"75802e86",
X"387382cc",
X"170c7382",
X"d015ff19",
X"59555676",
X"802e9b38",
X"83e0a852",
X"83e2c851",
X"94aa3f83",
X"e080088a",
X"3883e0b1",
X"335372fe",
X"d2387880",
X"2e893883",
X"e0a40851",
X"fcb83f83",
X"e0a40853",
X"7283e080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb53f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f696",
X"3f83e080",
X"08745387",
X"3d705355",
X"55f6b63f",
X"f7963f73",
X"51d33f63",
X"53745283",
X"e0800851",
X"fab83f92",
X"3d0d0471",
X"83e0800c",
X"0480c012",
X"83e0800c",
X"04803d0d",
X"7282c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"e0800c51",
X"823d0d04",
X"f93d0d79",
X"83e09808",
X"57578177",
X"27819638",
X"76881708",
X"27818e38",
X"75335574",
X"822e8938",
X"74832eb3",
X"3880fe39",
X"74547610",
X"83fe0653",
X"76882a8c",
X"17080552",
X"893dfc05",
X"5199c03f",
X"83e08008",
X"80df3802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d13984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"5199903f",
X"83e08008",
X"b038029f",
X"05330284",
X"059e0533",
X"71982b71",
X"902b0702",
X"8c059d05",
X"3370882b",
X"72078d3d",
X"337180ff",
X"fffe8006",
X"07515253",
X"57585683",
X"39815574",
X"83e0800c",
X"893d0d04",
X"fb3d0d83",
X"e09808fe",
X"19881208",
X"fe055556",
X"54805674",
X"73278d38",
X"82143375",
X"71299416",
X"08055753",
X"7583e080",
X"0c873d0d",
X"04fc3d0d",
X"7652800b",
X"83e09808",
X"70335152",
X"5370832e",
X"09810691",
X"38951233",
X"94133371",
X"982b7190",
X"2b075555",
X"519b1233",
X"9a133371",
X"882b0774",
X"0783e080",
X"0c55863d",
X"0d04fc3d",
X"0d7683e0",
X"98085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"fed63f83",
X"e0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183e080",
X"0c863d0d",
X"04fa3d0d",
X"7883e098",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fcb13f",
X"81527183",
X"e0800827",
X"a8388352",
X"83e08008",
X"88170827",
X"9c3883e0",
X"80088c16",
X"0c83e080",
X"0851fdbc",
X"3f83e080",
X"0890160c",
X"73752380",
X"527183e0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585e5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"9f269138",
X"7a51fdd2",
X"3f83e080",
X"0856807d",
X"34838139",
X"933d841c",
X"08705859",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"3880705a",
X"5c887f08",
X"5f5a7b81",
X"1d7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535e57",
X"557480e7",
X"3876ae2e",
X"09810683",
X"38815578",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675bb",
X"3888598b",
X"5affab39",
X"76982b55",
X"74802587",
X"3880f790",
X"173357ff",
X"9f175574",
X"99268938",
X"e0177081",
X"ff065855",
X"78811a70",
X"81ff0672",
X"1b535b57",
X"55767534",
X"fef8397b",
X"1e7f0c80",
X"5576a026",
X"83388155",
X"748b1934",
X"7a51fc82",
X"3f83e080",
X"0880f538",
X"a0547a22",
X"70852b83",
X"e0065455",
X"901b0852",
X"7c5193cb",
X"3f83e080",
X"085783e0",
X"80088181",
X"387c3355",
X"74802e80",
X"f4388b1d",
X"3370832a",
X"70810651",
X"565674b4",
X"388b7d84",
X"1d0883e0",
X"8008595b",
X"5b58ff18",
X"5877ff2e",
X"9a387970",
X"81055b33",
X"79708105",
X"5b337171",
X"31525656",
X"75802ee2",
X"38863975",
X"802e9638",
X"7a51fbe5",
X"3fff8639",
X"83e08008",
X"5683e080",
X"08b63883",
X"39765684",
X"1b088b11",
X"33515574",
X"a7388b1d",
X"3370842a",
X"70810651",
X"56567489",
X"38835694",
X"39815690",
X"397c51fa",
X"943f83e0",
X"8008881c",
X"0cfd8139",
X"7583e080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"5192903f",
X"835683e0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"5191e43f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"765191bb",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583e080",
X"0c8a3d0d",
X"04eb3d0d",
X"675a800b",
X"83e0980c",
X"90dd3f83",
X"e0800881",
X"06558256",
X"7483ee38",
X"7475538f",
X"3d705357",
X"59feca3f",
X"83e08008",
X"81ff0657",
X"76812e09",
X"810680d4",
X"38905483",
X"be537452",
X"755190cf",
X"3f83e080",
X"0880c938",
X"8f3d3355",
X"74802e80",
X"c93802bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"33710770",
X"587b575e",
X"525e5759",
X"57fdee3f",
X"83e08008",
X"81ff0657",
X"76832e09",
X"81068638",
X"815682f1",
X"3976802e",
X"86388656",
X"82e739a4",
X"548d5378",
X"5275518f",
X"e63f8156",
X"83e08008",
X"82d33802",
X"be053302",
X"8405bd05",
X"3371882b",
X"07595d77",
X"ab380280",
X"ce053302",
X"840580cd",
X"05337198",
X"2b71902b",
X"07973d33",
X"70882b72",
X"07029405",
X"80cb0533",
X"71075452",
X"5e575956",
X"02b70533",
X"78712902",
X"8805b605",
X"33028c05",
X"b5053371",
X"882b0770",
X"1d707f8c",
X"050c5f59",
X"57595d8e",
X"3d33821b",
X"3402b905",
X"33903d33",
X"71882b07",
X"5a5c7884",
X"1b2302bb",
X"05330284",
X"05ba0533",
X"71882b07",
X"565c74ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"07515253",
X"575e5c74",
X"76317831",
X"79842a90",
X"3d335471",
X"71315356",
X"56bfb33f",
X"83e08008",
X"82057088",
X"1c0c83e0",
X"8008e08a",
X"05565674",
X"83dffe26",
X"83388257",
X"83fff676",
X"27853883",
X"57893986",
X"5676802e",
X"80db3876",
X"7a347683",
X"2e098106",
X"b0380280",
X"d6053302",
X"840580d5",
X"05337198",
X"2b71902b",
X"07993d33",
X"70882b72",
X"07029405",
X"80d30533",
X"71077f90",
X"050c525e",
X"57585686",
X"39771b90",
X"1b0c841a",
X"228c1b08",
X"1971842a",
X"05941c0c",
X"5d800b81",
X"1b347983",
X"e0980c80",
X"567583e0",
X"800c973d",
X"0d04e93d",
X"0d83e098",
X"08568554",
X"75802e81",
X"8238800b",
X"81173499",
X"3de01146",
X"6a548a3d",
X"705458ec",
X"0551f6e6",
X"3f83e080",
X"085483e0",
X"800880df",
X"38893d33",
X"5473802e",
X"913802ab",
X"05337084",
X"2a810651",
X"5574802e",
X"86388354",
X"80c13976",
X"51f48a3f",
X"83e08008",
X"a0170c02",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"9c1c0c52",
X"78981b0c",
X"53565957",
X"810b8117",
X"34745473",
X"83e0800c",
X"993d0d04",
X"f53d0d7d",
X"7f617283",
X"e098085a",
X"5d5d595c",
X"807b0c85",
X"5775802e",
X"81e03881",
X"16338106",
X"55845774",
X"802e81d2",
X"38913974",
X"81173486",
X"39800b81",
X"17348157",
X"81c0399c",
X"16089817",
X"08315574",
X"78278338",
X"74587780",
X"2e81a938",
X"98160870",
X"83ff0656",
X"577480cf",
X"38821633",
X"ff057789",
X"2a067081",
X"ff065a55",
X"78a03876",
X"8738a016",
X"08558d39",
X"a4160851",
X"f0ea3f83",
X"e0800855",
X"817527ff",
X"a83874a4",
X"170ca416",
X"0851f284",
X"3f83e080",
X"085583e0",
X"8008802e",
X"ff893883",
X"e0800819",
X"a8170c98",
X"160883ff",
X"06848071",
X"31515577",
X"75278338",
X"77557483",
X"ffff0654",
X"98160883",
X"ff0653a8",
X"16085279",
X"577b8338",
X"7b577651",
X"8a8d3f83",
X"e08008fe",
X"d0389816",
X"08159817",
X"0c741a78",
X"76317c08",
X"177d0c59",
X"5afed339",
X"80577683",
X"e0800c8d",
X"3d0d04fa",
X"3d0d7883",
X"e0980855",
X"56855573",
X"802e81e1",
X"38811433",
X"81065384",
X"5572802e",
X"81d3389c",
X"14085372",
X"76278338",
X"72569814",
X"0857800b",
X"98150c75",
X"802e81b7",
X"38821433",
X"70892b56",
X"5376802e",
X"b5387452",
X"ff1651ba",
X"b53f83e0",
X"8008ff18",
X"76547053",
X"5853baa6",
X"3f83e080",
X"08732696",
X"38743070",
X"78067098",
X"170c7771",
X"31a41708",
X"52585153",
X"8939a014",
X"0870a416",
X"0c537476",
X"27b93872",
X"51eed93f",
X"83e08008",
X"53810b83",
X"e0800827",
X"8b388814",
X"0883e080",
X"08268838",
X"800b8115",
X"34b03983",
X"e08008a4",
X"150c9814",
X"08159815",
X"0c757531",
X"56c43998",
X"14081670",
X"98160c73",
X"5256efc8",
X"3f83e080",
X"088c3883",
X"e0800881",
X"15348155",
X"94398214",
X"33ff0576",
X"892a0683",
X"e0800805",
X"a8150c80",
X"557483e0",
X"800c883d",
X"0d04ef3d",
X"0d635685",
X"5583e098",
X"08802e80",
X"d238933d",
X"f4058417",
X"0c645388",
X"3d705376",
X"5257f1d2",
X"3f83e080",
X"085583e0",
X"8008b438",
X"883d3354",
X"73802ea1",
X"3802a705",
X"3370842a",
X"70810651",
X"55558355",
X"73802e97",
X"387651ee",
X"f83f83e0",
X"80088817",
X"0c7551ef",
X"a93f83e0",
X"80085574",
X"83e0800c",
X"933d0d04",
X"e43d0d6e",
X"a13d0840",
X"5e855683",
X"e0980880",
X"2e848538",
X"9e3df405",
X"841f0c7e",
X"98387d51",
X"eef83f83",
X"e0800856",
X"83ee3981",
X"4181f639",
X"834181f1",
X"39933d7f",
X"96054159",
X"807f8295",
X"055e5675",
X"6081ff05",
X"34834190",
X"1e08762e",
X"81d338a0",
X"547d2270",
X"852b83e0",
X"06545890",
X"1e085278",
X"5186983f",
X"83e08008",
X"4183e080",
X"08ffb838",
X"78335c7b",
X"802effb4",
X"388b1933",
X"70bf0671",
X"81065243",
X"5574802e",
X"80de387b",
X"81bf0655",
X"748f2480",
X"d3389a19",
X"33557480",
X"cb38f31d",
X"70585d81",
X"56758b2e",
X"09810685",
X"388e568b",
X"39759a2e",
X"09810683",
X"389c5675",
X"19707081",
X"05523371",
X"33811a82",
X"1a5f5b52",
X"5b557486",
X"38797734",
X"853980df",
X"7734777b",
X"57577aa0",
X"2e098106",
X"c0388156",
X"7b81e532",
X"7030709f",
X"2a515155",
X"7bae2e93",
X"3874802e",
X"8e386183",
X"2a708106",
X"51557480",
X"2e97387d",
X"51ede23f",
X"83e08008",
X"4183e080",
X"08873890",
X"1e08feaf",
X"38806034",
X"75802e88",
X"387c527f",
X"5183a53f",
X"60802e86",
X"38800b90",
X"1f0c6056",
X"60832e85",
X"386081d0",
X"38891f57",
X"901e0880",
X"2e81a838",
X"80567519",
X"70335155",
X"74a02ea0",
X"3874852e",
X"09810684",
X"3881e555",
X"74777081",
X"05593481",
X"167081ff",
X"06575587",
X"7627d738",
X"88193355",
X"74a02ea9",
X"38ae7770",
X"81055934",
X"88567519",
X"70335155",
X"74a02e95",
X"38747770",
X"81055934",
X"81167081",
X"ff065755",
X"8a7627e2",
X"388b1933",
X"7f880534",
X"9f19339e",
X"1a337198",
X"2b71902b",
X"079d1c33",
X"70882b72",
X"079c1e33",
X"7107640c",
X"52991d33",
X"981e3371",
X"882b0753",
X"51535759",
X"56747f84",
X"05239719",
X"33961a33",
X"71882b07",
X"5656747f",
X"86052380",
X"77347d51",
X"ebf33f83",
X"e0800883",
X"32703070",
X"72079f2c",
X"83e08008",
X"06525656",
X"961f3355",
X"748a3889",
X"1f52961f",
X"5181b13f",
X"7583e080",
X"0c9e3d0d",
X"04fd3d0d",
X"75775354",
X"73335170",
X"89387133",
X"5170802e",
X"a1387333",
X"72335253",
X"72712785",
X"38ff5194",
X"39707327",
X"85388151",
X"8b398114",
X"81135354",
X"d3398051",
X"7083e080",
X"0c853d0d",
X"04fd3d0d",
X"75775454",
X"72337081",
X"ff065252",
X"70802ea3",
X"387181ff",
X"068114ff",
X"bf125354",
X"52709926",
X"8938a012",
X"7081ff06",
X"53517174",
X"70810556",
X"34d23980",
X"7434853d",
X"0d04ffbd",
X"3d0d80c6",
X"3d0852a5",
X"3d705254",
X"ffb33f80",
X"c73d0852",
X"853d7052",
X"53ffa63f",
X"72527351",
X"fedf3f80",
X"c53d0d04",
X"fe3d0d74",
X"76535371",
X"70810553",
X"33517073",
X"70810555",
X"3470f038",
X"843d0d04",
X"fe3d0d74",
X"52807233",
X"52537073",
X"2e8d3881",
X"12811471",
X"33535452",
X"70f53872",
X"83e0800c",
X"843d0d04",
X"fc3d0d76",
X"557483e3",
X"88082eaf",
X"38805374",
X"5187cb3f",
X"83e08008",
X"81ff06ff",
X"147081ff",
X"06723070",
X"9f2a5152",
X"55535472",
X"802e8438",
X"71dd3873",
X"fe387483",
X"e3880c86",
X"3d0d04ff",
X"3d0dff0b",
X"83e3880c",
X"84af3f81",
X"51878f3f",
X"83e08008",
X"81ff0652",
X"71ee3881",
X"d63f7183",
X"e0800c83",
X"3d0d04fc",
X"3d0d7602",
X"8405a205",
X"22028805",
X"a605227a",
X"54555555",
X"ff823f72",
X"802ea038",
X"83e39c14",
X"33757081",
X"05573481",
X"147083ff",
X"ff06ff15",
X"7083ffff",
X"06565255",
X"52dd3980",
X"0b83e080",
X"0c863d0d",
X"04fc3d0d",
X"76787a11",
X"56535580",
X"5371742e",
X"93387215",
X"51703383",
X"e39c1334",
X"81128114",
X"5452ea39",
X"800b83e0",
X"800c863d",
X"0d04fd3d",
X"0d905483",
X"e3880851",
X"86fe3f83",
X"e0800881",
X"ff06ff15",
X"71307130",
X"7073079f",
X"2a729f2a",
X"06525552",
X"555372db",
X"38853d0d",
X"04ff3d0d",
X"83e39408",
X"1083e38c",
X"080780fe",
X"b8085271",
X"0c833d0d",
X"04800b83",
X"e3940ce1",
X"3f04810b",
X"83e3940c",
X"d83f04ed",
X"3f047183",
X"e3900c04",
X"803d0d80",
X"51f43f81",
X"0b83e394",
X"0c810b83",
X"e38c0cff",
X"b83f823d",
X"0d04803d",
X"0d723070",
X"74078025",
X"83e38c0c",
X"51ffa23f",
X"823d0d04",
X"fe3d0d02",
X"93053380",
X"febc0854",
X"730c80fe",
X"b8085271",
X"08708106",
X"515170f7",
X"38720870",
X"81ff0683",
X"e0800c51",
X"843d0d04",
X"803d0d81",
X"ff51cd3f",
X"83e08008",
X"81ff0683",
X"e0800c82",
X"3d0d04ff",
X"3d0d7490",
X"2b740780",
X"feac0852",
X"710c833d",
X"0d0404fb",
X"3d0d7802",
X"84059f05",
X"3370982b",
X"55575572",
X"80259b38",
X"7580ff06",
X"56805280",
X"f751e03f",
X"83e08008",
X"81ff0654",
X"73812680",
X"ff388051",
X"fee03fff",
X"9f3f8151",
X"fed83fff",
X"973f7551",
X"fee63f74",
X"982a51fe",
X"df3f7490",
X"2a7081ff",
X"065253fe",
X"d33f7488",
X"2a7081ff",
X"065253fe",
X"c73f7481",
X"ff0651fe",
X"bf3f8155",
X"7580c02e",
X"09810686",
X"38819555",
X"8d397580",
X"c82e0981",
X"06843881",
X"87557451",
X"fe9e3f8a",
X"55fec53f",
X"83e08008",
X"81ff0670",
X"982b5454",
X"7280258c",
X"38ff1570",
X"81ff0656",
X"5374e238",
X"7383e080",
X"0c873d0d",
X"04fa3d0d",
X"fdbe3f80",
X"51fdd33f",
X"8a54fe90",
X"3fff1470",
X"81ff0655",
X"5373f338",
X"73745355",
X"80c051fe",
X"a63f83e0",
X"800881ff",
X"06547381",
X"2e098106",
X"829f3883",
X"aa5280c8",
X"51fe8c3f",
X"83e08008",
X"81ff0653",
X"72812e09",
X"810681a8",
X"38745487",
X"3d741154",
X"56fdc53f",
X"83e08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e53802",
X"9a053353",
X"72812e09",
X"810681d9",
X"38029b05",
X"335380ce",
X"90547281",
X"aa2e8d38",
X"81c73980",
X"e4518afc",
X"3fff1454",
X"73802e81",
X"b838820a",
X"5281e951",
X"fda53f83",
X"e0800881",
X"ff065372",
X"de387252",
X"80fa51fd",
X"923f83e0",
X"800881ff",
X"06537281",
X"90387254",
X"731653fc",
X"d33f83e0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e8",
X"38873d33",
X"70862a70",
X"81065154",
X"548c5572",
X"80e33884",
X"5580de39",
X"745281e9",
X"51fccc3f",
X"83e08008",
X"81ff0653",
X"825581e9",
X"56817327",
X"86387355",
X"80c15680",
X"ce90548a",
X"3980e451",
X"89ee3fff",
X"14547380",
X"2ea93880",
X"527551fc",
X"9a3f83e0",
X"800881ff",
X"065372e1",
X"38848052",
X"80d051fc",
X"863f83e0",
X"800881ff",
X"06537280",
X"2e833880",
X"557483e3",
X"98348051",
X"fb803ffb",
X"bf3f883d",
X"0d04fb3d",
X"0d775480",
X"0b83e398",
X"3370832a",
X"70810651",
X"55575572",
X"752e0981",
X"06853873",
X"892b5473",
X"5280d151",
X"fbbd3f83",
X"e0800881",
X"ff065372",
X"bd3882b8",
X"c054fb80",
X"3f83e080",
X"0881ff06",
X"537281ff",
X"2e098106",
X"8938ff14",
X"5473e738",
X"9f397281",
X"fe2e0981",
X"06963883",
X"e79c5283",
X"e39c51fa",
X"ea3ffad0",
X"3ffacd3f",
X"83398155",
X"8051fa82",
X"3ffac13f",
X"7481ff06",
X"83e0800c",
X"873d0d04",
X"fb3d0d77",
X"83e39c56",
X"548151f9",
X"e53f83e3",
X"98337083",
X"2a708106",
X"51545672",
X"85387389",
X"2b547352",
X"80d851fa",
X"b63f83e0",
X"800881ff",
X"06537280",
X"e43881ff",
X"51f9cd3f",
X"81fe51f9",
X"c73f8480",
X"53747081",
X"05563351",
X"f9ba3fff",
X"137083ff",
X"ff065153",
X"72eb3872",
X"51f9a93f",
X"7251f9a4",
X"3ff9cd3f",
X"83e08008",
X"9f0653a7",
X"88547285",
X"2e8c3899",
X"3980e451",
X"87a63fff",
X"1454f9b0",
X"3f83e080",
X"0881ff2e",
X"843873e9",
X"388051f8",
X"dd3ff99c",
X"3f800b83",
X"e0800c87",
X"3d0d0471",
X"83e7a00c",
X"8880800b",
X"83e79c0c",
X"8480800b",
X"83e7a40c",
X"04f03d0d",
X"80fdc808",
X"54733383",
X"e7a83483",
X"a0805683",
X"e7a00816",
X"83e79c08",
X"17565474",
X"33743483",
X"e7a40816",
X"54807434",
X"81165675",
X"83a0a02e",
X"098106db",
X"3883a480",
X"5683e7a0",
X"081683e7",
X"9c081756",
X"54743374",
X"3483e7a4",
X"08165480",
X"74348116",
X"567583a4",
X"a02e0981",
X"06db3883",
X"a8805683",
X"e7a00816",
X"83e79c08",
X"17565474",
X"33743483",
X"e7a40816",
X"54807434",
X"81165675",
X"83a8902e",
X"098106db",
X"3880fdc8",
X"0854ff74",
X"34805683",
X"e7a00816",
X"83e7a408",
X"17555573",
X"33753481",
X"16567583",
X"a0802e09",
X"8106e438",
X"83b08056",
X"83e7a008",
X"1683e7a4",
X"08175555",
X"73337534",
X"81165675",
X"8480802e",
X"098106e4",
X"3886fd3f",
X"893d58a2",
X"5380f990",
X"527751ad",
X"8c3f8057",
X"8c805683",
X"e7a40816",
X"77195555",
X"73337534",
X"81168118",
X"585676a2",
X"2e098106",
X"e63880fd",
X"ec085486",
X"743480fd",
X"f0085480",
X"743480fd",
X"e8085480",
X"743480fd",
X"d80854af",
X"743480fd",
X"e40854bf",
X"743480fd",
X"e0085480",
X"743480fd",
X"dc08549f",
X"743480fd",
X"d4085480",
X"743480fd",
X"c00854e0",
X"743480fd",
X"b8085476",
X"743480fd",
X"b4085483",
X"743480fd",
X"bc085482",
X"7434923d",
X"0d04fe3d",
X"0d805383",
X"e7a40813",
X"83e7a008",
X"14525270",
X"33723481",
X"13537283",
X"a0802e09",
X"8106e438",
X"83b08053",
X"83e7a408",
X"1383e7a0",
X"08145252",
X"70337234",
X"81135372",
X"8480802e",
X"098106e4",
X"3883a080",
X"5383e7a4",
X"081383e7",
X"a0081452",
X"52703372",
X"34811353",
X"7283a0a0",
X"2e098106",
X"e43883a4",
X"805383e7",
X"a4081383",
X"e7a00814",
X"52527033",
X"72348113",
X"537283a4",
X"a02e0981",
X"06e43883",
X"a8805383",
X"e7a40813",
X"83e7a008",
X"14525270",
X"33723481",
X"13537283",
X"a8902e09",
X"8106e438",
X"80fdc808",
X"5183e7a8",
X"33713484",
X"3d0d0480",
X"3d0d80fe",
X"d0087008",
X"810683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d80fe",
X"d0087008",
X"70fe0676",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80fed008",
X"70087081",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80fed008",
X"700870fd",
X"06761007",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"fed00870",
X"0870822c",
X"bf0683e0",
X"800c5151",
X"823d0d04",
X"ff3d0d80",
X"fed00870",
X"0870fe83",
X"0676822b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80fed008",
X"70087088",
X"2c870683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80fed008",
X"700870f1",
X"ff067688",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d80fed0",
X"08700870",
X"8b2cbf06",
X"83e0800c",
X"5151823d",
X"0d04ff3d",
X"0d80fed0",
X"08700870",
X"f88fff06",
X"768b2b07",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"fee00870",
X"0870882c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fee00870",
X"0870892c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fee00870",
X"08708a2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"fee00870",
X"08708b2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"fd3d0d75",
X"81e62987",
X"2a80fec0",
X"0854730c",
X"853d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d848080",
X"53805288",
X"800a51ff",
X"b33f8180",
X"80538052",
X"82800a51",
X"c63f843d",
X"0d04803d",
X"0d8151fc",
X"ce3f7280",
X"2e8338d2",
X"3f8151fc",
X"f03f8051",
X"fceb3f80",
X"51fcb83f",
X"823d0d04",
X"fd3d0d75",
X"52805480",
X"ff722588",
X"38810bff",
X"80135354",
X"ffbf1251",
X"70992686",
X"38e01252",
X"9e39ff9f",
X"12519971",
X"279538d0",
X"12e01370",
X"54545189",
X"71278838",
X"8f732783",
X"38805273",
X"802e8538",
X"81801252",
X"7181ff06",
X"83e0800c",
X"853d0d04",
X"803d0d84",
X"d8c05180",
X"71708105",
X"53347084",
X"e0c02e09",
X"8106f038",
X"823d0d04",
X"fe3d0d02",
X"97053351",
X"ff863f83",
X"e0800881",
X"ff0683e7",
X"ac085452",
X"8073249b",
X"3883e7c8",
X"08137283",
X"e7cc0807",
X"53537173",
X"3483e7ac",
X"08810583",
X"e7ac0c84",
X"3d0d04fa",
X"3d0d8280",
X"0a1b5580",
X"57883dfc",
X"05547953",
X"74527851",
X"cbaa3f88",
X"3d0d04fe",
X"3d0d83e7",
X"c0085274",
X"51d2883f",
X"83e08008",
X"8c387653",
X"755283e7",
X"c00851c7",
X"3f843d0d",
X"04fe3d0d",
X"83e7c008",
X"53755274",
X"51ccc73f",
X"83e08008",
X"8d387753",
X"765283e7",
X"c00851ff",
X"a23f843d",
X"0d04fe3d",
X"0d83e7c4",
X"0851cbbb",
X"3f83e080",
X"08818080",
X"2e098106",
X"883883c1",
X"8080539b",
X"3983e7c4",
X"0851cb9f",
X"3f83e080",
X"0880d080",
X"2e098106",
X"933883c1",
X"b0805383",
X"e0800852",
X"83e7c408",
X"51fed83f",
X"843d0d04",
X"803d0dfa",
X"cc3f83e0",
X"80088429",
X"80fbe005",
X"700883e0",
X"800c5182",
X"3d0d04ee",
X"3d0d8043",
X"80428041",
X"80705a5b",
X"fdd23f80",
X"0b83e7ac",
X"0c800b83",
X"e7cc0c80",
X"fae051c6",
X"913f8180",
X"0b83e7cc",
X"0c80fae4",
X"51c6833f",
X"80d00b83",
X"e7ac0c78",
X"30707a07",
X"80257087",
X"2b83e7cc",
X"0c5155f9",
X"bb3f83e0",
X"80085280",
X"faec51c5",
X"dd3f80f8",
X"0b83e7ac",
X"0c788132",
X"70307072",
X"07802570",
X"872b83e7",
X"cc0c5156",
X"56fef13f",
X"83e08008",
X"5280faf8",
X"51c5b33f",
X"81a00b83",
X"e7ac0c78",
X"82327030",
X"70720780",
X"2570872b",
X"83e7cc0c",
X"515683e7",
X"c4085256",
X"c6cd3f83",
X"e0800852",
X"80fb8051",
X"c5843f81",
X"f00b83e7",
X"ac0c810b",
X"83e7b05b",
X"5883e7ac",
X"0882197a",
X"32703070",
X"72078025",
X"70872b83",
X"e7cc0c51",
X"578e3d70",
X"55ff1b54",
X"57575798",
X"c93f7970",
X"84055b08",
X"51c6843f",
X"745483e0",
X"80085377",
X"5280fb88",
X"51c4b73f",
X"a81783e7",
X"ac0c8118",
X"5877852e",
X"098106ff",
X"b0388390",
X"0b83e7ac",
X"0c788732",
X"70307072",
X"07802570",
X"872b83e7",
X"cc0c5156",
X"80fb9852",
X"56c4833f",
X"83e00b83",
X"e7ac0c78",
X"88327030",
X"70720780",
X"2570872b",
X"83e7cc0c",
X"515680fb",
X"ac5256c3",
X"e13f868d",
X"a051f9a0",
X"3f805291",
X"3d705255",
X"99bf3f83",
X"52745199",
X"b83f6119",
X"59788025",
X"85388059",
X"90398879",
X"25853888",
X"59873978",
X"882682b1",
X"3878822b",
X"5580f9b4",
X"150804f6",
X"f33f83e0",
X"80086157",
X"5575812e",
X"09810689",
X"3883e080",
X"08105590",
X"3975ff2e",
X"09810688",
X"3883e080",
X"08812c55",
X"90752585",
X"38905588",
X"39748024",
X"83388155",
X"7451f6d0",
X"3f81e639",
X"f6e33f83",
X"e0800861",
X"05557480",
X"25853880",
X"55883987",
X"75258338",
X"87557451",
X"f6df3f81",
X"c4396087",
X"3862802e",
X"81bb388a",
X"dd0b83e0",
X"9c0c83e7",
X"c40851ff",
X"b4d13ffb",
X"8d3f81a5",
X"39605680",
X"76259938",
X"89f60b83",
X"e09c0c83",
X"e7a41570",
X"085255ff",
X"b4b13f74",
X"08529139",
X"75802591",
X"3883e7a4",
X"150851c3",
X"c43f8052",
X"fd1951b8",
X"3962802e",
X"80eb3883",
X"e7a41570",
X"0883e7b0",
X"08720c83",
X"e7b00cfd",
X"1a705351",
X"558adf3f",
X"83e08008",
X"5680518a",
X"d53f83e0",
X"80085274",
X"5186ed3f",
X"75528051",
X"86e63fb5",
X"3962802e",
X"b0388add",
X"0b83e09c",
X"0c83e7c0",
X"0851ffb3",
X"c63f83e7",
X"c00851c2",
X"d23f9c80",
X"0a5380c0",
X"805283e0",
X"800851f9",
X"a63f8155",
X"8c396287",
X"387a802e",
X"fad23880",
X"557483e0",
X"800c943d",
X"0d04fe3d",
X"0df5cd3f",
X"83e08008",
X"802e8638",
X"805180f7",
X"39f5d53f",
X"83e08008",
X"80eb38f5",
X"fb3f83e0",
X"8008802e",
X"aa388151",
X"f3cd3fef",
X"983f800b",
X"83e7ac0c",
X"fa813f83",
X"e0800853",
X"ff0b83e7",
X"ac0cf1ea",
X"3f72be38",
X"7251f3ab",
X"3fbc39f5",
X"af3f83e0",
X"8008802e",
X"b1388151",
X"f3993fee",
X"e43f89f6",
X"0b83e09c",
X"0c83e7b0",
X"0851ffb2",
X"a23fff0b",
X"83e7ac0c",
X"f1b43f83",
X"e7b00852",
X"80518598",
X"3f8151f6",
X"993f843d",
X"0d04fc3d",
X"0d908080",
X"52868480",
X"8051c5a4",
X"3f83e080",
X"0880c338",
X"88e93f80",
X"fee451c9",
X"e43f83e0",
X"800883e7",
X"c4085480",
X"fbb45383",
X"e0800852",
X"55c4bf3f",
X"83e08008",
X"8438f886",
X"3f9c800a",
X"5480c080",
X"5380fbc0",
X"527451f7",
X"d03f8151",
X"f5c03f92",
X"f53f8151",
X"f5b83ffe",
X"913ffc39",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"0283e08c",
X"08fc050c",
X"800b83e7",
X"b00b83e0",
X"8c08f805",
X"0c83e08c",
X"08f4050c",
X"c39e3f83",
X"e0800886",
X"05fc0683",
X"e08c08f0",
X"050c0283",
X"e08c08f0",
X"0508310d",
X"833d7083",
X"e08c08f8",
X"05087084",
X"0583e08c",
X"08f8050c",
X"0c51ffbf",
X"ec3f83e0",
X"8c08f405",
X"08810583",
X"e08c08f4",
X"050c83e0",
X"8c08f405",
X"08862e09",
X"8106ffac",
X"38869480",
X"8051ecbb",
X"3fff0b83",
X"e7ac0c80",
X"0b83e7cc",
X"0c84d8c0",
X"0b83e7c8",
X"0c8151f0",
X"ea3f8151",
X"f1933f80",
X"51f18e3f",
X"8151f1b8",
X"3f8151f2",
X"953f8251",
X"f1df3f80",
X"d0e45280",
X"51ffbdaf",
X"3ffddb3f",
X"83e08c08",
X"fc05080d",
X"800b83e0",
X"800c873d",
X"0d83e08c",
X"0c04803d",
X"0d81ff51",
X"800b83e7",
X"d81234ff",
X"115170f4",
X"38823d0d",
X"04ff3d0d",
X"73703353",
X"51811133",
X"71347181",
X"1234833d",
X"0d04fb3d",
X"0d777956",
X"56807071",
X"55555271",
X"7525ac38",
X"72167033",
X"70147081",
X"ff065551",
X"51517174",
X"27893881",
X"127081ff",
X"06535171",
X"81147083",
X"ffff0655",
X"52547473",
X"24d63871",
X"83e0800c",
X"873d0d04",
X"fd3d0d75",
X"54ffb6d8",
X"3f83e080",
X"08802ef5",
X"3883e9f4",
X"08860570",
X"81ff0652",
X"53ffb4af",
X"3f8439fb",
X"9d3fffb6",
X"b73f83e0",
X"8008812e",
X"f238ffb5",
X"903f83e0",
X"80087434",
X"ffb5863f",
X"83e08008",
X"811534ff",
X"b4fb3f83",
X"e0800882",
X"1534ffb4",
X"f03f83e0",
X"80088315",
X"34ffb4e5",
X"3f83e080",
X"08841534",
X"8439fad6",
X"3fffb5f0",
X"3f83e080",
X"08802ef2",
X"38733383",
X"e7d83481",
X"143383e7",
X"d9348214",
X"3383e7da",
X"34831433",
X"83e7db34",
X"845283e7",
X"d851fe9e",
X"3f83e080",
X"0881ff06",
X"84153355",
X"5372742e",
X"0981068d",
X"38ffb4e0",
X"3f83e080",
X"08802e9a",
X"3883e9f4",
X"08a82e09",
X"81068938",
X"860b83e9",
X"f40c8739",
X"a80b83e9",
X"f40c80e4",
X"51f0993f",
X"853d0d04",
X"f43d0d7e",
X"60595580",
X"5d807582",
X"2b7183e9",
X"f8120c83",
X"ea8c175b",
X"5b577679",
X"3477772e",
X"83b83876",
X"527751ff",
X"be9e3f8e",
X"3dfc0554",
X"905383e9",
X"e0527751",
X"ffbdd93f",
X"7c567590",
X"2e098106",
X"83943883",
X"e9e051fc",
X"f83f83e9",
X"e251fcf1",
X"3f83e9e4",
X"51fcea3f",
X"7683e9f0",
X"0c7751ff",
X"bba53f80",
X"f9e85283",
X"e0800851",
X"ffa9f53f",
X"83e08008",
X"812e0981",
X"0680d438",
X"7683ea88",
X"0c820b83",
X"e9e034ff",
X"960b83e9",
X"e1347751",
X"ffbde43f",
X"83e08008",
X"5583e080",
X"08772588",
X"3883e080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"e9e23474",
X"83e9e334",
X"7683e9e4",
X"34ff800b",
X"83e9e534",
X"81903983",
X"e9e03383",
X"e9e13371",
X"882b0756",
X"5b7483ff",
X"ff2e0981",
X"0680e838",
X"fe800b83",
X"ea880c81",
X"0b83e9f0",
X"0cff0b83",
X"e9e034ff",
X"0b83e9e1",
X"347751ff",
X"bcf13f83",
X"e0800883",
X"ea900c83",
X"e0800855",
X"83e08008",
X"80258838",
X"83e08008",
X"8f055574",
X"842c7083",
X"ffff0670",
X"882a5851",
X"557583e9",
X"e2347483",
X"e9e33476",
X"83e9e434",
X"ff800b83",
X"e9e53481",
X"0b83e9ef",
X"34a53974",
X"85962e09",
X"810680fe",
X"387583ea",
X"880c7751",
X"ffbca53f",
X"83e9ef33",
X"83e08008",
X"07557483",
X"e9ef3483",
X"e9ef3381",
X"06557480",
X"2e833884",
X"5783e9e4",
X"3383e9e5",
X"3371882b",
X"07565c74",
X"81802e09",
X"8106a138",
X"83e9e233",
X"83e9e333",
X"71882b07",
X"565bad80",
X"75278738",
X"76820757",
X"9c397681",
X"07579639",
X"7482802e",
X"09810687",
X"38768307",
X"57873974",
X"81ff268a",
X"387783e9",
X"f81b0c76",
X"79348e3d",
X"0d04803d",
X"0d728429",
X"83e9f805",
X"700883e0",
X"800c5182",
X"3d0d04fe",
X"3d0d800b",
X"83e9dc0c",
X"800b83e9",
X"d80cff0b",
X"83e7d40c",
X"a80b83e9",
X"f40cae51",
X"ffaedc3f",
X"800b83e9",
X"f8545280",
X"73708405",
X"550c8112",
X"5271842e",
X"098106ef",
X"38843d0d",
X"04fe3d0d",
X"74028405",
X"96052253",
X"5371802e",
X"97387270",
X"81055433",
X"51ffaefa",
X"3fff1270",
X"83ffff06",
X"5152e639",
X"843d0d04",
X"fe3d0d02",
X"92052253",
X"82ac51eb",
X"ab3f80c3",
X"51ffaed6",
X"3f819651",
X"eb9e3f72",
X"5283e7d8",
X"51ffb23f",
X"725283e7",
X"d851f8d2",
X"3f83e080",
X"0881ff06",
X"51ffaeb2",
X"3f843d0d",
X"04ffb13d",
X"0d80d13d",
X"f80551f8",
X"fb3f83e9",
X"dc088105",
X"83e9dc0c",
X"80cf3d33",
X"cf117081",
X"ff065156",
X"56748326",
X"88ed3875",
X"8f06ff05",
X"567583e7",
X"d4082e9b",
X"38758326",
X"96387583",
X"e7d40c75",
X"842983e9",
X"f8057008",
X"53557551",
X"fa963f80",
X"762488c9",
X"38758429",
X"83e9f805",
X"55740880",
X"2e88ba38",
X"83e7d408",
X"842983e9",
X"f8057008",
X"02880582",
X"b9053352",
X"5b557480",
X"d22e84b1",
X"387480d2",
X"24903874",
X"bf2e9c38",
X"7480d02e",
X"81d73887",
X"f8397480",
X"d32e80d2",
X"387480d7",
X"2e81c638",
X"87e73902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"5656ffad",
X"b43f80c1",
X"51fface6",
X"3ff6cb3f",
X"860b83e7",
X"d8348152",
X"83e7d851",
X"ffaea13f",
X"8151fde4",
X"3f748938",
X"860b83e9",
X"f40c8739",
X"a80b83e9",
X"f40cffad",
X"803f80c1",
X"51ffacb2",
X"3ff6973f",
X"900b83e9",
X"ef338106",
X"56567480",
X"2e833898",
X"5683e9e4",
X"3383e9e5",
X"3371882b",
X"07565974",
X"81802e09",
X"81069c38",
X"83e9e233",
X"83e9e333",
X"71882b07",
X"5657ad80",
X"75278c38",
X"75818007",
X"56853975",
X"a0075675",
X"83e7d834",
X"ff0b83e7",
X"d934e00b",
X"83e7da34",
X"800b83e7",
X"db348452",
X"83e7d851",
X"ffad953f",
X"8451869e",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055659",
X"ffabf23f",
X"7951ffb6",
X"eb3f83e0",
X"8008802e",
X"8b3880ce",
X"51ffab96",
X"3f85f239",
X"80c151ff",
X"ab8c3fff",
X"ac943fff",
X"aa963f83",
X"ea880858",
X"8375259b",
X"3883e9e4",
X"3383e9e5",
X"3371882b",
X"07fc1771",
X"297a0583",
X"80055a51",
X"578d3974",
X"81802918",
X"ff800558",
X"81805780",
X"5676762e",
X"9338ffaa",
X"e83f83e0",
X"800883e7",
X"d8173481",
X"1656ea39",
X"ffaad63f",
X"83e08008",
X"81ff0677",
X"5383e7d8",
X"5256f4ba",
X"3f83e080",
X"0881ff06",
X"5575752e",
X"09810681",
X"8a38ffaa",
X"d83f80c1",
X"51ffaa8a",
X"3fffab92",
X"3f775279",
X"51ffb580",
X"3f805e80",
X"d13dfdf4",
X"05547653",
X"83e7d852",
X"7951ffb3",
X"8d3f0282",
X"b9053355",
X"81587480",
X"d72e0981",
X"06bd3880",
X"d13dfdf0",
X"05547653",
X"8f3d7053",
X"7a5259ff",
X"b4923f80",
X"5676762e",
X"a2387519",
X"83e7d817",
X"33713370",
X"72327030",
X"70802570",
X"307e0681",
X"1d5d5e51",
X"5151525b",
X"55db3982",
X"ac51e5e4",
X"3f77802e",
X"863880c3",
X"51843980",
X"ce51ffa9",
X"853fffaa",
X"8d3fffa8",
X"8f3f83dd",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055955",
X"80705d59",
X"ffa9a63f",
X"80c151ff",
X"a8d83f83",
X"e9f00879",
X"2e82de38",
X"83ea9008",
X"80fc0555",
X"80fd5274",
X"51868b3f",
X"83e08008",
X"5b778224",
X"b238ff18",
X"70872b83",
X"ffff8006",
X"80fc8005",
X"83e7d859",
X"57558180",
X"55757081",
X"05573377",
X"70810559",
X"34ff1570",
X"81ff0651",
X"5574ea38",
X"828d3977",
X"82e82e81",
X"ab387782",
X"e92e0981",
X"0681b238",
X"80fbd051",
X"ffaef33f",
X"78587787",
X"32703070",
X"72078025",
X"7a8a3270",
X"30707207",
X"80257307",
X"53545a51",
X"57557580",
X"2e973878",
X"78269238",
X"a00b83e7",
X"d81a3481",
X"197081ff",
X"065a55eb",
X"39811870",
X"81ff0659",
X"558a7827",
X"ffbc388f",
X"5883e7d3",
X"183383e7",
X"d81934ff",
X"187081ff",
X"06595577",
X"8426ea38",
X"9058800b",
X"83e7d819",
X"34811870",
X"81ff0670",
X"982b5259",
X"55748025",
X"e93880c6",
X"557a858f",
X"24843880",
X"c2557483",
X"e7d83480",
X"f10b83e7",
X"db34810b",
X"83e7dc34",
X"7a83e7d9",
X"347a882c",
X"557483e7",
X"da3480cb",
X"3982f078",
X"2580c438",
X"7780fd29",
X"fd97d305",
X"527951ff",
X"b1ae3f80",
X"d13dfdec",
X"055480fd",
X"5383e7d8",
X"527951ff",
X"b0e63f7b",
X"81195956",
X"7580fc24",
X"83387858",
X"77882c55",
X"7483e8d5",
X"347783e8",
X"d6347583",
X"e8d73481",
X"805980cc",
X"3983ea88",
X"08578378",
X"259b3883",
X"e9e43383",
X"e9e53371",
X"882b07fc",
X"1a712979",
X"05838005",
X"5951598d",
X"39778180",
X"2917ff80",
X"05578180",
X"59765279",
X"51ffb0bc",
X"3f80d13d",
X"fdec0554",
X"785383e7",
X"d8527951",
X"ffaff53f",
X"7851f6b8",
X"3fffa6aa",
X"3fffa4ac",
X"3f8b3983",
X"e9d80881",
X"0583e9d8",
X"0c80d13d",
X"0d04f6d9",
X"3feb9f3f",
X"f939fc3d",
X"0d767871",
X"842983e9",
X"f8057008",
X"51535353",
X"709e3880",
X"ce723480",
X"cf0b8113",
X"3480ce0b",
X"82133480",
X"c50b8313",
X"34708413",
X"3480e739",
X"83ea8c13",
X"335480d2",
X"72347382",
X"2a708106",
X"515180cf",
X"53708438",
X"80d75372",
X"811334a0",
X"0b821334",
X"73830651",
X"70812e9e",
X"38708124",
X"88387080",
X"2e8f389f",
X"3970822e",
X"92387083",
X"2e923893",
X"3980d855",
X"8e3980d3",
X"55893980",
X"cd558439",
X"80c45574",
X"83133480",
X"c40b8413",
X"34800b85",
X"1334863d",
X"0d04fd3d",
X"0d755480",
X"740c800b",
X"84150c80",
X"0b88150c",
X"80fdcc08",
X"70337081",
X"ff067081",
X"2a813271",
X"81327181",
X"06718106",
X"31841a0c",
X"56567083",
X"2a813271",
X"822a8132",
X"71810671",
X"81063179",
X"0c525551",
X"515180fd",
X"c4087033",
X"70098106",
X"88170c51",
X"51853d0d",
X"04fe3d0d",
X"74765452",
X"7151ff9a",
X"3f72812e",
X"a2388173",
X"268d3872",
X"822eab38",
X"72832e9f",
X"38e63971",
X"08e23884",
X"1208dd38",
X"881208d8",
X"38a03988",
X"1208812e",
X"098106cc",
X"38943988",
X"1208812e",
X"8d387108",
X"89388412",
X"08802eff",
X"b738843d",
X"0d0483e0",
X"8c080283",
X"e08c0cfd",
X"3d0d8053",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"83d43f83",
X"e0800870",
X"83e0800c",
X"54853d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cfd3d",
X"0d815383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"05085183",
X"a13f83e0",
X"80087083",
X"e0800c54",
X"853d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cf93d0d",
X"800b83e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"8025b938",
X"83e08c08",
X"88050830",
X"83e08c08",
X"88050c80",
X"0b83e08c",
X"08f4050c",
X"83e08c08",
X"fc05088a",
X"38810b83",
X"e08c08f4",
X"050c83e0",
X"8c08f405",
X"0883e08c",
X"08fc050c",
X"83e08c08",
X"8c050880",
X"25b93883",
X"e08c088c",
X"05083083",
X"e08c088c",
X"050c800b",
X"83e08c08",
X"f0050c83",
X"e08c08fc",
X"05088a38",
X"810b83e0",
X"8c08f005",
X"0c83e08c",
X"08f00508",
X"83e08c08",
X"fc050c80",
X"5383e08c",
X"088c0508",
X"5283e08c",
X"08880508",
X"5181df3f",
X"83e08008",
X"7083e08c",
X"08f8050c",
X"5483e08c",
X"08fc0508",
X"802e9038",
X"83e08c08",
X"f8050830",
X"83e08c08",
X"f8050c83",
X"e08c08f8",
X"05087083",
X"e0800c54",
X"893d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"800b83e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"80259938",
X"83e08c08",
X"88050830",
X"83e08c08",
X"88050c81",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"8c050880",
X"25903883",
X"e08c088c",
X"05083083",
X"e08c088c",
X"050c8153",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"bd3f83e0",
X"80087083",
X"e08c08f8",
X"050c5483",
X"e08c08fc",
X"0508802e",
X"903883e0",
X"8c08f805",
X"083083e0",
X"8c08f805",
X"0c83e08c",
X"08f80508",
X"7083e080",
X"0c54873d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cfd",
X"3d0d810b",
X"83e08c08",
X"fc050c80",
X"0b83e08c",
X"08f8050c",
X"83e08c08",
X"8c050883",
X"e08c0888",
X"050827b9",
X"3883e08c",
X"08fc0508",
X"802eae38",
X"800b83e0",
X"8c088c05",
X"0824a238",
X"83e08c08",
X"8c050810",
X"83e08c08",
X"8c050c83",
X"e08c08fc",
X"05081083",
X"e08c08fc",
X"050cffb8",
X"3983e08c",
X"08fc0508",
X"802e80e1",
X"3883e08c",
X"088c0508",
X"83e08c08",
X"88050826",
X"ad3883e0",
X"8c088805",
X"0883e08c",
X"088c0508",
X"3183e08c",
X"0888050c",
X"83e08c08",
X"f8050883",
X"e08c08fc",
X"05080783",
X"e08c08f8",
X"050c83e0",
X"8c08fc05",
X"08812a83",
X"e08c08fc",
X"050c83e0",
X"8c088c05",
X"08812a83",
X"e08c088c",
X"050cff95",
X"3983e08c",
X"08900508",
X"802e9338",
X"83e08c08",
X"88050870",
X"83e08c08",
X"f4050c51",
X"913983e0",
X"8c08f805",
X"087083e0",
X"8c08f405",
X"0c5183e0",
X"8c08f405",
X"0883e080",
X"0c853d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cff3d",
X"0d800b83",
X"e08c08fc",
X"050c83e0",
X"8c088805",
X"088106ff",
X"11700970",
X"83e08c08",
X"8c050806",
X"83e08c08",
X"fc050811",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"0508812a",
X"83e08c08",
X"88050c83",
X"e08c088c",
X"05081083",
X"e08c088c",
X"050c5151",
X"515183e0",
X"8c088805",
X"08802e84",
X"38ffab39",
X"83e08c08",
X"fc050870",
X"83e0800c",
X"51833d0d",
X"83e08c0c",
X"04fc3d0d",
X"7670797b",
X"55555555",
X"8f72278c",
X"38727507",
X"83065170",
X"802ea938",
X"ff125271",
X"ff2e9838",
X"72708105",
X"54337470",
X"81055634",
X"ff125271",
X"ff2e0981",
X"06ea3874",
X"83e0800c",
X"863d0d04",
X"74517270",
X"84055408",
X"71708405",
X"530c7270",
X"84055408",
X"71708405",
X"530c7270",
X"84055408",
X"71708405",
X"530c7270",
X"84055408",
X"71708405",
X"530cf012",
X"52718f26",
X"c9388372",
X"27953872",
X"70840554",
X"08717084",
X"05530cfc",
X"12527183",
X"26ed3870",
X"54ff8139",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00002af7",
X"00002b38",
X"00002b5a",
X"00002b79",
X"00002b79",
X"00002b79",
X"00002b79",
X"00002be9",
X"00002c1a",
X"25732025",
X"73000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"524f4d00",
X"42494e00",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"43617274",
X"72696467",
X"6520386b",
X"2073696d",
X"706c6500",
X"45786974",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"6e616d65",
X"20000000",
X"00000000",
X"00000000",
X"00003d1c",
X"00003d20",
X"00003d28",
X"00003d34",
X"00003d40",
X"00003d4c",
X"00003d58",
X"00003d5c",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"0001d20f",
X"0001d400",
X"0001d401",
X"0001d409",
X"0001d010",
X"0001d301",
X"0001d300",
X"0001d20a",
X"0001d01b",
X"0001d016",
X"0001d019",
X"0001d018",
X"0001d017",
X"0001d01a",
X"0001d403",
X"0001d402",
X"0001d40e",
X"0004007c",
X"00040078",
X"00040074",
X"00040068",
X"00040060",
X"0004005c",
X"00040058",
X"00040054",
X"00040050",
X"0004004c",
X"00040048",
X"00040044",
X"00040040",
X"00040034",
X"00040030",
X"0004002c",
X"00040028",
X"00040024",
X"00040020",
X"0004001c",
X"00040018",
X"00040014",
X"00040010",
X"0004000c",
X"00040008",
X"00040004",
X"00040000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"69383030",
X"00000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
