
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81e8",
X"9c738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81f0",
X"dc0c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757580f4",
X"e32d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7580f4a2",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80deb104",
X"fd3d0d75",
X"705254ae",
X"aa3f83c0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"c0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83c0",
X"8008732e",
X"a13883c0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183c0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83c2d008",
X"248a38b4",
X"fb3fff0b",
X"83c2d00c",
X"800b83c0",
X"800c04ff",
X"3d0d7352",
X"83c0ac08",
X"722e8d38",
X"d93f7151",
X"96a03f71",
X"83c0ac0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"55805681",
X"54bc1508",
X"762e0981",
X"06819138",
X"7451c83f",
X"7958757a",
X"2580f738",
X"83c38008",
X"70892a57",
X"83ff0678",
X"84807231",
X"56565773",
X"78258338",
X"73557583",
X"c2d0082e",
X"8438ff82",
X"3f83c2d0",
X"088025a6",
X"3875892b",
X"5198dc3f",
X"83c38008",
X"8f3dfc11",
X"555c5481",
X"52f81b51",
X"96c63f76",
X"1483c380",
X"0c7583c2",
X"d00c7453",
X"76527851",
X"b3a53f83",
X"c0800883",
X"c3800816",
X"83c3800c",
X"78763176",
X"1b5b5956",
X"778024ff",
X"8b38617a",
X"710c5475",
X"5475802e",
X"83388154",
X"7383c080",
X"0c8e3d0d",
X"04fc3d0d",
X"fe943f76",
X"51fea83f",
X"863dfc05",
X"53785277",
X"5195e93f",
X"7975710c",
X"5483c080",
X"085483c0",
X"8008802e",
X"83388154",
X"7383c080",
X"0c863d0d",
X"04fe3d0d",
X"7583c2d0",
X"08535380",
X"72248938",
X"71732e84",
X"38fdcf3f",
X"7451fde3",
X"3f725197",
X"ae3f83c0",
X"80085283",
X"c0800880",
X"2e833881",
X"527183c0",
X"800c843d",
X"0d04803d",
X"0d7280c0",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"3d0d72bc",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"c40b83c0",
X"800c04fd",
X"3d0d7577",
X"71547053",
X"5553a9fb",
X"3f82c813",
X"08bc150c",
X"82c01308",
X"80c0150c",
X"fce43f73",
X"5193ab3f",
X"7383c0ac",
X"0c83c080",
X"085383c0",
X"8008802e",
X"83388153",
X"7283c080",
X"0c853d0d",
X"04fd3d0d",
X"75775553",
X"fcb83f72",
X"802ea538",
X"bc130852",
X"7351a985",
X"3f83c080",
X"088f3877",
X"527251ff",
X"9a3f83c0",
X"8008538a",
X"3982cc13",
X"0853d839",
X"81537283",
X"c0800c85",
X"3d0d04fe",
X"3d0dff0b",
X"83c2d00c",
X"7483c0b0",
X"0c7583c2",
X"cc0cafd9",
X"3f83c080",
X"0881ff06",
X"52815371",
X"993883c2",
X"e8518e94",
X"3f83c080",
X"085283c0",
X"8008802e",
X"83387252",
X"71537283",
X"c0800c84",
X"3d0d04fa",
X"3d0d787a",
X"82c41208",
X"82c41208",
X"70722459",
X"56565757",
X"73732e09",
X"81069138",
X"80c01652",
X"80c01751",
X"a6f63f83",
X"c0800855",
X"7483c080",
X"0c883d0d",
X"04f63d0d",
X"7c5b807b",
X"715c5457",
X"7a772e8c",
X"38811a82",
X"cc140854",
X"5a72f638",
X"805980d9",
X"397a5481",
X"5780707b",
X"7b315a57",
X"55ff1853",
X"74732580",
X"c13882cc",
X"14085273",
X"51ff8c3f",
X"800b83c0",
X"800825a1",
X"3882cc14",
X"0882cc11",
X"0882cc16",
X"0c7482cc",
X"120c5375",
X"802e8638",
X"7282cc17",
X"0c725480",
X"577382cc",
X"15088117",
X"575556ff",
X"b8398119",
X"59800bff",
X"1b545478",
X"73258338",
X"81547681",
X"32707506",
X"515372ff",
X"90388c3d",
X"0d04f73d",
X"0d7b7d5a",
X"5a82d052",
X"83c2cc08",
X"5180e39e",
X"3f83c080",
X"0857f9da",
X"3f795283",
X"c2d45195",
X"b73f83c0",
X"80085480",
X"5383c080",
X"08732e09",
X"81068283",
X"3883c0b0",
X"080b0b81",
X"edbc5370",
X"5256a6b3",
X"3f0b0b81",
X"edbc5280",
X"c01651a6",
X"a63f75bc",
X"170c7382",
X"c0170c81",
X"0b82c417",
X"0c810b82",
X"c8170c73",
X"82cc170c",
X"ff1782d0",
X"17555781",
X"913983c0",
X"bc337082",
X"2a708106",
X"51545572",
X"81803874",
X"812a8106",
X"587780f6",
X"3874842a",
X"810682c4",
X"150c83c0",
X"bc338106",
X"82c8150c",
X"79527351",
X"a5cd3f73",
X"51a5e43f",
X"83c08008",
X"1453af73",
X"70810555",
X"3472bc15",
X"0c83c0bd",
X"527251a5",
X"ae3f83c0",
X"b40882c0",
X"150c83c0",
X"ca5280c0",
X"1451a59b",
X"3f78802e",
X"8d387351",
X"782d83c0",
X"8008802e",
X"99387782",
X"cc150c75",
X"802e8638",
X"7382cc17",
X"0c7382d0",
X"15ff1959",
X"55567680",
X"2e9b3883",
X"c0b45283",
X"c2d45194",
X"ad3f83c0",
X"80088a38",
X"83c0bd33",
X"5372fed2",
X"3878802e",
X"893883c0",
X"b00851fc",
X"b83f83c0",
X"b0085372",
X"83c0800c",
X"8b3d0d04",
X"ff3d0d80",
X"527351fd",
X"b53f833d",
X"0d04f03d",
X"0d627052",
X"54f6893f",
X"83c08008",
X"7453873d",
X"70535555",
X"f6a93ff7",
X"893f7351",
X"d33f6353",
X"745283c0",
X"800851fa",
X"b83f923d",
X"0d047183",
X"c0800c04",
X"80c01283",
X"c0800c04",
X"803d0d72",
X"82c01108",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"7282cc11",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d7282c4",
X"110883c0",
X"800c5182",
X"3d0d04f9",
X"3d0d7983",
X"c0900857",
X"57817727",
X"81963876",
X"88170827",
X"818e3875",
X"33557482",
X"2e893874",
X"832eb338",
X"80fe3974",
X"54761083",
X"fe065376",
X"882a8c17",
X"08055289",
X"3dfc0551",
X"aa873f83",
X"c0800880",
X"df38029d",
X"0533893d",
X"3371882b",
X"07565680",
X"d1398454",
X"76822b83",
X"fc065376",
X"872a8c17",
X"08055289",
X"3dfc0551",
X"a9d73f83",
X"c08008b0",
X"38029f05",
X"33028405",
X"9e053371",
X"982b7190",
X"2b07028c",
X"059d0533",
X"70882b72",
X"078d3d33",
X"7180ffff",
X"fe800607",
X"51525357",
X"58568339",
X"81557483",
X"c0800c89",
X"3d0d04fb",
X"3d0d83c0",
X"9008fe19",
X"881208fe",
X"05555654",
X"80567473",
X"278d3882",
X"14337571",
X"29941608",
X"05575375",
X"83c0800c",
X"873d0d04",
X"fc3d0d76",
X"52800b83",
X"c0900870",
X"33515253",
X"70832e09",
X"81069138",
X"95123394",
X"13337198",
X"2b71902b",
X"07555551",
X"9b12339a",
X"13337188",
X"2b077407",
X"83c0800c",
X"55863d0d",
X"04fc3d0d",
X"7683c090",
X"08555580",
X"75238815",
X"08537281",
X"2e883888",
X"14087326",
X"85388152",
X"b2397290",
X"38733352",
X"71832e09",
X"81068538",
X"90140853",
X"728c160c",
X"72802e8d",
X"387251fe",
X"d63f83c0",
X"80085285",
X"39901408",
X"52719016",
X"0c805271",
X"83c0800c",
X"863d0d04",
X"fa3d0d78",
X"83c09008",
X"71228105",
X"7083ffff",
X"06575457",
X"5573802e",
X"88389015",
X"08537286",
X"38835280",
X"e739738f",
X"06527180",
X"da388113",
X"90160c8c",
X"15085372",
X"9038830b",
X"84172257",
X"52737627",
X"80c638bf",
X"39821633",
X"ff057484",
X"2a065271",
X"b2387251",
X"fcb13f81",
X"527183c0",
X"800827a8",
X"38835283",
X"c0800888",
X"1708279c",
X"3883c080",
X"088c160c",
X"83c08008",
X"51fdbc3f",
X"83c08008",
X"90160c73",
X"75238052",
X"7183c080",
X"0c883d0d",
X"04f23d0d",
X"60626458",
X"5e5b7533",
X"5574a02e",
X"09810688",
X"38811670",
X"4456ef39",
X"62703356",
X"5674af2e",
X"09810684",
X"38811643",
X"800b881c",
X"0c627033",
X"5155749f",
X"2691387a",
X"51fdd23f",
X"83c08008",
X"56807d34",
X"83813993",
X"3d841c08",
X"7058595f",
X"8a55a076",
X"70810558",
X"34ff1555",
X"74ff2e09",
X"8106ef38",
X"80705a5c",
X"887f085f",
X"5a7b811d",
X"7081ff06",
X"60137033",
X"70af3270",
X"30a07327",
X"71802507",
X"5151525b",
X"535e5755",
X"7480e738",
X"76ae2e09",
X"81068338",
X"8155787a",
X"27750755",
X"74802e9f",
X"38798832",
X"703078ae",
X"32703070",
X"73079f2a",
X"53515751",
X"5675bb38",
X"88598b5a",
X"ffab3976",
X"982b5574",
X"80258738",
X"81e7ac17",
X"3357ff9f",
X"17557499",
X"268938e0",
X"177081ff",
X"06585578",
X"811a7081",
X"ff06721b",
X"535b5755",
X"767534fe",
X"f8397b1e",
X"7f0c8055",
X"76a02683",
X"38815574",
X"8b19347a",
X"51fc823f",
X"83c08008",
X"80f538a0",
X"547a2270",
X"852b83e0",
X"06545590",
X"1b08527c",
X"51a4923f",
X"83c08008",
X"5783c080",
X"08818138",
X"7c335574",
X"802e80f4",
X"388b1d33",
X"70832a70",
X"81065156",
X"5674b438",
X"8b7d841d",
X"0883c080",
X"08595b5b",
X"58ff1858",
X"77ff2e9a",
X"38797081",
X"055b3379",
X"7081055b",
X"33717131",
X"52565675",
X"802ee238",
X"86397580",
X"2e96387a",
X"51fbe53f",
X"ff863983",
X"c0800856",
X"83c08008",
X"b6388339",
X"7656841b",
X"088b1133",
X"515574a7",
X"388b1d33",
X"70842a70",
X"81065156",
X"56748938",
X"83569439",
X"81569039",
X"7c51fa94",
X"3f83c080",
X"08881c0c",
X"fd813975",
X"83c0800c",
X"903d0d04",
X"f83d0d7a",
X"7c595782",
X"5483fe53",
X"77527651",
X"a2d73f83",
X"5683c080",
X"0880ec38",
X"81173377",
X"3371882b",
X"07565682",
X"567482d4",
X"d52e0981",
X"0680d438",
X"7554b653",
X"77527651",
X"a2ab3f83",
X"c0800898",
X"38811733",
X"77337188",
X"2b0783c0",
X"80085256",
X"56748182",
X"c62eac38",
X"825480d2",
X"53775276",
X"51a2823f",
X"83c08008",
X"98388117",
X"33773371",
X"882b0783",
X"c0800852",
X"56567481",
X"82c62e83",
X"38815675",
X"83c0800c",
X"8a3d0d04",
X"eb3d0d67",
X"5a800b83",
X"c0900ca1",
X"a43f83c0",
X"80088106",
X"55825674",
X"83ef3874",
X"75538f3d",
X"70535759",
X"feca3f83",
X"c0800881",
X"ff065776",
X"812e0981",
X"0680d438",
X"905483be",
X"53745275",
X"51a1963f",
X"83c08008",
X"80c9388f",
X"3d335574",
X"802e80c9",
X"3802bf05",
X"33028405",
X"be053371",
X"982b7190",
X"2b07028c",
X"05bd0533",
X"70882b72",
X"07953d33",
X"71077058",
X"7b575e52",
X"5e575957",
X"fdee3f83",
X"c0800881",
X"ff065776",
X"832e0981",
X"06863881",
X"5682f239",
X"76802e86",
X"38865682",
X"e839a454",
X"8d537852",
X"7551a0ad",
X"3f815683",
X"c0800882",
X"d43802be",
X"05330284",
X"05bd0533",
X"71882b07",
X"595d77ab",
X"380280ce",
X"05330284",
X"0580cd05",
X"3371982b",
X"71902b07",
X"973d3370",
X"882b7207",
X"02940580",
X"cb053371",
X"0754525e",
X"57595602",
X"b7053378",
X"71290288",
X"05b60533",
X"028c05b5",
X"05337188",
X"2b07701d",
X"707f8c05",
X"0c5f5957",
X"595d8e3d",
X"33821b34",
X"02b90533",
X"903d3371",
X"882b075a",
X"5c78841b",
X"2302bb05",
X"33028405",
X"ba053371",
X"882b0756",
X"5c74ab38",
X"0280ca05",
X"33028405",
X"80c90533",
X"71982b71",
X"902b0796",
X"3d337088",
X"2b720702",
X"940580c7",
X"05337107",
X"51525357",
X"5e5c7476",
X"31783179",
X"842a903d",
X"33547171",
X"31535656",
X"80d4833f",
X"83c08008",
X"82057088",
X"1c0c83c0",
X"8008e08a",
X"05565674",
X"83dffe26",
X"83388257",
X"83fff676",
X"27853883",
X"57893986",
X"5676802e",
X"80db3876",
X"7a347683",
X"2e098106",
X"b0380280",
X"d6053302",
X"840580d5",
X"05337198",
X"2b71902b",
X"07993d33",
X"70882b72",
X"07029405",
X"80d30533",
X"71077f90",
X"050c525e",
X"57585686",
X"39771b90",
X"1b0c841a",
X"228c1b08",
X"1971842a",
X"05941c0c",
X"5d800b81",
X"1b347983",
X"c0900c80",
X"567583c0",
X"800c973d",
X"0d04e93d",
X"0d83c090",
X"08568554",
X"75802e81",
X"8238800b",
X"81173499",
X"3de01146",
X"6a548a3d",
X"705458ec",
X"0551f6e5",
X"3f83c080",
X"085483c0",
X"800880df",
X"38893d33",
X"5473802e",
X"913802ab",
X"05337084",
X"2a810651",
X"5574802e",
X"86388354",
X"80c13976",
X"51f4893f",
X"83c08008",
X"a0170c02",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"9c1c0c52",
X"78981b0c",
X"53565957",
X"810b8117",
X"34745473",
X"83c0800c",
X"993d0d04",
X"f53d0d7d",
X"7f617283",
X"c090085a",
X"5d5d595c",
X"807b0c85",
X"5775802e",
X"81e03881",
X"16338106",
X"55845774",
X"802e81d2",
X"38913974",
X"81173486",
X"39800b81",
X"17348157",
X"81c0399c",
X"16089817",
X"08315574",
X"78278338",
X"74587780",
X"2e81a938",
X"98160870",
X"83ff0656",
X"577480cf",
X"38821633",
X"ff057789",
X"2a067081",
X"ff065a55",
X"78a03876",
X"8738a016",
X"08558d39",
X"a4160851",
X"f0e93f83",
X"c0800855",
X"817527ff",
X"a83874a4",
X"170ca416",
X"0851f283",
X"3f83c080",
X"085583c0",
X"8008802e",
X"ff893883",
X"c0800819",
X"a8170c98",
X"160883ff",
X"06848071",
X"31515577",
X"75278338",
X"77557483",
X"ffff0654",
X"98160883",
X"ff0653a8",
X"16085279",
X"577b8338",
X"7b577651",
X"9ad33f83",
X"c08008fe",
X"d0389816",
X"08159817",
X"0c741a78",
X"76317c08",
X"177d0c59",
X"5afed339",
X"80577683",
X"c0800c8d",
X"3d0d04fa",
X"3d0d7883",
X"c0900855",
X"56855573",
X"802e81e3",
X"38811433",
X"81065384",
X"5572802e",
X"81d5389c",
X"14085372",
X"76278338",
X"72569814",
X"0857800b",
X"98150c75",
X"802e81b9",
X"38821433",
X"70892b56",
X"5376802e",
X"b7387452",
X"ff165180",
X"cf843f83",
X"c08008ff",
X"18765470",
X"53585380",
X"cef43f83",
X"c0800873",
X"26963874",
X"30707806",
X"7098170c",
X"777131a4",
X"17085258",
X"51538939",
X"a0140870",
X"a4160c53",
X"747627b9",
X"387251ee",
X"d63f83c0",
X"80085381",
X"0b83c080",
X"08278b38",
X"88140883",
X"c0800826",
X"8838800b",
X"811534b0",
X"3983c080",
X"08a4150c",
X"98140815",
X"98150c75",
X"753156c4",
X"39981408",
X"16709816",
X"0c735256",
X"efc53f83",
X"c080088c",
X"3883c080",
X"08811534",
X"81559439",
X"821433ff",
X"0576892a",
X"0683c080",
X"0805a815",
X"0c805574",
X"83c0800c",
X"883d0d04",
X"ef3d0d63",
X"56855583",
X"c0900880",
X"2e80d238",
X"933df405",
X"84170c64",
X"53883d70",
X"53765257",
X"f1cf3f83",
X"c0800855",
X"83c08008",
X"b438883d",
X"33547380",
X"2ea13802",
X"a7053370",
X"842a7081",
X"06515555",
X"83557380",
X"2e973876",
X"51eef53f",
X"83c08008",
X"88170c75",
X"51efa63f",
X"83c08008",
X"557483c0",
X"800c933d",
X"0d04e43d",
X"0d6ea13d",
X"08405e85",
X"5683c090",
X"08802e84",
X"85389e3d",
X"f405841f",
X"0c7e9838",
X"7d51eef5",
X"3f83c080",
X"085683ee",
X"39814181",
X"f6398341",
X"81f13993",
X"3d7f9605",
X"4159807f",
X"8295055e",
X"56756081",
X"ff053483",
X"41901e08",
X"762e81d3",
X"38a0547d",
X"2270852b",
X"83e00654",
X"58901e08",
X"52785196",
X"dc3f83c0",
X"80084183",
X"c08008ff",
X"b8387833",
X"5c7b802e",
X"ffb4388b",
X"193370bf",
X"06718106",
X"52435574",
X"802e80de",
X"387b81bf",
X"0655748f",
X"2480d338",
X"9a193355",
X"7480cb38",
X"f31d7058",
X"5d815675",
X"8b2e0981",
X"0685388e",
X"568b3975",
X"9a2e0981",
X"0683389c",
X"56751970",
X"70810552",
X"33713381",
X"1a821a5f",
X"5b525b55",
X"74863879",
X"77348539",
X"80df7734",
X"777b5757",
X"7aa02e09",
X"8106c038",
X"81567b81",
X"e5327030",
X"709f2a51",
X"51557bae",
X"2e933874",
X"802e8e38",
X"61832a70",
X"81065155",
X"74802e97",
X"387d51ed",
X"df3f83c0",
X"80084183",
X"c0800887",
X"38901e08",
X"feaf3880",
X"60347580",
X"2e88387c",
X"527f518e",
X"823f6080",
X"2e863880",
X"0b901f0c",
X"60566083",
X"2e853860",
X"81d03889",
X"1f57901e",
X"08802e81",
X"a8388056",
X"75197033",
X"515574a0",
X"2ea03874",
X"852e0981",
X"06843881",
X"e5557477",
X"70810559",
X"34811670",
X"81ff0657",
X"55877627",
X"d7388819",
X"335574a0",
X"2ea938ae",
X"77708105",
X"59348856",
X"75197033",
X"515574a0",
X"2e953874",
X"77708105",
X"59348116",
X"7081ff06",
X"57558a76",
X"27e2388b",
X"19337f88",
X"05349f19",
X"339e1a33",
X"71982b71",
X"902b079d",
X"1c337088",
X"2b72079c",
X"1e337107",
X"640c5299",
X"1d33981e",
X"3371882b",
X"07535153",
X"57595674",
X"7f840523",
X"97193396",
X"1a337188",
X"2b075656",
X"747f8605",
X"23807734",
X"7d51ebf0",
X"3f83c080",
X"08833270",
X"30707207",
X"9f2c83c0",
X"80080652",
X"5656961f",
X"3355748a",
X"38891f52",
X"961f518c",
X"8e3f7583",
X"c0800c9e",
X"3d0d04f4",
X"3d0d7e8f",
X"3dec1156",
X"56589053",
X"f0155277",
X"51e0d23f",
X"83c08008",
X"80d63878",
X"902e0981",
X"0680cd38",
X"02ab0533",
X"81f0e40b",
X"81f0e433",
X"5758568c",
X"3974762e",
X"8a388417",
X"70335657",
X"74f33876",
X"33705755",
X"74802eac",
X"38821722",
X"708a2b90",
X"3dec0556",
X"70555656",
X"96800a52",
X"7751e081",
X"3f83c080",
X"08863878",
X"752e8538",
X"80568539",
X"81173356",
X"7583c080",
X"0c8e3d0d",
X"04fc3d0d",
X"76705255",
X"8b953f83",
X"c0800815",
X"ff055473",
X"752e8e38",
X"73335372",
X"ae2e8638",
X"ff1454ef",
X"39775281",
X"14518aad",
X"3f83c080",
X"08307083",
X"c0800807",
X"802583c0",
X"800c5386",
X"3d0d04fc",
X"3d0d7670",
X"5255e6ee",
X"3f83c080",
X"08548153",
X"83c08008",
X"80c13874",
X"51e6b13f",
X"83c08008",
X"81edcc53",
X"83c08008",
X"5253ff91",
X"3f83c080",
X"08a13881",
X"edd05272",
X"51ff823f",
X"83c08008",
X"923881ed",
X"d4527251",
X"fef33f83",
X"c0800880",
X"2e833881",
X"54735372",
X"83c0800c",
X"863d0d04",
X"fd3d0d75",
X"705254e6",
X"8d3f8153",
X"83c08008",
X"98387351",
X"e5d63f83",
X"c3980852",
X"83c08008",
X"51feba3f",
X"83c08008",
X"537283c0",
X"800c853d",
X"0d04df3d",
X"0da43d08",
X"70525edb",
X"f43f83c0",
X"80083395",
X"3d565473",
X"963881f4",
X"b4527451",
X"898d3f9a",
X"397d5278",
X"51defc3f",
X"84d0397d",
X"51dbda3f",
X"83c08008",
X"527451db",
X"8a3f8043",
X"80428041",
X"804083c3",
X"a0085294",
X"3d70525d",
X"e1e43f83",
X"c0800859",
X"800b83c0",
X"8008555b",
X"83c08008",
X"7b2e9438",
X"811b7452",
X"5be4e63f",
X"83c08008",
X"5483c080",
X"08ee3880",
X"5aff5f79",
X"09709f2c",
X"7b065b54",
X"7a7a2484",
X"38ff1b5a",
X"f61a7009",
X"709f2c72",
X"067bff12",
X"5a5a5255",
X"55807525",
X"95387651",
X"e4ab3f83",
X"c0800876",
X"ff185855",
X"57738024",
X"ed38747f",
X"2e8638a1",
X"b53f745f",
X"78ff1b70",
X"585d5880",
X"7a259538",
X"7751e481",
X"3f83c080",
X"0876ff18",
X"58555873",
X"8024ed38",
X"800b83c7",
X"d00c800b",
X"83c8980c",
X"81edd851",
X"8d8c3f81",
X"800b83c8",
X"980c81ed",
X"e0518cfe",
X"3fa80b83",
X"c7d00c76",
X"802e80e4",
X"3883c7d0",
X"08777932",
X"70307072",
X"07802570",
X"872b83c8",
X"980c5156",
X"78535656",
X"e3b83f83",
X"c0800880",
X"2e883881",
X"ede8518c",
X"c53f7651",
X"e2fa3f83",
X"c0800852",
X"81ef8851",
X"8cb43f76",
X"51e3823f",
X"83c08008",
X"83c7d008",
X"55577574",
X"258638a8",
X"1656f739",
X"7583c7d0",
X"0c86f076",
X"24ff9838",
X"87980b83",
X"c7d00c77",
X"802eb138",
X"7751e2b8",
X"3f83c080",
X"08785255",
X"e2d83f81",
X"edf05483",
X"c080088d",
X"38873980",
X"763481d0",
X"3981edec",
X"54745373",
X"5281edc0",
X"518bd33f",
X"805481ed",
X"c8518bca",
X"3f811454",
X"73a82e09",
X"8106ef38",
X"868da051",
X"9da83f80",
X"52903d70",
X"525780c4",
X"f93f8352",
X"765180c4",
X"f13f6281",
X"8f386180",
X"2e80fb38",
X"7b5473ff",
X"2e963878",
X"802e818a",
X"387851e1",
X"dc3f83c0",
X"8008ff15",
X"5559e739",
X"78802e80",
X"f5387851",
X"e1d83f83",
X"c0800880",
X"2efc8e38",
X"7851e1a0",
X"3f83c080",
X"085281ed",
X"bc5183e0",
X"3f83c080",
X"08a3387c",
X"5185983f",
X"83c08008",
X"5574ff16",
X"56548074",
X"25ae3874",
X"1d703355",
X"5673af2e",
X"fecd38e9",
X"397851e0",
X"e13f83c0",
X"8008527c",
X"5184d03f",
X"8f397f88",
X"29601005",
X"7a056105",
X"5afc9039",
X"62802efb",
X"d1388052",
X"765180c3",
X"d13fa33d",
X"0d04803d",
X"0d9088b8",
X"337081ff",
X"0670842a",
X"81327081",
X"06515151",
X"5170802e",
X"8d38a80b",
X"9088b834",
X"b80b9088",
X"b8347083",
X"c0800c82",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067085",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d3898",
X"0b9088b8",
X"34b80b90",
X"88b83470",
X"83c0800c",
X"823d0d04",
X"930b9088",
X"bc34ff0b",
X"9088a834",
X"04ff3d0d",
X"028f0533",
X"52800b90",
X"88bc348a",
X"519aef3f",
X"df3f80f8",
X"0b9088a0",
X"34800b90",
X"888834fa",
X"12527190",
X"88803480",
X"0b908898",
X"34719088",
X"90349088",
X"b8528072",
X"34b87234",
X"833d0d04",
X"803d0d02",
X"8b053351",
X"709088b4",
X"34febf3f",
X"83c08008",
X"802ef638",
X"823d0d04",
X"803d0d84",
X"39a6af3f",
X"fed93f83",
X"c0800880",
X"2ef33890",
X"88b43370",
X"81ff0683",
X"c0800c51",
X"823d0d04",
X"803d0da3",
X"0b9088bc",
X"34ff0b90",
X"88a83490",
X"88b851a8",
X"7134b871",
X"34823d0d",
X"04803d0d",
X"9088bc33",
X"70982b70",
X"802583c0",
X"800c5151",
X"823d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"832a8132",
X"70810651",
X"51515170",
X"802ee838",
X"b00b9088",
X"b834b80b",
X"9088b834",
X"823d0d04",
X"803d0d90",
X"80ac0881",
X"0683c080",
X"0c823d0d",
X"04fd3d0d",
X"75775454",
X"80732594",
X"38737081",
X"05553352",
X"81edf451",
X"87843fff",
X"1353e939",
X"853d0d04",
X"fd3d0d75",
X"77535473",
X"33517089",
X"38713351",
X"70802ea1",
X"38733372",
X"33525372",
X"71278538",
X"ff519439",
X"70732785",
X"3881518b",
X"39811481",
X"135354d3",
X"39805170",
X"83c0800c",
X"853d0d04",
X"fd3d0d75",
X"77545472",
X"337081ff",
X"06525270",
X"802ea338",
X"7181ff06",
X"8114ffbf",
X"12535452",
X"70992689",
X"38a01270",
X"81ff0653",
X"51717470",
X"81055634",
X"d2398074",
X"34853d0d",
X"04ffbd3d",
X"0d80c63d",
X"0852a53d",
X"705254ff",
X"b33f80c7",
X"3d085285",
X"3d705253",
X"ffa63f72",
X"527351fe",
X"df3f80c5",
X"3d0d04fe",
X"3d0d7476",
X"53537170",
X"81055333",
X"51707370",
X"81055534",
X"70f03884",
X"3d0d04fe",
X"3d0d7452",
X"80723352",
X"5370732e",
X"8d388112",
X"81147133",
X"53545270",
X"f5387283",
X"c0800c84",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"bbdc3f83",
X"c080087a",
X"27ee3874",
X"802e80dd",
X"38745275",
X"51bbc73f",
X"83c08008",
X"75537652",
X"54bbcb3f",
X"83c08008",
X"7a537552",
X"56bbaf3f",
X"83c08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"c08008c5",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9f",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fc813f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd53f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbb13f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83c0940c",
X"7183c098",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383c094",
X"085283c0",
X"980851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"bdbe5351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fc3d",
X"0d765574",
X"83c3ac08",
X"2eaf3880",
X"53745187",
X"c13f83c0",
X"800881ff",
X"06ff1470",
X"81ff0672",
X"30709f2a",
X"51525553",
X"5472802e",
X"843871dd",
X"3873fe38",
X"7483c3ac",
X"0c863d0d",
X"04ff3d0d",
X"ff0b83c3",
X"ac0c84a5",
X"3f815187",
X"853f83c0",
X"800881ff",
X"065271ee",
X"3881d33f",
X"7183c080",
X"0c833d0d",
X"04fc3d0d",
X"76028405",
X"a2052202",
X"8805a605",
X"227a5455",
X"5555ff82",
X"3f72802e",
X"a03883c3",
X"c0143375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552dd",
X"39800b83",
X"c0800c86",
X"3d0d04fc",
X"3d0d7678",
X"7a115653",
X"55805371",
X"742e9338",
X"72155170",
X"3383c3c0",
X"13348112",
X"81145452",
X"ea39800b",
X"83c0800c",
X"863d0d04",
X"fd3d0d90",
X"5483c3ac",
X"085186f4",
X"3f83c080",
X"0881ff06",
X"ff157130",
X"71307073",
X"079f2a72",
X"9f2a0652",
X"55525553",
X"72db3885",
X"3d0d0480",
X"3d0d83c3",
X"b8081083",
X"c3b00807",
X"9080a80c",
X"823d0d04",
X"800b83c3",
X"b80ce43f",
X"04810b83",
X"c3b80cdb",
X"3f04ed3f",
X"047183c3",
X"b40c0480",
X"3d0d8051",
X"f43f810b",
X"83c3b80c",
X"810b83c3",
X"b00cffbb",
X"3f823d0d",
X"04803d0d",
X"72307074",
X"07802583",
X"c3b00c51",
X"ffa53f82",
X"3d0d0480",
X"3d0d028b",
X"05339080",
X"a40c9080",
X"a8087081",
X"06515170",
X"f5389080",
X"a4087081",
X"ff0683c0",
X"800c5182",
X"3d0d0480",
X"3d0d81ff",
X"51d13f83",
X"c0800881",
X"ff0683c0",
X"800c823d",
X"0d04803d",
X"0d73902b",
X"73079080",
X"b40c823d",
X"0d0404fb",
X"3d0d7802",
X"84059f05",
X"3370982b",
X"55575572",
X"80259b38",
X"7580ff06",
X"56805280",
X"f751e03f",
X"83c08008",
X"81ff0654",
X"73812680",
X"ff388051",
X"fee73fff",
X"a23f8151",
X"fedf3fff",
X"9a3f7551",
X"feed3f74",
X"982a51fe",
X"e63f7490",
X"2a7081ff",
X"065253fe",
X"da3f7488",
X"2a7081ff",
X"065253fe",
X"ce3f7481",
X"ff0651fe",
X"c63f8155",
X"7580c02e",
X"09810686",
X"38819555",
X"8d397580",
X"c82e0981",
X"06843881",
X"87557451",
X"fea53f8a",
X"55fec83f",
X"83c08008",
X"81ff0670",
X"982b5454",
X"7280258c",
X"38ff1570",
X"81ff0656",
X"5374e238",
X"7383c080",
X"0c873d0d",
X"04fa3d0d",
X"fdc53f80",
X"51fdda3f",
X"8a54fe93",
X"3fff1470",
X"81ff0655",
X"5373f338",
X"73745355",
X"80c051fe",
X"a63f83c0",
X"800881ff",
X"06547381",
X"2e098106",
X"829f3883",
X"aa5280c8",
X"51fe8c3f",
X"83c08008",
X"81ff0653",
X"72812e09",
X"810681a8",
X"38745487",
X"3d741154",
X"56fdc83f",
X"83c08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e53802",
X"9a053353",
X"72812e09",
X"810681d9",
X"38029b05",
X"335380ce",
X"90547281",
X"aa2e8d38",
X"81c73980",
X"e4518b9a",
X"3fff1454",
X"73802e81",
X"b838820a",
X"5281e951",
X"fda53f83",
X"c0800881",
X"ff065372",
X"de387252",
X"80fa51fd",
X"923f83c0",
X"800881ff",
X"06537281",
X"90387254",
X"731653fc",
X"d63f83c0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e8",
X"38873d33",
X"70862a70",
X"81065154",
X"548c5572",
X"80e33884",
X"5580de39",
X"745281e9",
X"51fccc3f",
X"83c08008",
X"81ff0653",
X"825581e9",
X"56817327",
X"86387355",
X"80c15680",
X"ce90548a",
X"3980e451",
X"8a8c3fff",
X"14547380",
X"2ea93880",
X"527551fc",
X"9a3f83c0",
X"800881ff",
X"065372e1",
X"38848052",
X"80d051fc",
X"863f83c0",
X"800881ff",
X"06537280",
X"2e833880",
X"557483c3",
X"bc348051",
X"fb873ffb",
X"c23f883d",
X"0d04fb3d",
X"0d775480",
X"0b83c3bc",
X"3370832a",
X"70810651",
X"55575572",
X"752e0981",
X"06853873",
X"892b5473",
X"5280d151",
X"fbbd3f83",
X"c0800881",
X"ff065372",
X"bd3882b8",
X"c054fb83",
X"3f83c080",
X"0881ff06",
X"537281ff",
X"2e098106",
X"8938ff14",
X"5473e738",
X"9f397281",
X"fe2e0981",
X"06963883",
X"c7c05283",
X"c3c051fa",
X"ed3ffad3",
X"3ffad03f",
X"83398155",
X"8051fa89",
X"3ffac43f",
X"7481ff06",
X"83c0800c",
X"873d0d04",
X"fb3d0d77",
X"83c3c056",
X"548151f9",
X"ec3f83c3",
X"bc337083",
X"2a708106",
X"51545672",
X"85387389",
X"2b547352",
X"80d851fa",
X"b63f83c0",
X"800881ff",
X"06537280",
X"e43881ff",
X"51f9d43f",
X"81fe51f9",
X"ce3f8480",
X"53747081",
X"05563351",
X"f9c13fff",
X"137083ff",
X"ff065153",
X"72eb3872",
X"51f9b03f",
X"7251f9ab",
X"3ff9d03f",
X"83c08008",
X"9f0653a7",
X"88547285",
X"2e8c3899",
X"3980e451",
X"87c43fff",
X"1454f9b3",
X"3f83c080",
X"0881ff2e",
X"843873e9",
X"388051f8",
X"e43ff99f",
X"3f800b83",
X"c0800c87",
X"3d0d0471",
X"83c7c40c",
X"8880800b",
X"83c7c00c",
X"8480800b",
X"83c7c80c",
X"04fd3d0d",
X"77701755",
X"7705ff1a",
X"535371ff",
X"2e943873",
X"70810555",
X"33517073",
X"70810555",
X"34ff1252",
X"e939853d",
X"0d04fb3d",
X"0d87a681",
X"0b83c7c4",
X"08565675",
X"3383a680",
X"1634a054",
X"83a08053",
X"83c7c408",
X"5283c7c0",
X"0851ffb1",
X"3fa05483",
X"a4805383",
X"c7c40852",
X"83c7c008",
X"51ff9e3f",
X"905483a8",
X"805383c7",
X"c4085283",
X"c7c00851",
X"ff8b3fa0",
X"53805283",
X"c7c80883",
X"a0800551",
X"86953fa0",
X"53805283",
X"c7c80883",
X"a4800551",
X"86853f90",
X"53805283",
X"c7c80883",
X"a8800551",
X"85f53fff",
X"763483a0",
X"80548053",
X"83c7c408",
X"5283c7c8",
X"0851fec5",
X"3f80d080",
X"5483b080",
X"5383c7c4",
X"085283c7",
X"c80851fe",
X"b03f87ba",
X"3fa25480",
X"5383c7c8",
X"088c8005",
X"5281f1d8",
X"51fe9a3f",
X"860b87a8",
X"8334800b",
X"87a88234",
X"800b87a0",
X"9a34af0b",
X"87a09634",
X"bf0b87a0",
X"9734800b",
X"87a09834",
X"9f0b87a0",
X"9934800b",
X"87a09b34",
X"e00b87a8",
X"8934a20b",
X"87a88034",
X"830b87a4",
X"8f34820b",
X"87a88134",
X"873d0d04",
X"fc3d0d83",
X"a0805480",
X"5383c7c8",
X"085283c7",
X"c40851fd",
X"b83f80d0",
X"805483b0",
X"805383c7",
X"c8085283",
X"c7c40851",
X"fda33fa0",
X"5483a080",
X"5383c7c8",
X"085283c7",
X"c40851fd",
X"903fa054",
X"83a48053",
X"83c7c808",
X"5283c7c4",
X"0851fcfd",
X"3f905483",
X"a8805383",
X"c7c80852",
X"83c7c408",
X"51fcea3f",
X"83c7c408",
X"5583a680",
X"153387a6",
X"8134863d",
X"0d04fa3d",
X"0d787052",
X"55c1e33f",
X"83ffff0b",
X"83c08008",
X"25a93874",
X"51c1e43f",
X"83c08008",
X"9e3883c0",
X"80085788",
X"3dfc0554",
X"84808053",
X"83c7c408",
X"527451ff",
X"bf963fff",
X"bedc3f88",
X"3d0d04fa",
X"3d0d7870",
X"5255c1a2",
X"3f83ffff",
X"0b83c080",
X"08259638",
X"8057883d",
X"fc055484",
X"80805383",
X"c7c40852",
X"7451c095",
X"3f883d0d",
X"04803d0d",
X"90809008",
X"810683c0",
X"800c823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087081",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fd0676",
X"1007720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870822c",
X"bf0683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe830676",
X"822b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087088",
X"2c870683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f1ff06",
X"76882b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"912cbf06",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fc87",
X"ffff0676",
X"912b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087099",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70ffbf0a",
X"0676992b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90808008",
X"70882c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"0870892c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708a",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8b2c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708c2cbf",
X"0683c080",
X"0c51823d",
X"0d04fe3d",
X"0d7481e6",
X"29872a90",
X"80a00c84",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70810554",
X"34ff1151",
X"f039843d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"8405540c",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"84808053",
X"80528880",
X"0a51ffb3",
X"3f818080",
X"53805282",
X"800a51c6",
X"3f843d0d",
X"04803d0d",
X"8151fcaa",
X"3f72802e",
X"90388051",
X"fdfe3fcd",
X"3f83c7cc",
X"3351fdf4",
X"3f8151fc",
X"bb3f8051",
X"fcb63f80",
X"51fc873f",
X"823d0d04",
X"fd3d0d75",
X"52805480",
X"ff722588",
X"38810bff",
X"80135354",
X"ffbf1251",
X"70992686",
X"38e01252",
X"b039ff9f",
X"12519971",
X"27a738d0",
X"12e01354",
X"51708926",
X"85387252",
X"9839728f",
X"26853872",
X"528f3971",
X"ba2e0981",
X"0685389a",
X"52833980",
X"5273802e",
X"85388180",
X"12527181",
X"ff0683c0",
X"800c853d",
X"0d04803d",
X"0d84d8c0",
X"51807170",
X"81055334",
X"7084e0c0",
X"2e098106",
X"f038823d",
X"0d04fe3d",
X"0d029705",
X"3351fef4",
X"3f83c080",
X"0881ff06",
X"83c7d008",
X"54528073",
X"249b3883",
X"c8940813",
X"7283c898",
X"08075353",
X"71733483",
X"c7d00881",
X"0583c7d0",
X"0c843d0d",
X"04fa3d0d",
X"82800a1b",
X"55805788",
X"3dfc0554",
X"79537452",
X"7851ffba",
X"ac3f883d",
X"0d04fe3d",
X"0d83c7e8",
X"08527451",
X"c1903f83",
X"c080088c",
X"38765375",
X"5283c7e8",
X"0851c63f",
X"843d0d04",
X"fe3d0d83",
X"c7e80853",
X"75527451",
X"ffbbce3f",
X"83c08008",
X"8d387753",
X"765283c7",
X"e80851ff",
X"a03f843d",
X"0d04fe3d",
X"0d83c7e8",
X"0851ffba",
X"c13f83c0",
X"80088180",
X"802e0981",
X"06883883",
X"c1808053",
X"9c3983c7",
X"e80851ff",
X"baa43f83",
X"c0800880",
X"d0802e09",
X"81069338",
X"83c1b080",
X"5383c080",
X"085283c7",
X"e80851fe",
X"d43f843d",
X"0d04803d",
X"0df9fc3f",
X"83c08008",
X"842981f1",
X"fc057008",
X"83c0800c",
X"51823d0d",
X"04ed3d0d",
X"80448043",
X"80428041",
X"80705a5b",
X"fdcc3f80",
X"0b83c7d0",
X"0c800b83",
X"c8980c81",
X"eec051e9",
X"c53f8180",
X"0b83c898",
X"0c81eec4",
X"51e9b73f",
X"80d00b83",
X"c7d00c78",
X"30707a07",
X"80257087",
X"2b83c898",
X"0c5155f8",
X"ed3f83c0",
X"80085281",
X"eecc51e9",
X"913f80f8",
X"0b83c7d0",
X"0c788132",
X"70307072",
X"07802570",
X"872b83c8",
X"980c5156",
X"569eed3f",
X"83c08008",
X"5281eedc",
X"51e8e73f",
X"81a00b83",
X"c7d00c78",
X"82327030",
X"70720780",
X"2570872b",
X"83c8980c",
X"515656fe",
X"c53f83c0",
X"80085281",
X"eeec51e8",
X"bd3f81c8",
X"0b83c7d0",
X"0c788332",
X"70307072",
X"07802570",
X"872b83c8",
X"980c5156",
X"83c7e808",
X"5256ffb5",
X"983f83c0",
X"80085281",
X"eef451e8",
X"8d3f8298",
X"0b83c7d0",
X"0c810b83",
X"c7d45b58",
X"83c7d008",
X"83197a32",
X"70307072",
X"07802570",
X"872b83c8",
X"980c5157",
X"8e3d7055",
X"ff1b5457",
X"57579caf",
X"3f797084",
X"055b0851",
X"ffb4ce3f",
X"745483c0",
X"80085377",
X"5281eefc",
X"51e7bf3f",
X"a81783c7",
X"d00c8118",
X"5877852e",
X"098106ff",
X"af3883b8",
X"0b83c7d0",
X"0c788832",
X"70307072",
X"07802570",
X"872b83c8",
X"980c5156",
X"56f7b93f",
X"81ef8c55",
X"83c08008",
X"802e8f38",
X"83c7e408",
X"51ffb3f9",
X"3f83c080",
X"08557452",
X"81ef9451",
X"e6ec3f84",
X"880b83c7",
X"d00c7889",
X"32703070",
X"72078025",
X"70872b83",
X"c8980c51",
X"5681efa0",
X"5256e6ca",
X"3f84b00b",
X"83c7d00c",
X"788a3270",
X"30707207",
X"80257087",
X"2b83c898",
X"0c515681",
X"efac5256",
X"e6a83f85",
X"800b83c7",
X"d00c788b",
X"32703070",
X"72078025",
X"70872b83",
X"c8980c51",
X"5681efc8",
X"5256e686",
X"3f868da0",
X"51f7ef3f",
X"8052913d",
X"7052559f",
X"c13f8352",
X"74519fba",
X"3f635574",
X"83e13861",
X"19597880",
X"25853874",
X"5991398c",
X"79258638",
X"8c5983c5",
X"39788b26",
X"83bf3878",
X"822b5581",
X"e9ac1508",
X"04f58f3f",
X"83c08008",
X"61575575",
X"812e0981",
X"06893883",
X"c0800810",
X"55903975",
X"ff2e0981",
X"06883883",
X"c0800881",
X"2c559075",
X"25853890",
X"55883974",
X"80248338",
X"81557451",
X"f4e93f82",
X"f4399aef",
X"3f83c080",
X"08610555",
X"74802585",
X"38805588",
X"39877525",
X"83388755",
X"74518ed2",
X"3f82d239",
X"f4d93f83",
X"c0800861",
X"05557480",
X"25853880",
X"55883986",
X"75258338",
X"86557451",
X"f4d23f82",
X"b0396087",
X"3862802e",
X"82a73883",
X"c39c0883",
X"c3980cad",
X"ec0b83c3",
X"a00c83c7",
X"e80851d5",
X"9d3ff9ca",
X"3f828a39",
X"60568076",
X"259838ad",
X"8b0b83c3",
X"a00c83c7",
X"c4157008",
X"5255d4fe",
X"3f740852",
X"92397580",
X"25923883",
X"c7c41508",
X"51ffb0fb",
X"3f8052fc",
X"1951b839",
X"62802e81",
X"d03883c7",
X"c4157008",
X"83c7d408",
X"720c83c7",
X"d40cfc1a",
X"70535155",
X"8d9f3f83",
X"c0800856",
X"80518d95",
X"3f83c080",
X"08527451",
X"89ae3f75",
X"52805189",
X"a73f8199",
X"39605580",
X"7525b838",
X"83c3a808",
X"83c3980c",
X"adec0b83",
X"c3a00c83",
X"c7e40851",
X"d4883f83",
X"c7e40851",
X"d1a93f83",
X"c0800881",
X"ff067052",
X"55f3b23f",
X"74802e80",
X"e0388155",
X"80e33974",
X"802580d5",
X"3883c7e4",
X"0851ffaf",
X"ea3f8051",
X"f3933f80",
X"c4396280",
X"2ebf3883",
X"c3a40883",
X"c3980cad",
X"ec0b83c3",
X"a00c83c7",
X"ec0851d3",
X"b53f7889",
X"2e098106",
X"8b3883c7",
X"ec0851f0",
X"f63f9639",
X"788a2e09",
X"81068e38",
X"83c7ec08",
X"51f0a33f",
X"84396287",
X"387a802e",
X"f8ae3880",
X"557483c0",
X"800c953d",
X"0d04fe3d",
X"0d83c884",
X"51818395",
X"3f83c7f4",
X"5181838d",
X"3ff2ee3f",
X"83c08008",
X"802e8638",
X"8051818a",
X"39f2f33f",
X"83c08008",
X"80fe38f3",
X"933f83c0",
X"8008802e",
X"b9388151",
X"f0d03f80",
X"51f2a93f",
X"ecc83f80",
X"0b83c7d0",
X"0cf7c63f",
X"83c08008",
X"53ff0b83",
X"c7d00cee",
X"bb3f7280",
X"cb3883c7",
X"cc3351f2",
X"833f7251",
X"f0a03f80",
X"c039f2bb",
X"3f83c080",
X"08802eb5",
X"388151f0",
X"8d3f8051",
X"f1e63fec",
X"853fad8b",
X"0b83c3a0",
X"0c83c7d4",
X"0851d1e6",
X"3fff0b83",
X"c7d00ced",
X"f73f83c7",
X"d4085280",
X"5186d13f",
X"8151f3ad",
X"3f843d0d",
X"04fb3d0d",
X"805283c8",
X"845180f2",
X"9c3f8152",
X"83c7f451",
X"80f2923f",
X"800b83c7",
X"cc349080",
X"80528684",
X"808051ff",
X"b1c53f83",
X"c0800881",
X"a03883c7",
X"f0085181",
X"88c83f8a",
X"993f81f4",
X"9c51ffb5",
X"fb3f83c0",
X"8008559c",
X"800a5480",
X"c0805381",
X"efd05283",
X"c0800851",
X"f4f63f83",
X"c7e80853",
X"81efe052",
X"7451ffb0",
X"c43f83c0",
X"80088438",
X"f5843f83",
X"c7ec0853",
X"81efec52",
X"7451ffb0",
X"ac3f83c0",
X"8008b638",
X"873dfc05",
X"54848080",
X"5386a880",
X"805283c7",
X"ec0851ff",
X"aeb73f83",
X"c0800893",
X"38758480",
X"802e0981",
X"06893881",
X"0b83c7cc",
X"34873980",
X"0b83c7cc",
X"3483c7cc",
X"3351eff0",
X"3f8151f1",
X"dc3f93ca",
X"3f8151f1",
X"d43f8151",
X"fcf43ffa",
X"3983c08c",
X"080283c0",
X"8c0cfb3d",
X"0d0281ef",
X"f80b83c3",
X"9c0c81ef",
X"fc0b83c3",
X"940c81f0",
X"800b83c3",
X"a80c81f0",
X"840b83c3",
X"a40c83c0",
X"8c08fc05",
X"0c800b83",
X"c7d40b83",
X"c08c08f8",
X"050c83c0",
X"8c08f405",
X"0cffaebf",
X"3f83c080",
X"088605fc",
X"0683c08c",
X"08f0050c",
X"0283c08c",
X"08f00508",
X"310d833d",
X"7083c08c",
X"08f80508",
X"70840583",
X"c08c08f8",
X"050c0c51",
X"ffab803f",
X"83c08c08",
X"f4050881",
X"0583c08c",
X"08f4050c",
X"83c08c08",
X"f4050888",
X"2e098106",
X"ffab3886",
X"94808051",
X"e8993fff",
X"0b83c7d0",
X"0c800b83",
X"c8980c84",
X"d8c00b83",
X"c8940c81",
X"51ecbf3f",
X"8151ece4",
X"3f8051ec",
X"df3f8151",
X"ed853f82",
X"51edad3f",
X"8051edd5",
X"3f8051ed",
X"ff3f80d1",
X"ae528051",
X"dcfd3ffc",
X"bc3f83c0",
X"8c08fc05",
X"080d800b",
X"83c0800c",
X"873d0d83",
X"c08c0c04",
X"803d0d81",
X"ff51800b",
X"83c8a812",
X"34ff1151",
X"70f43882",
X"3d0d04ff",
X"3d0d7370",
X"33535181",
X"11337134",
X"71811234",
X"833d0d04",
X"ff3d0d83",
X"cac408a8",
X"2e098106",
X"8b3883ca",
X"dc0883ca",
X"c40c8739",
X"a80b83ca",
X"c40c83ca",
X"c4088605",
X"7081ff06",
X"5252d385",
X"3f833d0d",
X"04fb3d0d",
X"77795656",
X"80707155",
X"55527175",
X"25ac3872",
X"16703370",
X"147081ff",
X"06555151",
X"51717427",
X"89388112",
X"7081ff06",
X"53517181",
X"147083ff",
X"ff065552",
X"54747324",
X"d6387183",
X"c0800c87",
X"3d0d04fb",
X"3d0d7756",
X"8939f9c6",
X"3f8351ed",
X"ad3fd48c",
X"3f83c080",
X"08802eee",
X"3883cac4",
X"08860570",
X"81ff0652",
X"53d2923f",
X"810b9088",
X"d434f99e",
X"3f8351ed",
X"853f9088",
X"d4337081",
X"ff065553",
X"73802eea",
X"3873862a",
X"70810651",
X"5372ffbe",
X"3873982b",
X"53807324",
X"80de38d2",
X"fc3f83c0",
X"80085583",
X"c0800880",
X"cf387416",
X"75822b54",
X"549088c0",
X"13337434",
X"81155574",
X"852e0981",
X"06e83875",
X"3383c8a8",
X"34811633",
X"83c8a934",
X"82163383",
X"c8aa3483",
X"163383c8",
X"ab348452",
X"83c8a851",
X"fe933f83",
X"c0800881",
X"ff068417",
X"33555372",
X"742e8738",
X"fdce3ffe",
X"d13980e4",
X"51ebf73f",
X"873d0d04",
X"f43d0d7e",
X"60595580",
X"5d807582",
X"2b7183ca",
X"c8120c83",
X"cae0175b",
X"5b577679",
X"3477772e",
X"83b73876",
X"527751ff",
X"a99b3f8e",
X"3dfc0554",
X"905383ca",
X"b0527751",
X"ffa8d63f",
X"7c567590",
X"2e098106",
X"83933883",
X"cab051fc",
X"de3f83ca",
X"b251fcd7",
X"3f83cab4",
X"51fcd03f",
X"7683cac0",
X"0c7751ff",
X"a69b3f81",
X"edd05283",
X"c0800851",
X"c8bb3f83",
X"c0800881",
X"2e098106",
X"80d43876",
X"83cad80c",
X"820b83ca",
X"b034ff96",
X"0b83cab1",
X"347751ff",
X"a8e83f83",
X"c0800855",
X"83c08008",
X"77258838",
X"83c08008",
X"8f055574",
X"842c7083",
X"ffff0670",
X"882a5851",
X"557583ca",
X"b2347483",
X"cab33476",
X"83cab434",
X"ff800b83",
X"cab53481",
X"903983ca",
X"b03383ca",
X"b1337188",
X"2b07565b",
X"7483ffff",
X"2e098106",
X"80e838fe",
X"800b83ca",
X"d80c810b",
X"83cac00c",
X"ff0b83ca",
X"b034ff0b",
X"83cab134",
X"7751ffa7",
X"f53f83c0",
X"800883ca",
X"e40c83c0",
X"80085583",
X"c0800880",
X"25883883",
X"c080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583cab2",
X"347483ca",
X"b3347683",
X"cab434ff",
X"800b83ca",
X"b534810b",
X"83cabf34",
X"a5397485",
X"962e0981",
X"0680fe38",
X"7583cad8",
X"0c7751ff",
X"a7a93f83",
X"cabf3383",
X"c0800807",
X"557483ca",
X"bf3483ca",
X"bf338106",
X"5574802e",
X"83388457",
X"83cab433",
X"83cab533",
X"71882b07",
X"565c7481",
X"802e0981",
X"06a13883",
X"cab23383",
X"cab33371",
X"882b0756",
X"5bad8075",
X"27873876",
X"8207579c",
X"39768107",
X"57963974",
X"82802e09",
X"81068738",
X"76830757",
X"87397481",
X"ff268a38",
X"7783cac8",
X"1b0c7679",
X"348e3d0d",
X"04803d0d",
X"72842983",
X"cac80570",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d727083",
X"c8a00c70",
X"842981f3",
X"d0057008",
X"83cadc0c",
X"5151823d",
X"0d04fe3d",
X"0d8151de",
X"3f800b83",
X"caac0c80",
X"0b83caa8",
X"0cff0b83",
X"c8a40ca8",
X"0b83cac4",
X"0cae51cc",
X"c03f800b",
X"83cac854",
X"52807370",
X"8405550c",
X"81125271",
X"842e0981",
X"06ef3884",
X"3d0d04fe",
X"3d0d7402",
X"84059605",
X"22535371",
X"802e9638",
X"72708105",
X"543351cc",
X"cb3fff12",
X"7083ffff",
X"065152e7",
X"39843d0d",
X"04fe3d0d",
X"02920522",
X"5382ac51",
X"e6ec3f80",
X"c351cca8",
X"3f819651",
X"e6e03f72",
X"5283c8a8",
X"51ffb43f",
X"725283c8",
X"a851f8cd",
X"3f83c080",
X"0881ff06",
X"51cc853f",
X"843d0d04",
X"ffb13d0d",
X"80d13df8",
X"0551f8f7",
X"3f83caac",
X"08810583",
X"caac0c80",
X"cf3d33cf",
X"117081ff",
X"06515656",
X"74832688",
X"e638758f",
X"06ff0556",
X"7583c8a4",
X"082e9b38",
X"75832696",
X"387583c8",
X"a40c7584",
X"2983cac8",
X"05700853",
X"557551f9",
X"fb3f8076",
X"2488c238",
X"75842983",
X"cac80555",
X"7408802e",
X"88b33883",
X"c8a40884",
X"2983cac8",
X"05700802",
X"880582b9",
X"0533525b",
X"557480d2",
X"2e84b038",
X"7480d224",
X"903874bf",
X"2e9c3874",
X"80d02e81",
X"d53887f2",
X"397480d3",
X"2e80d338",
X"7480d72e",
X"81c43887",
X"e1390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290556",
X"56cb813f",
X"80c151ca",
X"bb3ff698",
X"3f83cadf",
X"3383c8a8",
X"34815283",
X"c8a851cb",
X"d83f8151",
X"fde73f74",
X"8b3883ca",
X"dc0883ca",
X"c40c8739",
X"a80b83ca",
X"c40ccacc",
X"3f80c151",
X"ca863ff5",
X"e33f900b",
X"83cabf33",
X"81065656",
X"74802e83",
X"38985683",
X"cab43383",
X"cab53371",
X"882b0756",
X"59748180",
X"2e098106",
X"9c3883ca",
X"b23383ca",
X"b3337188",
X"2b075657",
X"ad807527",
X"8c387581",
X"80075685",
X"3975a007",
X"567583c8",
X"a834ff0b",
X"83c8a934",
X"e00b83c8",
X"aa34800b",
X"83c8ab34",
X"845283c8",
X"a851cacd",
X"3f845186",
X"9b390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290556",
X"59c9c13f",
X"7951ffa1",
X"d63f83c0",
X"8008802e",
X"8a3880ce",
X"51c8ed3f",
X"85f13980",
X"c151c8e4",
X"3fc9d53f",
X"c88e3f83",
X"cad80858",
X"8375259b",
X"3883cab4",
X"3383cab5",
X"3371882b",
X"07fc1771",
X"297a0583",
X"80055a51",
X"578d3974",
X"81802918",
X"ff800558",
X"81805780",
X"5676762e",
X"9238c8c0",
X"3f83c080",
X"0883c8a8",
X"17348116",
X"56eb39c8",
X"af3f83c0",
X"800881ff",
X"06775383",
X"c8a85256",
X"f4bf3f83",
X"c0800881",
X"ff065575",
X"752e0981",
X"06819538",
X"9451e2aa",
X"3fc8a93f",
X"80c151c7",
X"e33fc8d4",
X"3f775279",
X"51ff9fe9",
X"3f805e80",
X"d13dfdf4",
X"05547653",
X"83c8a852",
X"7951ff9d",
X"ef3f0282",
X"b9053355",
X"81597480",
X"d72e0981",
X"0680c538",
X"77527951",
X"ff9fba3f",
X"80d13dfd",
X"f0055476",
X"538f3d70",
X"537a5258",
X"ff9ef23f",
X"80567676",
X"2ea23875",
X"1883c8a8",
X"17337133",
X"70723270",
X"30708025",
X"70307f06",
X"811d5d5f",
X"51515152",
X"5b55db39",
X"82ac51e1",
X"a53f7880",
X"2e863880",
X"c3518439",
X"80ce51c6",
X"d73fc7c8",
X"3fc6813f",
X"83d83902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"59558070",
X"5d5980e4",
X"51e0ef3f",
X"c6ee3f80",
X"c151c6a8",
X"3f83cac0",
X"08792e82",
X"d63883ca",
X"e40880fc",
X"055580fd",
X"52745185",
X"c13f83c0",
X"80085b77",
X"8224b238",
X"ff187087",
X"2b83ffff",
X"800681f2",
X"9c0583c8",
X"a8595755",
X"81805575",
X"70810557",
X"33777081",
X"055934ff",
X"157081ff",
X"06515574",
X"ea388285",
X"397782e8",
X"2e81a338",
X"7782e92e",
X"09810681",
X"aa387858",
X"77873270",
X"30707207",
X"80257a8a",
X"32703070",
X"72078025",
X"73075354",
X"5a515755",
X"75802e97",
X"38787826",
X"9238a00b",
X"83c8a81a",
X"34811970",
X"81ff065a",
X"55eb3981",
X"187081ff",
X"0659558a",
X"7827ffbc",
X"388f5883",
X"c8a31833",
X"83c8a819",
X"34ff1870",
X"81ff0659",
X"55778426",
X"ea389058",
X"800b83c8",
X"a8193481",
X"187081ff",
X"0670982b",
X"52595574",
X"8025e938",
X"80c6557a",
X"858f2484",
X"3880c255",
X"7483c8a8",
X"3480f10b",
X"83c8ab34",
X"810b83c8",
X"ac347a83",
X"c8a9347a",
X"882c5574",
X"83c8aa34",
X"80cb3982",
X"f0782580",
X"c4387780",
X"fd29fd97",
X"d3055279",
X"51ff9c95",
X"3f80d13d",
X"fdec0554",
X"80fd5383",
X"c8a85279",
X"51ff9bcd",
X"3f7b8119",
X"59567580",
X"fc248338",
X"78587788",
X"2c557483",
X"c9a53477",
X"83c9a634",
X"7583c9a7",
X"34818059",
X"80cc3983",
X"cad80857",
X"8378259b",
X"3883cab4",
X"3383cab5",
X"3371882b",
X"07fc1a71",
X"29790583",
X"80055951",
X"598d3977",
X"81802917",
X"ff800557",
X"81805976",
X"527951ff",
X"9ba33f80",
X"d13dfdec",
X"05547853",
X"83c8a852",
X"7951ff9a",
X"dc3f7851",
X"f6bf3fc3",
X"eb3fc2a4",
X"3f8b3983",
X"caa80881",
X"0583caa8",
X"0c80d13d",
X"0d04f6e0",
X"3ffc39fc",
X"3d0d7678",
X"71842983",
X"cac80570",
X"08515353",
X"53709e38",
X"80ce7234",
X"80cf0b81",
X"133480ce",
X"0b821334",
X"80c50b83",
X"13347084",
X"133480e7",
X"3983cae0",
X"13335480",
X"d2723473",
X"822a7081",
X"06515180",
X"cf537084",
X"3880d753",
X"72811334",
X"a00b8213",
X"34738306",
X"5170812e",
X"9e387081",
X"24883870",
X"802e8f38",
X"9f397082",
X"2e923870",
X"832e9238",
X"933980d8",
X"558e3980",
X"d3558939",
X"80cd5584",
X"3980c455",
X"74831334",
X"80c40b84",
X"1334800b",
X"85133486",
X"3d0d0483",
X"c8a00883",
X"c0800c04",
X"803d0d83",
X"c8a00884",
X"2981f3f0",
X"05700883",
X"c0800c51",
X"823d0d04",
X"fc3d0d76",
X"78535481",
X"53805587",
X"39711073",
X"10545273",
X"72265172",
X"802ea738",
X"70802e86",
X"38718025",
X"e8387280",
X"2e983871",
X"74268938",
X"73723175",
X"74075654",
X"72812a72",
X"812a5353",
X"e5397351",
X"78833874",
X"517083c0",
X"800c863d",
X"0d04fe3d",
X"0d805375",
X"527451ff",
X"a33f843d",
X"0d04fe3d",
X"0d815375",
X"527451ff",
X"933f843d",
X"0d04fb3d",
X"0d777955",
X"55805674",
X"76258638",
X"74305581",
X"56738025",
X"88387330",
X"76813257",
X"54805373",
X"527451fe",
X"e73f83c0",
X"80085475",
X"802e8738",
X"83c08008",
X"30547383",
X"c0800c87",
X"3d0d04fa",
X"3d0d787a",
X"57558057",
X"74772586",
X"38743055",
X"8157759f",
X"2c548153",
X"75743274",
X"31527451",
X"feaa3f83",
X"c0800854",
X"76802e87",
X"3883c080",
X"08305473",
X"83c0800c",
X"883d0d04",
X"fc3d0d76",
X"5580750c",
X"800b8416",
X"0c800b88",
X"160c800b",
X"8c160c83",
X"c8845180",
X"e9833f83",
X"c7f45180",
X"e8fb3f87",
X"a6803370",
X"81ff0670",
X"71842a06",
X"515152d9",
X"a03f7181",
X"2a813272",
X"81327181",
X"06718106",
X"3184180c",
X"54547183",
X"2a813272",
X"822a8132",
X"70810672",
X"7131780c",
X"51535387",
X"a0903387",
X"a0913370",
X"81ff0670",
X"73068132",
X"81068819",
X"0c515353",
X"83c08008",
X"802e80c2",
X"3883c080",
X"08812a70",
X"810683c0",
X"80088106",
X"3184170c",
X"5283c080",
X"08832a83",
X"c0800882",
X"2a718106",
X"71810631",
X"770c5353",
X"83c08008",
X"842a8106",
X"88160c83",
X"c0800885",
X"2a81068c",
X"160c863d",
X"0d04fe3d",
X"0d747654",
X"527151fe",
X"ab3f7281",
X"2ea23881",
X"73268d38",
X"72822ea8",
X"3872832e",
X"9c38e639",
X"7108e238",
X"841208dd",
X"38881208",
X"d838a539",
X"88120881",
X"2e9e3891",
X"39881208",
X"812e9538",
X"71089138",
X"8412088c",
X"388c1208",
X"812e0981",
X"06ffb238",
X"843d0d04",
X"fb3d0d78",
X"0284059f",
X"05335556",
X"800b81eb",
X"c8565381",
X"732b7406",
X"5271802e",
X"83388152",
X"74708205",
X"56227073",
X"902b0790",
X"809c0c51",
X"81135372",
X"882e0981",
X"06d93880",
X"5383caec",
X"13335170",
X"81ff2eb2",
X"38701081",
X"e9e80570",
X"22555180",
X"73177033",
X"701081e9",
X"e8057022",
X"51515152",
X"5273712e",
X"91388112",
X"5271862e",
X"098106f1",
X"38739080",
X"9c0c8113",
X"5372862e",
X"098106ff",
X"b8388053",
X"72167033",
X"51517081",
X"ff2e9438",
X"701081e9",
X"e8057022",
X"70848080",
X"0790809c",
X"0c515181",
X"13537286",
X"2e098106",
X"d7388053",
X"72165170",
X"3383caec",
X"14348113",
X"5372862e",
X"098106ec",
X"38873d0d",
X"0404ff3d",
X"0d740284",
X"058f0533",
X"52527088",
X"38719080",
X"940c8e39",
X"70812e09",
X"81068638",
X"71908098",
X"0c833d0d",
X"04fb3d0d",
X"029f0533",
X"79982b70",
X"982c7c98",
X"2b70982c",
X"83cb8815",
X"70337098",
X"2b70982c",
X"51585c5a",
X"51555154",
X"5470732e",
X"09810694",
X"3883cae8",
X"14337098",
X"2b70982c",
X"51525670",
X"722eb138",
X"72753471",
X"83cae815",
X"3483cae9",
X"3383cb89",
X"3371982b",
X"71902b07",
X"83cae833",
X"70882b72",
X"0783cb88",
X"33710790",
X"80b80c52",
X"59535452",
X"873d0d04",
X"fe3d0d74",
X"81113371",
X"3371882b",
X"0783c080",
X"0c535184",
X"3d0d0483",
X"caf43383",
X"c0800c04",
X"f53d0d02",
X"bb053302",
X"8405bf05",
X"33028805",
X"80c30533",
X"028c0580",
X"c6052266",
X"5c5a5e5c",
X"567a557b",
X"548953a1",
X"527d5180",
X"dedc3f83",
X"c0800881",
X"ff0683c0",
X"800c8d3d",
X"0d0483c0",
X"8c080283",
X"c08c0cf5",
X"3d0d83c0",
X"8c088805",
X"0883c08c",
X"088f0533",
X"83c08c08",
X"92052202",
X"8c057390",
X"0583c08c",
X"08e8050c",
X"83c08c08",
X"f8050c83",
X"c08c08f0",
X"050c83c0",
X"8c08ec05",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08f005",
X"0883c08c",
X"08e0050c",
X"83c08c08",
X"fc050c83",
X"c08c08f0",
X"05088927",
X"8a38890b",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"05088605",
X"87fffc06",
X"83c08c08",
X"e0050c02",
X"83c08c08",
X"e0050831",
X"0d853d70",
X"5583c08c",
X"08ec0508",
X"5483c08c",
X"08f00508",
X"5383c08c",
X"08f40508",
X"5283c08c",
X"08e4050c",
X"80e8b53f",
X"83c08008",
X"81ff0683",
X"c08c08e4",
X"050883c0",
X"8c08ec05",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"e0050880",
X"2e8c3883",
X"c08c08f8",
X"05080d89",
X"c83983c0",
X"8c08f005",
X"08802e89",
X"a63883c0",
X"8c08ec05",
X"08810533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508842e",
X"a938840b",
X"83c08c08",
X"e0050825",
X"88c73883",
X"c08c08e0",
X"0508852e",
X"859b3883",
X"c08c08e0",
X"0508a12e",
X"87ad3888",
X"ac39800b",
X"83c08c08",
X"ec050885",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08fc050c",
X"83c08c08",
X"e0050883",
X"2e098106",
X"88833883",
X"c08c08e8",
X"05088105",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e0050881",
X"2687e638",
X"810b83c0",
X"8c08e005",
X"0880d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08fc",
X"050c83c0",
X"8c08ec05",
X"08820533",
X"83c08c08",
X"e0050887",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088b",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"e005088c",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088d",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"e005088e",
X"052383c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088a",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"70940508",
X"fcffff06",
X"7194050c",
X"83c08c08",
X"e0050c83",
X"c08c08ec",
X"05088605",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"f4050c83",
X"c08c08e0",
X"050883c0",
X"8c08fc05",
X"082e0981",
X"06b63883",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c83",
X"c08c08fc",
X"050883c0",
X"8c08e005",
X"088b0534",
X"83c08c08",
X"ec050887",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"812e8f38",
X"83c08c08",
X"e0050882",
X"2eb73884",
X"8c3983c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c820b",
X"83c08c08",
X"e005088a",
X"053483d9",
X"3983c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08fc0508",
X"83c08c08",
X"e005088a",
X"053483a1",
X"3983c08c",
X"08fc0508",
X"802e8395",
X"3883c08c",
X"08ec0508",
X"83053383",
X"0683c08c",
X"08e0050c",
X"83c08c08",
X"e0050883",
X"2e098106",
X"82f33883",
X"c08c08ec",
X"05088205",
X"3370982b",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c83c0",
X"8c08e005",
X"08802582",
X"cc3883c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c83c0",
X"8c08ec05",
X"08860533",
X"83c08c08",
X"e0050880",
X"d6053483",
X"c08c08e0",
X"05088405",
X"83c08c08",
X"ec050882",
X"05338f06",
X"83c08c08",
X"e4050c83",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0883c08c",
X"08e00508",
X"3483c08c",
X"08ec0508",
X"84053383",
X"c08c08e0",
X"05088105",
X"34800b83",
X"c08c08e0",
X"05088205",
X"3483c08c",
X"08e00508",
X"08ff83ff",
X"06828007",
X"83c08c08",
X"e005080c",
X"83c08c08",
X"e8050881",
X"05338105",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"050883c0",
X"8c08e805",
X"08810534",
X"81833983",
X"c08c08fc",
X"0508802e",
X"80f73883",
X"c08c08ec",
X"05088605",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e00508a2",
X"2e098106",
X"80d73883",
X"c08c08ec",
X"05088805",
X"3383c08c",
X"08ec0508",
X"87053371",
X"82802905",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c5283c0",
X"8c08e405",
X"0c83c08c",
X"08f4050c",
X"83c08c08",
X"e4050883",
X"c08c08e0",
X"05088805",
X"2383c08c",
X"08ec0508",
X"3383c08c",
X"08f00508",
X"71317083",
X"ffff0683",
X"c08c08f0",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08ec0508",
X"0583c08c",
X"08ec050c",
X"f6d03983",
X"c08c08f8",
X"05080d83",
X"c08c08f0",
X"050883c0",
X"8c08e005",
X"0c83c08c",
X"08f80508",
X"0d83c08c",
X"08e00508",
X"83c0800c",
X"8d3d0d83",
X"c08c0c04",
X"83c08c08",
X"0283c08c",
X"0ce73d0d",
X"83c08c08",
X"88050802",
X"840583c0",
X"8c08e805",
X"0c83c08c",
X"08d4050c",
X"800b83cb",
X"903483c0",
X"8c08d405",
X"08900583",
X"c08c08c4",
X"050c800b",
X"83c08c08",
X"c4050834",
X"800b83c0",
X"8c08c405",
X"08810534",
X"800b83c0",
X"8c08c805",
X"0c83c08c",
X"08c80508",
X"80d82983",
X"c08c08c4",
X"05080583",
X"c08c08ff",
X"b8050c80",
X"0b83c08c",
X"08ffb805",
X"0880d805",
X"0c83c08c",
X"08ffb805",
X"08840583",
X"c08c08ff",
X"b8050c83",
X"c08c08c8",
X"050883c0",
X"8c08ffb8",
X"05083488",
X"0b83c08c",
X"08ffb805",
X"08810534",
X"800b83c0",
X"8c08ffb8",
X"05088205",
X"3483c08c",
X"08ffb805",
X"0808ffa1",
X"ff06a080",
X"0783c08c",
X"08ffb805",
X"080c83c0",
X"8c08c805",
X"08810570",
X"81ff0683",
X"c08c08c8",
X"050c83c0",
X"8c08ffb8",
X"050c810b",
X"83c08c08",
X"c8050827",
X"fedb3883",
X"c08c08ec",
X"05705483",
X"c08c08cc",
X"050c9252",
X"83c08c08",
X"d4050851",
X"80dbdc3f",
X"83c08008",
X"81ff0670",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffbc0508",
X"91c63883",
X"c08c08f4",
X"0551f18c",
X"3f83c080",
X"0883ffff",
X"0683c08c",
X"08f60552",
X"83c08c08",
X"e0050cf0",
X"f33f83c0",
X"800883ff",
X"ff0683c0",
X"8c08fd05",
X"3383c08c",
X"08ffbc05",
X"0883c08c",
X"08c8050c",
X"83c08c08",
X"c0050c83",
X"c08c08dc",
X"050c83c0",
X"8c08c805",
X"0883c08c",
X"08c00508",
X"2780fe38",
X"83c08c08",
X"cc050854",
X"83c08c08",
X"c8050853",
X"895283c0",
X"8c08d405",
X"085180da",
X"e33f83c0",
X"800881ff",
X"0683c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffbc05",
X"0883eb38",
X"83c08c08",
X"ee0551ef",
X"f33f83c0",
X"800883ff",
X"ff065383",
X"c08c08c8",
X"05085283",
X"c08c08d4",
X"050851f0",
X"b53f83c0",
X"8c08c805",
X"08810570",
X"81ff0683",
X"c08c08c8",
X"050c83c0",
X"8c08ffb8",
X"050cfef2",
X"3983c08c",
X"08c40508",
X"81053383",
X"c08c08c0",
X"050c83c0",
X"8c08c005",
X"08839e38",
X"83c08c08",
X"c0050883",
X"c08c08ff",
X"b8050c83",
X"c08c08e0",
X"050888de",
X"2e098106",
X"8b38810b",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"dc050885",
X"8e2e0981",
X"0682c538",
X"817083c0",
X"8c08ffb8",
X"05080683",
X"c08c08ff",
X"b8050c83",
X"c08c08c8",
X"050c83c0",
X"8c08ffb8",
X"0508802e",
X"829e3883",
X"c08c08c8",
X"050883c0",
X"8c08c405",
X"08810534",
X"83c08c08",
X"c0050883",
X"c08c08c4",
X"05088705",
X"3483c08c",
X"08c00508",
X"83c08c08",
X"c405088b",
X"053483c0",
X"8c08c005",
X"0883c08c",
X"08c40508",
X"8c053483",
X"0b83c08c",
X"08c40508",
X"8d053483",
X"c08c08c0",
X"050883c0",
X"8c08c405",
X"088e0523",
X"830b83c0",
X"8c08c405",
X"088a0534",
X"83c08c08",
X"c4050894",
X"05088380",
X"800783c0",
X"8c08c405",
X"0894050c",
X"83caf433",
X"7083c08c",
X"08c80508",
X"0583c08c",
X"08ffb805",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffb805",
X"0883caf4",
X"3483c08c",
X"08ffbc05",
X"0883c08c",
X"08c40508",
X"94053483",
X"c08c08c8",
X"050883c0",
X"8c08c405",
X"0880d605",
X"3483c08c",
X"08c80508",
X"83c08c08",
X"c4050884",
X"05348e0b",
X"83c08c08",
X"c4050885",
X"053483c0",
X"8c08c005",
X"0883c08c",
X"08c40508",
X"86053483",
X"c08c08c4",
X"05088405",
X"08ff83ff",
X"06828007",
X"83c08c08",
X"c4050884",
X"050ca239",
X"81db0b83",
X"c08c08ff",
X"b8050c8c",
X"c33983c0",
X"8c08ffbc",
X"050883c0",
X"8c08ffb8",
X"050c8cb0",
X"3983c08c",
X"08f10533",
X"5283c08c",
X"08d40508",
X"5180d6e8",
X"3f800b83",
X"c08c08c4",
X"05088105",
X"3383c08c",
X"08ffb805",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"c8050883",
X"c08c08ff",
X"b8050827",
X"8acb3883",
X"c08c08c8",
X"050880d8",
X"297083c0",
X"8c08c405",
X"08057088",
X"05708305",
X"3383c08c",
X"08ffb805",
X"0c83c08c",
X"08cc050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"d8050c83",
X"c08c08ff",
X"b8050888",
X"893883c0",
X"8c08ffbc",
X"05088d05",
X"3383c08c",
X"08d0050c",
X"83c08c08",
X"d0050887",
X"ed3883c0",
X"8c08cc05",
X"08220284",
X"05718605",
X"87fffc06",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"e4050c83",
X"c08c08c0",
X"050c0283",
X"c08c08ff",
X"b8050831",
X"0d893d70",
X"5983c08c",
X"08c00508",
X"5883c08c",
X"08ffbc05",
X"08870533",
X"5783c08c",
X"08ffb805",
X"0ca25583",
X"c08c08d0",
X"05085486",
X"53818152",
X"83c08c08",
X"d4050851",
X"80c99b3f",
X"83c08008",
X"81ff0683",
X"c08c08d0",
X"050c83c0",
X"8c08d005",
X"0881c038",
X"83c08c08",
X"ffbc0508",
X"96055383",
X"c08c08c0",
X"05085283",
X"c08c08ff",
X"b8050851",
X"accf3f83",
X"c0800881",
X"ff0683c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"0508802e",
X"81853883",
X"c08c08ff",
X"bc050894",
X"0583c08c",
X"08ffbc05",
X"08960533",
X"70862a83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08c0",
X"050c83c0",
X"8c08ffb8",
X"0508832e",
X"09810680",
X"c63883c0",
X"8c08ffb8",
X"050883c0",
X"8c08cc05",
X"08820534",
X"83caf433",
X"70810583",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"b8050883",
X"caf43483",
X"c08c08ff",
X"bc050883",
X"c08c08c0",
X"05083483",
X"c08c08e4",
X"05080d83",
X"c08c08d0",
X"050881ff",
X"0683c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffbc05",
X"08fbe338",
X"83c08c08",
X"d8050883",
X"c08c08c4",
X"05080588",
X"05708205",
X"335183c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"0508832e",
X"09810680",
X"e33883c0",
X"8c08ffbc",
X"050883c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"05088105",
X"7081ff06",
X"5183c08c",
X"08ffb805",
X"0c810b83",
X"c08c08ff",
X"b8050827",
X"dd38800b",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"81057081",
X"ff065183",
X"c08c08ff",
X"b8050c97",
X"0b83c08c",
X"08ffb805",
X"0827dd38",
X"83c08c08",
X"e0050880",
X"f9327030",
X"70802551",
X"5183c08c",
X"08ffb805",
X"0c83c08c",
X"08dc0508",
X"912e0981",
X"0680f938",
X"83c08c08",
X"ffb80508",
X"802e80ec",
X"3883c08c",
X"08c80508",
X"80e23885",
X"0b83c08c",
X"08c40508",
X"a60534a0",
X"0b83c08c",
X"08c40508",
X"a7053485",
X"0b83c08c",
X"08c40508",
X"a8053480",
X"c00b83c0",
X"8c08c405",
X"08a90534",
X"860b83c0",
X"8c08c405",
X"08aa0534",
X"900b83c0",
X"8c08c405",
X"08ab0534",
X"860b83c0",
X"8c08c405",
X"08ac0534",
X"a00b83c0",
X"8c08c405",
X"08ad0534",
X"83c08c08",
X"e0050889",
X"d8327030",
X"70802551",
X"5183c08c",
X"08ffb805",
X"0c83c08c",
X"08dc0508",
X"83edec2e",
X"09810680",
X"f6388170",
X"83c08c08",
X"ffb80508",
X"0683c08c",
X"08ffb805",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffb805",
X"08802e80",
X"ce3883c0",
X"8c08c805",
X"0880c438",
X"840b83c0",
X"8c08c405",
X"08aa0534",
X"80c00b83",
X"c08c08c4",
X"0508ab05",
X"34840b83",
X"c08c08c4",
X"0508ac05",
X"34900b83",
X"c08c08c4",
X"0508ad05",
X"3483c08c",
X"08ffbc05",
X"0883c08c",
X"08c40508",
X"8c053483",
X"c08c08e0",
X"050880f9",
X"32703070",
X"80255151",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"dc050886",
X"2e098106",
X"80c33881",
X"7083c08c",
X"08ffb805",
X"080683c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb8",
X"0508802e",
X"9c3883c0",
X"8c08c805",
X"08933883",
X"c08c08ff",
X"bc050883",
X"c08c08c4",
X"05088d05",
X"3483c08c",
X"08e00508",
X"b4b43270",
X"30708025",
X"515183c0",
X"8c08ffb8",
X"050c83c0",
X"8c08dc05",
X"0890892e",
X"098106a2",
X"3883c08c",
X"08ffb805",
X"08802e96",
X"3883c08c",
X"08c80508",
X"8d38820b",
X"83c08c08",
X"c405088d",
X"053483c0",
X"8c08c805",
X"0880d829",
X"83c08c08",
X"c4050805",
X"70840570",
X"83053383",
X"c08c08ff",
X"b8050c83",
X"c08c08cc",
X"050c83c0",
X"8c08c005",
X"0c805880",
X"5783c08c",
X"08ffb805",
X"08568055",
X"80548a53",
X"a15283c0",
X"8c08d405",
X"085180c1",
X"cd3f83c0",
X"800881ff",
X"06703070",
X"9f2a5183",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"bc0508a0",
X"2e8c3883",
X"c08c08ff",
X"b80508f5",
X"dd3883c0",
X"8c08c005",
X"088b0533",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"802eb438",
X"83c08c08",
X"cc050883",
X"053383c0",
X"8c08ffb8",
X"050c8058",
X"805783c0",
X"8c08ffb8",
X"05085680",
X"5580548b",
X"53a15283",
X"c08c08d4",
X"05085180",
X"c0c83f83",
X"c08c08c8",
X"05088105",
X"7081ff06",
X"83c08c08",
X"c4050881",
X"05335283",
X"c08c08c8",
X"050c83c0",
X"8c08ffb8",
X"050cf5a4",
X"39800b83",
X"c08c08c8",
X"050c83c0",
X"8c08c805",
X"0880d829",
X"83c08c08",
X"d4050805",
X"709a0533",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb80508",
X"822e0981",
X"06a93883",
X"cb905681",
X"55805483",
X"c08c08ff",
X"b8050853",
X"83c08c08",
X"ffbc0508",
X"97053352",
X"83c08c08",
X"d4050851",
X"e0ae3f83",
X"c08c08c8",
X"05088105",
X"7081ff06",
X"83c08c08",
X"c8050c83",
X"c08c08ff",
X"b8050c81",
X"0b83c08c",
X"08c80508",
X"27fefb38",
X"810b83c0",
X"8c08c405",
X"0834800b",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"e805080d",
X"83c08c08",
X"ffb80508",
X"83c0800c",
X"9b3d0d83",
X"c08c0c04",
X"f43d0d90",
X"1f59800b",
X"811a3355",
X"5b7a7427",
X"81ad387a",
X"80d82919",
X"8a113355",
X"5573832e",
X"09810681",
X"88389415",
X"33578052",
X"7651dde6",
X"3f805380",
X"527651de",
X"843fb3bc",
X"3f83c080",
X"085c8058",
X"7781c429",
X"1c871133",
X"55557380",
X"2e80c038",
X"740881e9",
X"dc2e0981",
X"06b53880",
X"755b5675",
X"80d8291a",
X"9a113355",
X"5573832e",
X"09810692",
X"38a41570",
X"33555576",
X"74278738",
X"ff145473",
X"75348116",
X"7081ff06",
X"57548176",
X"27d13881",
X"187081ff",
X"0659548f",
X"7827ffa4",
X"3883caf4",
X"33ff0554",
X"7383caf4",
X"34811b70",
X"81ff0681",
X"1b335f5c",
X"547c7b26",
X"fed53880",
X"0b83c080",
X"0c8e3d0d",
X"0483c08c",
X"080283c0",
X"8c0ce63d",
X"0d83c08c",
X"08880508",
X"02840571",
X"90057033",
X"7083c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08cc050c",
X"83c08c08",
X"dc050c83",
X"c08c08e0",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"9ee43880",
X"0b83c08c",
X"08cc0508",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08d4",
X"050c83c0",
X"8c08d405",
X"0883c08c",
X"08ffa405",
X"08259eac",
X"3883c08c",
X"08d40508",
X"80d82983",
X"c08c08cc",
X"05080584",
X"05708605",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffa405",
X"08802e9d",
X"b838b0e2",
X"3f83c08c",
X"08ffbc05",
X"0880d405",
X"0883c080",
X"08269da1",
X"380283c0",
X"8c08ffbc",
X"05088105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08d8050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"fc052383",
X"c08c08ff",
X"a4050886",
X"0583fc06",
X"83c08c08",
X"ffa4050c",
X"0283c08c",
X"08ffa405",
X"08310d85",
X"3d705583",
X"c08c08fc",
X"055483c0",
X"8c08ffbc",
X"05085383",
X"c08c08e0",
X"05085283",
X"c08c08c0",
X"050cb8ba",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"9bea3883",
X"c08c08ff",
X"bc050887",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"80d53883",
X"c08c08ff",
X"bc050886",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508822e",
X"098106b3",
X"3883c08c",
X"08fc0522",
X"83c08c08",
X"ffa4050c",
X"870b83c0",
X"8c08ffa4",
X"05082797",
X"3883c08c",
X"08c00508",
X"82055283",
X"c08c08c0",
X"05083351",
X"d7ba3f83",
X"c08c08ff",
X"bc050886",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508832e",
X"0981069a",
X"d33883c0",
X"8c08ffbc",
X"05089205",
X"83c08c08",
X"ffbc0508",
X"89053383",
X"c08c08ff",
X"a4050c83",
X"c08c08c4",
X"050c83c0",
X"8c08ffa4",
X"0508832e",
X"b63883c0",
X"8c08c405",
X"08820533",
X"83c08c08",
X"fc052283",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a8050883",
X"c08c08ff",
X"ac050826",
X"99ee3880",
X"0b83c08c",
X"08e4050c",
X"800b83c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa4",
X"0508832e",
X"09810688",
X"993883c0",
X"8c08c005",
X"083383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffb0",
X"05082e09",
X"810687d2",
X"3883c08c",
X"08c00508",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050894",
X"2e098106",
X"87b03883",
X"c08c08c0",
X"05088205",
X"33708106",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffb00508",
X"2e8a3888",
X"0b83c08c",
X"08e4050c",
X"83c08c08",
X"ffa80508",
X"812a7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"913883c0",
X"8c08e405",
X"08840783",
X"c08c08e4",
X"050c83c0",
X"8c08ffa8",
X"0508822a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9138",
X"83c08c08",
X"e4050882",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"ffa80508",
X"832a7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"913883c0",
X"8c08e405",
X"08810783",
X"c08c08e4",
X"050c83c0",
X"8c08c005",
X"08830533",
X"70982b83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050880",
X"25913883",
X"c08c08e4",
X"05089007",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"a8050881",
X"ff067085",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"08802e91",
X"3883c08c",
X"08e40508",
X"a00783c0",
X"8c08e405",
X"0c83c08c",
X"08ffa805",
X"08842a70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e923883",
X"c08c08e4",
X"050880c0",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"ffa80508",
X"862a7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"923883c0",
X"8c08e405",
X"08818007",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"a8050881",
X"0683c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e92",
X"3883c08c",
X"08e40508",
X"82800783",
X"c08c08e4",
X"050c83c0",
X"8c08ffa8",
X"0508812a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9238",
X"83c08c08",
X"e4050884",
X"800783c0",
X"8c08e405",
X"0c83c08c",
X"08c00508",
X"84053370",
X"982b83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa4",
X"05088025",
X"923883c0",
X"8c08e405",
X"08888007",
X"83c08c08",
X"e4050c83",
X"c08c08c0",
X"05088505",
X"3370982b",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa40508",
X"80259238",
X"83c08c08",
X"e4050890",
X"800783c0",
X"8c08e405",
X"0c83c08c",
X"08c00508",
X"82053370",
X"81ff0670",
X"852a7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"923883c0",
X"8c08e405",
X"08a08007",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"a8050884",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e93",
X"3883c08c",
X"08e40508",
X"80c08007",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"a8050886",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e93",
X"3883c08c",
X"08e40508",
X"81808007",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"ac050898",
X"2b83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802593",
X"3883c08c",
X"08e40508",
X"82808007",
X"83c08c08",
X"e4050c83",
X"c08c08c0",
X"05088705",
X"33818005",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"f8052383",
X"c08c08c0",
X"05088905",
X"33818005",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"fa052385",
X"eb39800b",
X"83c08c08",
X"e4050c81",
X"800b83c0",
X"8c08f805",
X"2381800b",
X"83c08c08",
X"fa052385",
X"cb3983c0",
X"8c08ffb0",
X"05081083",
X"c08c0805",
X"f80583c0",
X"8c08ffb0",
X"05088429",
X"83c08c08",
X"ffb00508",
X"100583c0",
X"8c08c405",
X"08057084",
X"05703383",
X"c08c08c0",
X"05080570",
X"3383c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb405",
X"0883c08c",
X"08ffb805",
X"082383c0",
X"8c08ffa8",
X"05088105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08902e09",
X"8106be38",
X"83c08c08",
X"ffa80508",
X"3383c08c",
X"08c00508",
X"05810570",
X"33708280",
X"2983c08c",
X"08ffb405",
X"08055151",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffb80508",
X"2383c08c",
X"08ffac05",
X"08860522",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa80508",
X"a23883c0",
X"8c08ffac",
X"05088805",
X"2283c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"0881ff2e",
X"80e53883",
X"c08c08ff",
X"b8050822",
X"7083c08c",
X"08ffa805",
X"08317082",
X"80297131",
X"83c08c08",
X"ffac0508",
X"88052270",
X"83c08c08",
X"ffa80508",
X"31707335",
X"5383c08c",
X"08ffa805",
X"0c83c08c",
X"08ffac05",
X"0c5183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffb8",
X"05082383",
X"c08c08ff",
X"b0050881",
X"057081ff",
X"0683c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa405",
X"0c810b83",
X"c08c08ff",
X"b0050827",
X"fce03883",
X"c08c08f8",
X"052283c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508bf26",
X"913883c0",
X"8c08e405",
X"08820783",
X"c08c08e4",
X"050c81c0",
X"0b83c08c",
X"08ffa405",
X"08279138",
X"83c08c08",
X"e4050881",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"fa052283",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a40508bf",
X"26913883",
X"c08c08e4",
X"05088807",
X"83c08c08",
X"e4050c81",
X"c00b83c0",
X"8c08ffa4",
X"05082791",
X"3883c08c",
X"08e40508",
X"840783c0",
X"8c08e405",
X"0c800b83",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"b0050810",
X"83c08c08",
X"c4050805",
X"70900570",
X"3383c08c",
X"08c00508",
X"05703372",
X"81053370",
X"72065153",
X"5183c08c",
X"08ffa805",
X"0c5183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"9b38900b",
X"83c08c08",
X"ffb00508",
X"2b83c08c",
X"08e40508",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"ffb00508",
X"81057081",
X"ff0683c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa4",
X"050c970b",
X"83c08c08",
X"ffb00508",
X"27fef438",
X"83c08c08",
X"ffbc0508",
X"90053383",
X"c08c08e4",
X"050883c0",
X"8c08ffa4",
X"050c83c0",
X"8c08c405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffbc05",
X"088c0508",
X"2e85e038",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffbc0508",
X"8c050c83",
X"c08c08ff",
X"bc050889",
X"053383c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa8",
X"0508802e",
X"859a3883",
X"c08c08e4",
X"0583c08c",
X"08ffa405",
X"0883c08c",
X"08ffa405",
X"088f0683",
X"c08c08e4",
X"050c83c0",
X"8c08ffb0",
X"050c83c0",
X"8c08d005",
X"0c83c08c",
X"08ffa805",
X"08822e09",
X"810681c2",
X"38800b83",
X"c08c08ff",
X"a4050886",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffa805",
X"082e8c38",
X"81c00b83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"b0050887",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e94",
X"3883c08c",
X"08ffa805",
X"08819032",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffb00508",
X"842a7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"943883c0",
X"8c08ffa8",
X"050880d0",
X"3283c08c",
X"08ffa805",
X"0c83c08c",
X"08ffb005",
X"0883c08c",
X"08ffa805",
X"083283c0",
X"8c08ffb0",
X"050c800b",
X"83c08c08",
X"f0050c80",
X"0b83c08c",
X"08f40523",
X"800b81eb",
X"d83383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffb8",
X"05082e82",
X"d33883c0",
X"8c08f005",
X"81ebd80b",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"c8050c83",
X"c08c08ff",
X"ac050833",
X"83c08c08",
X"ffac0508",
X"81053381",
X"722b8172",
X"2b077083",
X"c08c08ff",
X"b0050806",
X"5283c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffa805",
X"082e0981",
X"0681be38",
X"83c08c08",
X"ffb80508",
X"852680f6",
X"3883c08c",
X"08ffac05",
X"08820533",
X"7081ff06",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa40508",
X"802e80ca",
X"3883c08c",
X"08ffb805",
X"0883c08c",
X"08ffb805",
X"08810570",
X"81ff0683",
X"c08c08c8",
X"05087305",
X"5383c08c",
X"08ffb805",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb405",
X"0883c08c",
X"08ffa405",
X"083483c0",
X"8c08ffac",
X"05088305",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e9d",
X"38810b83",
X"c08c08ff",
X"a405082b",
X"83c08c08",
X"d0050808",
X"0783c08c",
X"08d00508",
X"0c83c08c",
X"08ffac05",
X"08840570",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa405",
X"08fdc838",
X"83c08c08",
X"f0055280",
X"51c2a93f",
X"83c08c08",
X"e4050852",
X"83c08c08",
X"c4050851",
X"c3e43f83",
X"c08c08fb",
X"05337081",
X"800a2981",
X"0a057098",
X"2c5583c0",
X"8c08ffa4",
X"050c83c0",
X"8c08f905",
X"33708180",
X"0a29810a",
X"0570982c",
X"5583c08c",
X"08ffa405",
X"0c83c08c",
X"08c40508",
X"5383c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa805",
X"0cc3ba3f",
X"83c08c08",
X"ffbc0508",
X"88053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e84e138",
X"83c08c08",
X"ffbc0508",
X"90053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050881",
X"2684c138",
X"807081ec",
X"980b81ec",
X"980b8105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffb405",
X"082e81ae",
X"3883c08c",
X"08ffac05",
X"08842983",
X"c08c08ff",
X"a8050805",
X"703383c0",
X"8c08c005",
X"08057033",
X"72810533",
X"70720651",
X"535183c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"aa38810b",
X"83c08c08",
X"ffac0508",
X"2b83c08c",
X"08ffb405",
X"08077083",
X"ffff0683",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"ac050881",
X"057081ff",
X"0681ec98",
X"71842971",
X"05708105",
X"33515383",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a40508fe",
X"d43883c0",
X"8c08ffbc",
X"05088a05",
X"2283c08c",
X"08c0050c",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"c005082e",
X"82ae3880",
X"0b83c08c",
X"08e8050c",
X"800b83c0",
X"8c08ec05",
X"23807083",
X"c08c08e8",
X"0583c08c",
X"08ffb805",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffb005",
X"0c81af39",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffac0508",
X"2c708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e80",
X"e73883c0",
X"8c08ffb0",
X"050883c0",
X"8c08ffb0",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ffb80508",
X"730583c0",
X"8c08ffbc",
X"05089005",
X"3383c08c",
X"08ffac05",
X"08842905",
X"535383c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050881ec",
X"9a053383",
X"c08c08ff",
X"a4050834",
X"83c08c08",
X"ffac0508",
X"81057081",
X"ff0683c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa4",
X"050c8f0b",
X"83c08c08",
X"ffac0508",
X"2783c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb005",
X"0885268c",
X"3883c08c",
X"08ffa405",
X"08fea938",
X"83c08c08",
X"e8055280",
X"51ffbcd8",
X"3f83c08c",
X"08ffb405",
X"0883c08c",
X"08ffbc05",
X"088a0523",
X"83c08c08",
X"ffbc0508",
X"80d20533",
X"83c08c08",
X"ffbc0508",
X"80d40508",
X"0583c08c",
X"08ffbc05",
X"0880d405",
X"0c83c08c",
X"08d80508",
X"0d83c08c",
X"08d40508",
X"81800a29",
X"81800a05",
X"70982c83",
X"c08c08cc",
X"05088105",
X"3383c08c",
X"08ffa805",
X"0c5183c0",
X"8c08d405",
X"0c83c08c",
X"08ffa805",
X"0883c08c",
X"08d40508",
X"24e1d638",
X"800b83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08dc05",
X"080d83c0",
X"8c08ffa8",
X"050883c0",
X"800c9c3d",
X"0d83c08c",
X"0c04f33d",
X"0d02bf05",
X"33028405",
X"80c30533",
X"83cb9033",
X"5a5b5979",
X"802e8d38",
X"78780657",
X"76802e8e",
X"38818a39",
X"78780657",
X"76802e81",
X"803883cb",
X"9033707a",
X"07585879",
X"88387809",
X"70790651",
X"577683cb",
X"90349298",
X"3f83c080",
X"085e805c",
X"8f5d7d1c",
X"87113358",
X"5876802e",
X"80c23877",
X"0881e9dc",
X"2e098106",
X"b738805b",
X"815a7d1c",
X"701c9a11",
X"33595959",
X"76822e09",
X"81069538",
X"83cb9056",
X"81558054",
X"76539718",
X"33527851",
X"ffbda93f",
X"ff1a80d8",
X"1c5c5a79",
X"8025cf38",
X"ff1d81c4",
X"1d5d5d7c",
X"8025ffa6",
X"388f3d0d",
X"04e93d0d",
X"696c0288",
X"0580ea05",
X"225c5a5b",
X"80707141",
X"5e58ff78",
X"797a7b7c",
X"7d464c4a",
X"45405d43",
X"62993d34",
X"62028405",
X"80dd0534",
X"77792280",
X"ffff0654",
X"45727923",
X"79782e88",
X"87387a70",
X"81055c33",
X"70842a71",
X"8c067082",
X"2a5a5656",
X"8306ff1b",
X"7083ffff",
X"065c5456",
X"80547574",
X"2e91387a",
X"7081055c",
X"33ff1b70",
X"83ffff06",
X"5c545481",
X"76279b38",
X"7381ff06",
X"7b708105",
X"5d335574",
X"82802905",
X"ff1b7083",
X"ffff065c",
X"54548276",
X"27aa3873",
X"83ffff06",
X"7b708105",
X"5d337090",
X"2b72077d",
X"7081055f",
X"3370982b",
X"7207fe1f",
X"7083ffff",
X"06405252",
X"52525454",
X"7e802e80",
X"c4387686",
X"f738748a",
X"2e098106",
X"9438811f",
X"7081ff06",
X"811e7081",
X"ff065f52",
X"405386dc",
X"39748c2e",
X"09810686",
X"d338ff1f",
X"7081ff06",
X"ff1e7081",
X"ff065f52",
X"40537b63",
X"2586bd38",
X"ff4386b8",
X"3976812e",
X"83bb3876",
X"81248938",
X"76802e8d",
X"3886a539",
X"76822e84",
X"a638869c",
X"39f81553",
X"72842684",
X"95387284",
X"2981ecd8",
X"05537208",
X"0464802e",
X"80cd3878",
X"22838080",
X"06537283",
X"80802e09",
X"8106bc38",
X"80567564",
X"27a43875",
X"1e7083ff",
X"ff067710",
X"1b901172",
X"832a5851",
X"57515373",
X"75347287",
X"0681712b",
X"51537281",
X"16348116",
X"7081ff06",
X"57539776",
X"27cc387f",
X"84074080",
X"0b993d43",
X"56611670",
X"3370982b",
X"70982c51",
X"51515380",
X"732480fb",
X"38607329",
X"1e7083ff",
X"ff067a22",
X"83808006",
X"52585372",
X"8380802e",
X"09810680",
X"de386088",
X"32703070",
X"72078025",
X"63903270",
X"30707207",
X"80257307",
X"53545851",
X"55537380",
X"2ebd3876",
X"87065372",
X"b6387584",
X"29761005",
X"79118411",
X"79832a57",
X"57515373",
X"75346081",
X"16346586",
X"14236688",
X"14237587",
X"387f8107",
X"408d3975",
X"812e0981",
X"0685387f",
X"82074081",
X"167081ff",
X"06575381",
X"7627fee5",
X"38636129",
X"1e7083ff",
X"ff065f53",
X"80704642",
X"ff028405",
X"80dd0534",
X"ff0b993d",
X"3483f539",
X"811c7081",
X"ff065d53",
X"80427381",
X"2e098106",
X"8e387781",
X"800a2981",
X"800a0558",
X"80d33973",
X"802e8938",
X"73822e09",
X"81068d38",
X"7c81800a",
X"2981800a",
X"055da439",
X"815f83b8",
X"39ff1c70",
X"81ff065d",
X"537b6325",
X"8338ff43",
X"7c802e92",
X"387c8180",
X"0a2981ff",
X"0a055d7c",
X"982c5d83",
X"93397780",
X"2e923877",
X"81800a29",
X"81ff0a05",
X"5877982c",
X"5882fd39",
X"7753839e",
X"39748926",
X"80f43874",
X"842981ec",
X"ec055372",
X"08047387",
X"2e82e138",
X"73852e82",
X"db387388",
X"2e82d538",
X"738c2e82",
X"cf387389",
X"2e098106",
X"86388145",
X"82c23973",
X"812e0981",
X"0682b938",
X"62802582",
X"b3387b98",
X"2b70982c",
X"514382a8",
X"397383ff",
X"ff064682",
X"9f397383",
X"ffff0647",
X"82963973",
X"81ff0641",
X"828e3973",
X"811a3482",
X"87397381",
X"ff064481",
X"ff397e53",
X"82a03974",
X"812e81e3",
X"38748124",
X"89387480",
X"2e8d3881",
X"e7397482",
X"2e81d838",
X"81de3974",
X"567b8338",
X"81567453",
X"73862e09",
X"81069738",
X"75810653",
X"72802e8e",
X"38782282",
X"ffff06fe",
X"80800753",
X"b6397b83",
X"38815373",
X"822e0981",
X"06973872",
X"81065372",
X"802e8e38",
X"782281ff",
X"ff068180",
X"80075393",
X"397b9638",
X"fc145372",
X"81268e38",
X"7822ff80",
X"80075372",
X"792380e5",
X"39805573",
X"812e0981",
X"06833873",
X"55775377",
X"802e8938",
X"74810653",
X"7280ca38",
X"72d01554",
X"55728126",
X"83388155",
X"77802eb9",
X"38748106",
X"5372802e",
X"b0387822",
X"83808006",
X"53728380",
X"802e0981",
X"069f3873",
X"b02e0981",
X"06873861",
X"993d3491",
X"3973b12e",
X"09810689",
X"38610284",
X"0580dd05",
X"34618105",
X"538c3961",
X"74318105",
X"53843961",
X"14537283",
X"ffff0642",
X"79f7fb38",
X"7d832a53",
X"72821a34",
X"78228380",
X"80065372",
X"8380802e",
X"09810688",
X"3881537f",
X"872e8338",
X"80537283",
X"c0800c99",
X"3d0d04fd",
X"3d0d7583",
X"11338212",
X"3371982b",
X"71902b07",
X"81143370",
X"882b7207",
X"75337107",
X"83c0800c",
X"52535456",
X"5452853d",
X"0d04f63d",
X"0d02b705",
X"33028405",
X"bb053302",
X"8805bf05",
X"335b5b5b",
X"80588057",
X"78882b7a",
X"07568055",
X"7a548153",
X"a3527c51",
X"92cc3f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f63d",
X"0d02b705",
X"33028405",
X"bb053302",
X"8805bf05",
X"335b5b5b",
X"80588057",
X"78882b7a",
X"07568055",
X"7a548353",
X"a3527c51",
X"92903f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f73d",
X"0d02b305",
X"33028405",
X"b6052260",
X"5a585680",
X"55805480",
X"5381a352",
X"7b5191e2",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8b3d0d04",
X"ee3d0d64",
X"90115c5c",
X"807b3480",
X"0b841c0c",
X"800b881c",
X"34810b89",
X"1c34880b",
X"8a1c3480",
X"0b8b1c34",
X"881b08c1",
X"06810788",
X"1c0c8f3d",
X"70545d88",
X"527b519c",
X"923f83c0",
X"800881ff",
X"06705b59",
X"7881a938",
X"903d335e",
X"81db5a7d",
X"892e0981",
X"06819938",
X"7c539252",
X"7b519beb",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"8182387c",
X"58885778",
X"56a95578",
X"54865381",
X"a0527b51",
X"90d03f83",
X"c0800881",
X"ff06705b",
X"597880e0",
X"3802ba05",
X"337b347c",
X"5478537d",
X"527b519b",
X"d33f83c0",
X"800881ff",
X"06705b59",
X"7880c138",
X"02bd0533",
X"527b519b",
X"eb3f83c0",
X"800881ff",
X"06705b59",
X"78aa3881",
X"7b335a5a",
X"79792699",
X"38805479",
X"5388527b",
X"51fdbb3f",
X"811a7081",
X"ff067c33",
X"525b59e4",
X"39810b88",
X"1c34805a",
X"7983c080",
X"0c943d0d",
X"04800b83",
X"c0800c04",
X"f93d0d79",
X"028405ab",
X"05338e3d",
X"70545858",
X"58ffb094",
X"3f8a3d8a",
X"0551ffb0",
X"8b3f7551",
X"fc8d3f83",
X"c0800884",
X"86812ebe",
X"3883c080",
X"08848681",
X"26993883",
X"c0800884",
X"82802e80",
X"e63883c0",
X"80088482",
X"812e9f38",
X"81b43983",
X"c0800880",
X"c082832e",
X"80f43883",
X"c0800880",
X"c086832e",
X"80e83881",
X"993983c0",
X"9c335580",
X"5674762e",
X"09810681",
X"8b387454",
X"76539152",
X"7751fbd6",
X"3f745476",
X"53905277",
X"51fbcb3f",
X"74547653",
X"84527751",
X"fbfc3f81",
X"0b83c09c",
X"3481b156",
X"80de3980",
X"54765391",
X"527751fb",
X"a93f8054",
X"76539052",
X"7751fb9e",
X"3f800b83",
X"c09c3476",
X"52871833",
X"5197963f",
X"b5398054",
X"76539452",
X"7751fb82",
X"3f805476",
X"53905277",
X"51faf73f",
X"7551ffae",
X"bf3f83c0",
X"8008892a",
X"81065376",
X"52871833",
X"5190cd3f",
X"800b83c0",
X"9c348056",
X"7583c080",
X"0c893d0d",
X"04f23d0d",
X"6090115a",
X"58800b88",
X"1a337159",
X"56567476",
X"2e82a538",
X"82ac3f84",
X"190883c0",
X"80082682",
X"95387833",
X"5a810b8e",
X"3d23903d",
X"f81155f4",
X"05539918",
X"5277518a",
X"e53f83c0",
X"800881ff",
X"06705755",
X"74772e09",
X"810681d9",
X"38863974",
X"5681d239",
X"81568257",
X"8e3d3377",
X"06557480",
X"2ebb3880",
X"0b8d3d34",
X"903df005",
X"54845375",
X"527751fa",
X"cd3f83c0",
X"800881ff",
X"0655749d",
X"387b5375",
X"527751fc",
X"e73f83c0",
X"800881ff",
X"06557481",
X"b12e818b",
X"3874ffb3",
X"38761081",
X"fc068117",
X"7081ff06",
X"58565787",
X"7627ffa8",
X"38815675",
X"7a2680eb",
X"38800b8d",
X"3d348c3d",
X"70555784",
X"53755277",
X"51f9f73f",
X"83c08008",
X"81ff0655",
X"7480c138",
X"7651ffac",
X"bb3f83c0",
X"80088287",
X"06557482",
X"812e0981",
X"06aa3802",
X"ae053381",
X"07557402",
X"8405ae05",
X"347b5375",
X"527751fb",
X"eb3f83c0",
X"800881ff",
X"06557481",
X"b12e9038",
X"74feb838",
X"81167081",
X"ff065755",
X"ff913980",
X"567581ff",
X"0656973f",
X"83c08008",
X"8fd00584",
X"1a0c7557",
X"7683c080",
X"0c903d0d",
X"04049080",
X"a00883c0",
X"800c04ff",
X"3d0d7387",
X"e82951ff",
X"80a03f83",
X"3d0d0404",
X"83cb940b",
X"83c0800c",
X"04fd3d0d",
X"75775454",
X"800b83ca",
X"f434728a",
X"38909080",
X"0b84150c",
X"90397281",
X"2e098106",
X"88389098",
X"800b8415",
X"0c841408",
X"83cb8c0c",
X"800b8815",
X"0c800b8c",
X"150c83cb",
X"8c085382",
X"0b878014",
X"348151ff",
X"9e3f83cb",
X"8c085380",
X"0b881434",
X"83cb8c08",
X"53810b87",
X"80143483",
X"cb8c0853",
X"800b8c14",
X"3483cb8c",
X"0853800b",
X"a4143491",
X"7434800b",
X"83c0a034",
X"800b83c0",
X"a434800b",
X"83c0a834",
X"80547381",
X"c42983cb",
X"98055380",
X"0b831434",
X"81147081",
X"ff065553",
X"8f7427e6",
X"38853d0d",
X"04fe3d0d",
X"74768211",
X"3370bf06",
X"81712bff",
X"05565151",
X"52539071",
X"278338ff",
X"52765171",
X"712383cb",
X"8c085187",
X"13339012",
X"34800b83",
X"c0a43480",
X"0b83c0a8",
X"34881333",
X"8a143352",
X"5271802e",
X"aa387081",
X"ff065184",
X"52708338",
X"70527183",
X"c0a4348a",
X"13337030",
X"70802584",
X"2b708807",
X"51515253",
X"7083c0a8",
X"34903970",
X"81ff0651",
X"70833898",
X"527183c0",
X"a834800b",
X"83c0800c",
X"843d0d04",
X"f13d0d61",
X"6568028c",
X"0580cb05",
X"33029005",
X"80ce0522",
X"02940580",
X"d6052242",
X"40415a40",
X"40fd8b3f",
X"83c08008",
X"a788055b",
X"8070715b",
X"5b528394",
X"3983cb8c",
X"08517d94",
X"123483c0",
X"a4338107",
X"55807054",
X"567f8626",
X"80ea387f",
X"842981ed",
X"a00583cb",
X"8c085351",
X"70080480",
X"0b841334",
X"a1397733",
X"70307080",
X"25837131",
X"51515253",
X"70841334",
X"8d39810b",
X"841334b8",
X"39830b84",
X"13348170",
X"5456ad39",
X"810b8413",
X"34a23977",
X"33703070",
X"80258371",
X"31515152",
X"53708413",
X"34807833",
X"52527083",
X"38815271",
X"78348153",
X"74880755",
X"83c0a833",
X"83cb8c08",
X"5257810b",
X"81d01234",
X"83cb8c08",
X"51810b81",
X"9012347e",
X"802eae38",
X"72802ea9",
X"387eff1e",
X"52547083",
X"ffff0653",
X"7283ffff",
X"2e973873",
X"70810555",
X"3383cb8c",
X"08535170",
X"81c01334",
X"ff1351de",
X"3983cb8c",
X"08a81133",
X"53517688",
X"123483cb",
X"8c085174",
X"713481ff",
X"52913983",
X"cb8c08a0",
X"11337081",
X"06515253",
X"708f38fa",
X"fd3f7a83",
X"c0800826",
X"e6388188",
X"39810ba0",
X"143483cb",
X"8c08a811",
X"3380ff06",
X"70780752",
X"53517080",
X"2e80ed38",
X"71862a70",
X"81065151",
X"70802e91",
X"38807833",
X"52537083",
X"38815372",
X"783480e0",
X"3971842a",
X"70810651",
X"5170802e",
X"9b388119",
X"7083ffff",
X"067d3070",
X"9f2a5152",
X"5a51787c",
X"2e098106",
X"af38a439",
X"71832a70",
X"81065151",
X"70802e93",
X"38811a70",
X"81ff065b",
X"5179832e",
X"09810690",
X"388a3971",
X"a3065170",
X"802e8538",
X"71519239",
X"f9e43f7a",
X"83c08008",
X"26fce238",
X"7181bf06",
X"517083c0",
X"800c913d",
X"0d04f63d",
X"0d02b305",
X"33028405",
X"b7053302",
X"8805ba05",
X"22595959",
X"800b8c3d",
X"348c3dfc",
X"05568055",
X"80547653",
X"77527851",
X"fbf23f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f33d",
X"0d7f6264",
X"028c0580",
X"c2052272",
X"22811533",
X"425f415e",
X"59598078",
X"237d5378",
X"33528151",
X"ffa03f83",
X"c0800881",
X"ff065675",
X"802e8638",
X"755481ad",
X"3983cb8c",
X"08a81133",
X"821b3370",
X"862a7081",
X"0673982b",
X"5351575c",
X"56577980",
X"25833881",
X"5673762e",
X"873881f0",
X"54818239",
X"818c1733",
X"7081ff06",
X"79227d71",
X"31902b70",
X"902c7009",
X"709f2c72",
X"06705252",
X"53515357",
X"57547574",
X"24833875",
X"55748480",
X"8029fc80",
X"80057090",
X"2c515574",
X"ff2e9438",
X"83cb8c08",
X"81801133",
X"5154737c",
X"7081055e",
X"34db3977",
X"22760554",
X"73782379",
X"09709f2a",
X"70810682",
X"1c3381bf",
X"0671862b",
X"07515151",
X"5473821a",
X"347c7626",
X"8a387722",
X"547a7426",
X"febb3880",
X"547383c0",
X"800c8f3d",
X"0d04f93d",
X"0d7a5780",
X"0b893d23",
X"893dfc05",
X"53765279",
X"51f8da3f",
X"83c08008",
X"81ff0670",
X"57557496",
X"387c547b",
X"53883d22",
X"527651fd",
X"e53f83c0",
X"800881ff",
X"06567583",
X"c0800c89",
X"3d0d04f0",
X"3d0d6266",
X"02880580",
X"ce052241",
X"5d5e8002",
X"840580d2",
X"05227f81",
X"0533ff11",
X"5a5d5a5d",
X"81da5876",
X"bf2680e9",
X"3878802e",
X"80e1387a",
X"58787b27",
X"83387858",
X"821e3370",
X"872a585a",
X"76923d34",
X"923dfc05",
X"5677557b",
X"547e537d",
X"33528251",
X"f8de3f83",
X"c0800881",
X"ff065d80",
X"0b923d33",
X"585a7680",
X"2e833881",
X"5a821e33",
X"80ff067a",
X"872b0757",
X"76821f34",
X"7c913878",
X"78317083",
X"ffff0679",
X"1e5e5a57",
X"ff9b397c",
X"587783c0",
X"800c923d",
X"0d04f83d",
X"0d7b0284",
X"05b20522",
X"5858800b",
X"8a3d238a",
X"3dfc0553",
X"77527a51",
X"f6f73f83",
X"c0800881",
X"ff067057",
X"55749638",
X"7d547653",
X"893d2252",
X"7751feaf",
X"3f83c080",
X"0881ff06",
X"567583c0",
X"800c8a3d",
X"0d04ec3d",
X"0d666e02",
X"880580df",
X"0533028c",
X"0580e305",
X"33029005",
X"80e70533",
X"02940580",
X"eb053302",
X"980580ee",
X"05224143",
X"415f5c40",
X"570280f2",
X"0522963d",
X"23963df0",
X"05538417",
X"70537752",
X"59f6863f",
X"83c08008",
X"81ff0658",
X"7781e538",
X"777a8180",
X"06584080",
X"77258338",
X"81407994",
X"3d347b02",
X"840580c9",
X"05347c02",
X"840580ca",
X"05347d02",
X"840580cb",
X"05347a95",
X"3d347a88",
X"2a577602",
X"840580cd",
X"0534953d",
X"22577602",
X"840580ce",
X"05347688",
X"2a577602",
X"840580cf",
X"05347792",
X"3d34963d",
X"ec115757",
X"8855f417",
X"54923d22",
X"53775277",
X"51f6953f",
X"83c08008",
X"81ff0658",
X"7780ed38",
X"7e802e80",
X"cb38923d",
X"22790858",
X"587f802e",
X"9c387681",
X"80800779",
X"0c7e5496",
X"3dfc0553",
X"7783ffff",
X"06527851",
X"f9fc3f99",
X"39768280",
X"8007790c",
X"7e54953d",
X"22537783",
X"ffff0652",
X"7851fc8f",
X"3f83c080",
X"0881ff06",
X"58779d38",
X"923d2253",
X"80527f30",
X"70802584",
X"71315351",
X"57f9873f",
X"83c08008",
X"81ff0658",
X"7783c080",
X"0c963d0d",
X"04f63d0d",
X"7c028405",
X"b705335b",
X"5b805880",
X"57805680",
X"55795485",
X"5380527a",
X"51fda33f",
X"83c08008",
X"81ff0659",
X"78853879",
X"871c3478",
X"83c0800c",
X"8c3d0d04",
X"f93d0d02",
X"a7053302",
X"8405ab05",
X"33028805",
X"af053358",
X"5957800b",
X"83cb9b33",
X"54547274",
X"2e9f3881",
X"147081ff",
X"06555373",
X"8f2681b6",
X"387381c4",
X"2983cb98",
X"05831133",
X"515372e3",
X"387381c4",
X"2983cb94",
X"0555800b",
X"87163476",
X"88163475",
X"8a163477",
X"89163480",
X"750c83cb",
X"8c088c16",
X"0c800b84",
X"1634880b",
X"85163480",
X"0b861634",
X"841508ff",
X"a1ff06a0",
X"80078416",
X"0c811470",
X"81ff0653",
X"537451fe",
X"bc3f83c0",
X"800881ff",
X"06705553",
X"7280cd38",
X"8a397308",
X"750c7254",
X"80c23972",
X"81f49055",
X"5681f490",
X"08802eb2",
X"38758429",
X"14700876",
X"53700851",
X"5454722d",
X"83c08008",
X"81ff0653",
X"72802ece",
X"38811670",
X"81ff0681",
X"f4907184",
X"29115356",
X"57537208",
X"d0388054",
X"7383c080",
X"0c893d0d",
X"04f93d0d",
X"7957800b",
X"84180883",
X"cb8c0c58",
X"f0883f88",
X"170883c0",
X"80082783",
X"ed38effa",
X"3f83c080",
X"08810588",
X"180c83cb",
X"8c08b811",
X"337081ff",
X"06515154",
X"73812ea4",
X"38738124",
X"88387378",
X"2e8a38b8",
X"3973822e",
X"9538b139",
X"763381f0",
X"06547390",
X"2ea63891",
X"7734a139",
X"73587633",
X"81f00654",
X"73902e09",
X"81069138",
X"efa83f83",
X"c0800881",
X"c8058c18",
X"0ca07734",
X"80567581",
X"c42983cb",
X"9b113355",
X"5573802e",
X"aa3883cb",
X"94157008",
X"56547480",
X"2e9d3888",
X"1508802e",
X"96388c14",
X"0883cb8c",
X"082e0981",
X"06893873",
X"51881508",
X"54732d81",
X"167081ff",
X"0657548f",
X"7627ffba",
X"38763354",
X"73b02e81",
X"993873b0",
X"248f3873",
X"912eab38",
X"73a02e80",
X"f53882a6",
X"397380d0",
X"2e81e438",
X"7380d024",
X"8b387380",
X"c02e8199",
X"38828f39",
X"7381802e",
X"81fb3882",
X"85398056",
X"7581c429",
X"83cb9811",
X"83113356",
X"59557380",
X"2ea83883",
X"cb941570",
X"08565474",
X"802e9b38",
X"8c140883",
X"cb8c082e",
X"0981068e",
X"38735184",
X"15085473",
X"2d800b83",
X"19348116",
X"7081ff06",
X"57548f76",
X"27ffb938",
X"92773481",
X"b539edc2",
X"3f8c1708",
X"83c08008",
X"2781a738",
X"b0773481",
X"a13983cb",
X"8c085480",
X"0b8c1534",
X"83cb8c08",
X"54840b88",
X"153480c0",
X"7734ed96",
X"3f83c080",
X"08b2058c",
X"180c80fa",
X"39ed873f",
X"8c170883",
X"c0800827",
X"80ec3883",
X"cb8c0854",
X"810b8c15",
X"3483cb8c",
X"0854800b",
X"88153483",
X"cb8c0854",
X"880ba015",
X"34ecdb3f",
X"83c08008",
X"94058c18",
X"0c80d077",
X"34bc3983",
X"cb8c08a0",
X"11337083",
X"2a708106",
X"51515555",
X"73802ea6",
X"38880ba0",
X"1634ecae",
X"3f8c1708",
X"83c08008",
X"279438ff",
X"8077348e",
X"39775380",
X"528051fa",
X"8b3fff90",
X"773483cb",
X"8c08a011",
X"3370832a",
X"70810651",
X"51555573",
X"802e8638",
X"880ba016",
X"34893d0d",
X"04f43d0d",
X"02bb0533",
X"028405bf",
X"05335d5d",
X"800b83cb",
X"980b83cb",
X"940b8c11",
X"72718814",
X"755c5a5b",
X"5f5c595b",
X"58831533",
X"5372802e",
X"81883873",
X"33537c73",
X"2e098106",
X"80fc3881",
X"1433537b",
X"732e0981",
X"0680ef38",
X"750883cb",
X"8c082e09",
X"810680e2",
X"38805675",
X"81c42983",
X"cb9c1170",
X"33831e33",
X"5b575553",
X"74782e09",
X"81069738",
X"83cba013",
X"0879082e",
X"0981068a",
X"38811433",
X"527451fe",
X"f83f8116",
X"7081ff06",
X"57538f76",
X"27c53880",
X"77085454",
X"72742e91",
X"38765184",
X"13085372",
X"2d83c080",
X"0881ff06",
X"54800b83",
X"1b347353",
X"a9398118",
X"81c41681",
X"c41681c4",
X"1981c41f",
X"81c41e81",
X"c41d6081",
X"c405415d",
X"5e5f5956",
X"56588f78",
X"25feca38",
X"80537283",
X"c0800c8e",
X"3d0d04f8",
X"3d0d02ae",
X"05227d59",
X"57805681",
X"55805486",
X"53818052",
X"7a51f4ee",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8a3d0d04",
X"f73d0d02",
X"b2052202",
X"8405b705",
X"33605a5b",
X"57805682",
X"55795486",
X"53818052",
X"7b51f4be",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8b3d0d04",
X"f83d0d02",
X"af053359",
X"80588057",
X"80568055",
X"78548953",
X"80527a51",
X"f4943f83",
X"c0800881",
X"ff0683c0",
X"800c8a3d",
X"0d04ffb8",
X"3d0d80cb",
X"3d087053",
X"81f0cc52",
X"56feadba",
X"3f83c080",
X"0880f338",
X"7551fea7",
X"a53f83ff",
X"ff0b83c0",
X"80082580",
X"e1387551",
X"fea7a43f",
X"83c08008",
X"5583c080",
X"0880cf38",
X"82805383",
X"c0800852",
X"8a3d7052",
X"57fee8fb",
X"3f745275",
X"51fea6b5",
X"3f805980",
X"ca3dfdfc",
X"05548280",
X"53765275",
X"51fea4bc",
X"3f811555",
X"7488802e",
X"098106e1",
X"38805275",
X"51fea68d",
X"3f800b83",
X"e3d80c75",
X"83e3d40c",
X"8739800b",
X"83e3d40c",
X"80ca3d0d",
X"04ff3d0d",
X"73700853",
X"51029305",
X"33723470",
X"08810571",
X"0c833d0d",
X"04ffb83d",
X"0d80cb3d",
X"70708405",
X"52085856",
X"83e3d408",
X"802e80fa",
X"388a3d70",
X"5a765577",
X"5481e6ed",
X"5380cb3d",
X"fdfc0552",
X"55fed2cb",
X"3f805280",
X"ca3dfdfc",
X"0551ffad",
X"3f83e3d8",
X"085283e3",
X"d40851fe",
X"a5933f80",
X"587451fe",
X"d0913f80",
X"ca3dfdf8",
X"055483c0",
X"80085374",
X"5283e3d4",
X"0851fea3",
X"8f3f83e3",
X"d8081883",
X"e3d80c80",
X"ca3dfdf8",
X"05548153",
X"81f0d852",
X"83e3d408",
X"51fea2f0",
X"3f83e3d8",
X"081883e3",
X"d80c80ca",
X"3d0d0400",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002bdd",
X"00002c1e",
X"00002c40",
X"00002c62",
X"00002c88",
X"00002c88",
X"00002c88",
X"00002c88",
X"00002cf9",
X"00002d4e",
X"00002d4e",
X"00002d8e",
X"0000435c",
X"00004d7c",
X"00004e45",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3f00",
X"0c0c4000",
X"0a0a4100",
X"0b0b4100",
X"07074100",
X"0a0b4300",
X"080b4200",
X"04044500",
X"05054400",
X"0e0f2900",
X"06060004",
X"08080004",
X"09090004",
X"0a0f4300",
X"090f4200",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"00006001",
X"00006308",
X"00006114",
X"00006308",
X"00006151",
X"000061a2",
X"000061e1",
X"000061ea",
X"00006308",
X"00006308",
X"00006308",
X"00006308",
X"000061f3",
X"000061fb",
X"00006202",
X"00006408",
X"00006501",
X"00006615",
X"0000690b",
X"00006926",
X"00006912",
X"00006926",
X"0000692d",
X"00006938",
X"0000693f",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"43505520",
X"54757262",
X"6f3a2564",
X"78000000",
X"44726976",
X"65205475",
X"72626f3a",
X"25730000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"4c6f6164",
X"206d656d",
X"6f727900",
X"53617665",
X"206d656d",
X"6f727920",
X"28666f72",
X"20646562",
X"75676769",
X"6e672900",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"66726565",
X"7a65722e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"4d454d00",
X"5374616e",
X"64617264",
X"00000000",
X"46617374",
X"28362900",
X"46617374",
X"28352900",
X"46617374",
X"28342900",
X"46617374",
X"28332900",
X"46617374",
X"28322900",
X"46617374",
X"28312900",
X"46617374",
X"28302900",
X"2f757362",
X"2e6c6f67",
X"00000000",
X"0a000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"000076fc",
X"00007700",
X"00007708",
X"00007714",
X"00007720",
X"0000772c",
X"00007738",
X"0000773c",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00000028",
X"00000006",
X"00000005",
X"00000004",
X"00000003",
X"00000002",
X"00000001",
X"00000000",
X"00007808",
X"00007814",
X"0000781c",
X"00007824",
X"0000782c",
X"00007834",
X"0000783c",
X"00007844",
X"00007694",
X"000074dc",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"69383030",
X"00000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
