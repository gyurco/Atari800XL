
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81ca",
X"d0738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81d1",
X"e00c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757581c4",
X"ff2d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7581c393",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80dea704",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"775193c4",
X"3f83c080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3381d1e8",
X"0b81d1e8",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"52775192",
X"f33f83c0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583c0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"55b3aa3f",
X"83c08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"811451b2",
X"c23f83c0",
X"80083070",
X"83c08008",
X"07802583",
X"c0800c53",
X"863d0d04",
X"fc3d0d76",
X"70525599",
X"e03f83c0",
X"80085481",
X"5383c080",
X"0880c738",
X"745199a3",
X"3f83c080",
X"080b0b81",
X"cffc5383",
X"c0800852",
X"53ff8f3f",
X"83c08008",
X"a5380b0b",
X"81d08052",
X"7251fefe",
X"3f83c080",
X"0894380b",
X"0b81d084",
X"527251fe",
X"ed3f83c0",
X"8008802e",
X"83388154",
X"73537283",
X"c0800c86",
X"3d0d04fd",
X"3d0d7570",
X"525498f9",
X"3f815383",
X"c0800898",
X"38735198",
X"c23f83c0",
X"b0085283",
X"c0800851",
X"feb43f83",
X"c0800853",
X"7283c080",
X"0c853d0d",
X"04df3d0d",
X"a43d0870",
X"525e8ee7",
X"3f83c080",
X"0833953d",
X"56547396",
X"3881d384",
X"527451b1",
X"9c3f9a39",
X"7d527851",
X"91e83f84",
X"e3397d51",
X"8ecd3f83",
X"c0800852",
X"74518dfd",
X"3f804380",
X"42804180",
X"4083c0b8",
X"0852943d",
X"70525d94",
X"d03f83c0",
X"80085980",
X"0b83c080",
X"08555b83",
X"c080087b",
X"2e943881",
X"1b74525b",
X"97d23f83",
X"c0800854",
X"83c08008",
X"ee38805a",
X"ff5f7909",
X"709f2c7b",
X"065b547a",
X"7a248438",
X"ff1b5af6",
X"1a700970",
X"9f2c7206",
X"7bff125a",
X"5a525555",
X"80752595",
X"38765197",
X"973f83c0",
X"800876ff",
X"18585557",
X"738024ed",
X"38747f2e",
X"873880c3",
X"853f745f",
X"78ff1b70",
X"585d5880",
X"7a259538",
X"775196ec",
X"3f83c080",
X"0876ff18",
X"58555873",
X"8024ed38",
X"800b83c7",
X"cc0c800b",
X"83c8900c",
X"0b0b81d0",
X"88518bbe",
X"3f81800b",
X"83c8900c",
X"0b0b81d0",
X"90518bae",
X"3fa80b83",
X"c7cc0c76",
X"802e80e8",
X"3883c7cc",
X"08777932",
X"70307072",
X"07802570",
X"872b83c8",
X"900c5156",
X"78535656",
X"969f3f83",
X"c0800880",
X"2e8a380b",
X"0b81d098",
X"518af33f",
X"765195df",
X"3f83c080",
X"08520b0b",
X"81d1ac51",
X"8ae03f76",
X"5195e53f",
X"83c08008",
X"83c7cc08",
X"55577574",
X"258638a8",
X"1656f739",
X"7583c7cc",
X"0c86f076",
X"24ff9438",
X"87980b83",
X"c7cc0c77",
X"802eb738",
X"7751959b",
X"3f83c080",
X"08785255",
X"95bb3f0b",
X"0b81d0a0",
X"5483c080",
X"088f3887",
X"39807634",
X"81d8390b",
X"0b81d09c",
X"54745373",
X"520b0b81",
X"cfec5189",
X"f93f8054",
X"0b0b81cf",
X"f45189ee",
X"3f811454",
X"73a82e09",
X"8106ed38",
X"868da051",
X"befb3f80",
X"52903d70",
X"525780d2",
X"943f8352",
X"765180d2",
X"8c3f6281",
X"91386180",
X"2e80fd38",
X"7b5473ff",
X"2e963878",
X"802e818c",
X"38785194",
X"b73f83c0",
X"8008ff15",
X"5559e739",
X"78802e80",
X"f7387851",
X"94b33f83",
X"c0800880",
X"2efbfd38",
X"785193fb",
X"3f83c080",
X"08520b0b",
X"81cff851",
X"abdc3f83",
X"c08008a3",
X"387c51ad",
X"943f83c0",
X"80085574",
X"ff165654",
X"807425ae",
X"38741d70",
X"33555673",
X"af2efec5",
X"38e93978",
X"5193ba3f",
X"83c08008",
X"527c51ac",
X"cc3f8f39",
X"7f882960",
X"10057a05",
X"61055afb",
X"fd396280",
X"2efbbe38",
X"80527651",
X"80d0ea3f",
X"a33d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"842a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"a80b9088",
X"b834b80b",
X"9088b834",
X"7083c080",
X"0c823d0d",
X"04803d0d",
X"9088b833",
X"7081ff06",
X"70852a81",
X"32708106",
X"51515151",
X"70802e8d",
X"38980b90",
X"88b834b8",
X"0b9088b8",
X"347083c0",
X"800c823d",
X"0d04930b",
X"9088bc34",
X"ff0b9088",
X"a83404ff",
X"3d0d028f",
X"05335280",
X"0b9088bc",
X"348a51bc",
X"c03fdf3f",
X"80f80b90",
X"88a03480",
X"0b908888",
X"34fa1252",
X"71908880",
X"34800b90",
X"88983471",
X"90889034",
X"9088b852",
X"807234b8",
X"7234833d",
X"0d04803d",
X"0d028b05",
X"33517090",
X"88b434fe",
X"bf3f83c0",
X"8008802e",
X"f638823d",
X"0d04803d",
X"0d853980",
X"c9ba3ffe",
X"d83f83c0",
X"8008802e",
X"f2389088",
X"b4337081",
X"ff0683c0",
X"800c5182",
X"3d0d0480",
X"3d0da30b",
X"9088bc34",
X"ff0b9088",
X"a8349088",
X"b851a871",
X"34b87134",
X"823d0d04",
X"803d0d90",
X"88bc3370",
X"81c00670",
X"30708025",
X"83c0800c",
X"51515182",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067083",
X"2a813270",
X"81065151",
X"51517080",
X"2ee838b0",
X"0b9088b8",
X"34b80b90",
X"88b83482",
X"3d0d0480",
X"3d0d9080",
X"ac088106",
X"83c0800c",
X"823d0d04",
X"fd3d0d75",
X"77545480",
X"73259438",
X"73708105",
X"55335281",
X"d0a45185",
X"a13fff13",
X"53e93985",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"81ade23f",
X"83c08008",
X"7a27ed38",
X"74802e80",
X"e0387452",
X"755181ad",
X"cc3f83c0",
X"80087553",
X"76525481",
X"adf23f83",
X"c080087a",
X"53755256",
X"81adb23f",
X"83c08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"c08008c2",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9c",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fbfd3f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd13f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbad3f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83c0900c",
X"7183c094",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383c090",
X"085283c0",
X"940851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"99e65351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fd3d",
X"0d757052",
X"54a3c63f",
X"83c08008",
X"14537274",
X"2e9238ff",
X"13703353",
X"5371af2e",
X"098106ee",
X"38811353",
X"7283c080",
X"0c853d0d",
X"04fd3d0d",
X"75777053",
X"5454c73f",
X"83c08008",
X"732ea138",
X"83c08008",
X"733152ff",
X"125271ff",
X"2e8f3872",
X"70810554",
X"33747081",
X"055634eb",
X"39ff1454",
X"80743485",
X"3d0d0480",
X"3d0d7251",
X"ff903f82",
X"3d0d0471",
X"83c0800c",
X"04803d0d",
X"72518071",
X"34810bbc",
X"120c800b",
X"80c0120c",
X"823d0d04",
X"800b83c2",
X"e408248a",
X"38a4b03f",
X"ff0b83c2",
X"e40c800b",
X"83c0800c",
X"04ff3d0d",
X"735283c0",
X"c008722e",
X"8d38d93f",
X"71519699",
X"3f7183c0",
X"c00c833d",
X"0d04f43d",
X"0d7e6062",
X"5c5a5581",
X"54bc1508",
X"81913874",
X"51cf3f79",
X"58807a25",
X"80f73883",
X"c3940870",
X"892a5783",
X"ff067884",
X"80723156",
X"56577378",
X"25833873",
X"557583c2",
X"e4082e84",
X"38ff893f",
X"83c2e408",
X"8025a638",
X"75892b51",
X"98dc3f83",
X"c394088f",
X"3dfc1155",
X"5c548152",
X"f81b5196",
X"c63f7614",
X"83c3940c",
X"7583c2e4",
X"0c745376",
X"527851a2",
X"e13f83c0",
X"800883c3",
X"94081683",
X"c3940c78",
X"7631761b",
X"5b595677",
X"8024ff8b",
X"38617a71",
X"0c547554",
X"75802e83",
X"38815473",
X"83c0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"9b3f7651",
X"feaf3f86",
X"3dfc0553",
X"78527751",
X"95e93f79",
X"75710c54",
X"83c08008",
X"5483c080",
X"08802e83",
X"38815473",
X"83c0800c",
X"863d0d04",
X"fe3d0d75",
X"83c2e408",
X"53538072",
X"24893871",
X"732e8438",
X"fdd63f74",
X"51fdea3f",
X"725197ae",
X"3f83c080",
X"085283c0",
X"8008802e",
X"83388152",
X"7183c080",
X"0c843d0d",
X"04803d0d",
X"7280c011",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d72bc11",
X"0883c080",
X"0c51823d",
X"0d0480c4",
X"0b83c080",
X"0c04fd3d",
X"0d757771",
X"54705355",
X"539f9e3f",
X"82c81308",
X"bc150c82",
X"c0130880",
X"c0150cfc",
X"eb3f7351",
X"93ab3f73",
X"83c0c00c",
X"83c08008",
X"5383c080",
X"08802e83",
X"38815372",
X"83c0800c",
X"853d0d04",
X"fd3d0d75",
X"775553fc",
X"bf3f7280",
X"2ea538bc",
X"13085273",
X"519ea83f",
X"83c08008",
X"8f387752",
X"7251ff9a",
X"3f83c080",
X"08538a39",
X"82cc1308",
X"53d83981",
X"537283c0",
X"800c853d",
X"0d04fe3d",
X"0dff0b83",
X"c2e40c74",
X"83c0c40c",
X"7583c2e0",
X"0c9f953f",
X"83c08008",
X"81ff0652",
X"81537199",
X"3883c2fc",
X"518e943f",
X"83c08008",
X"5283c080",
X"08802e83",
X"38725271",
X"537283c0",
X"800c843d",
X"0d04fa3d",
X"0d787a82",
X"c4120882",
X"c4120870",
X"72245956",
X"56575773",
X"732e0981",
X"06913880",
X"c0165280",
X"c017519c",
X"993f83c0",
X"80085574",
X"83c0800c",
X"883d0d04",
X"f63d0d7c",
X"5b807b71",
X"5c54577a",
X"772e8c38",
X"811a82cc",
X"1408545a",
X"72f63880",
X"5980d939",
X"7a548157",
X"80707b7b",
X"315a5755",
X"ff185374",
X"732580c1",
X"3882cc14",
X"08527351",
X"ff8c3f80",
X"0b83c080",
X"0825a138",
X"82cc1408",
X"82cc1108",
X"82cc160c",
X"7482cc12",
X"0c537580",
X"2e863872",
X"82cc170c",
X"72548057",
X"7382cc15",
X"08811757",
X"5556ffb8",
X"39811959",
X"800bff1b",
X"54547873",
X"25833881",
X"54768132",
X"70750651",
X"5372ff90",
X"388c3d0d",
X"04f73d0d",
X"7b7d5a5a",
X"82d05283",
X"c2e00851",
X"81a0ea3f",
X"83c08008",
X"57f9e13f",
X"795283c2",
X"e85195b7",
X"3f83c080",
X"08548053",
X"83c08008",
X"732e0981",
X"06828338",
X"83c0c408",
X"0b0b81cf",
X"f8537052",
X"569bd63f",
X"0b0b81cf",
X"f85280c0",
X"16519bc9",
X"3f75bc17",
X"0c7382c0",
X"170c810b",
X"82c4170c",
X"810b82c8",
X"170c7382",
X"cc170cff",
X"1782d017",
X"55578191",
X"3983c0d0",
X"3370822a",
X"70810651",
X"54557281",
X"80387481",
X"2a810658",
X"7780f638",
X"74842a81",
X"0682c415",
X"0c83c0d0",
X"33810682",
X"c8150c79",
X"5273519a",
X"f03f7351",
X"9b873f83",
X"c0800814",
X"53af7370",
X"81055534",
X"72bc150c",
X"83c0d152",
X"72519ad1",
X"3f83c0c8",
X"0882c015",
X"0c83c0de",
X"5280c014",
X"519abe3f",
X"78802e8d",
X"38735178",
X"2d83c080",
X"08802e99",
X"387782cc",
X"150c7580",
X"2e863873",
X"82cc170c",
X"7382d015",
X"ff195955",
X"5676802e",
X"9b3883c0",
X"c85283c2",
X"e85194ad",
X"3f83c080",
X"088a3883",
X"c0d13353",
X"72fed238",
X"78802e89",
X"3883c0c4",
X"0851fcb8",
X"3f83c0c4",
X"08537283",
X"c0800c8b",
X"3d0d04ff",
X"3d0d8052",
X"7351fdb5",
X"3f833d0d",
X"04f03d0d",
X"62705254",
X"f6903f83",
X"c0800874",
X"53873d70",
X"535555f6",
X"b03ff790",
X"3f7351d3",
X"3f635374",
X"5283c080",
X"0851fab8",
X"3f923d0d",
X"047183c0",
X"800c0480",
X"c01283c0",
X"800c0480",
X"3d0d7282",
X"c0110883",
X"c0800c51",
X"823d0d04",
X"803d0d72",
X"82cc1108",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"7282c411",
X"0883c080",
X"0c51823d",
X"0d04f93d",
X"0d7983c0",
X"98085757",
X"81772781",
X"96387688",
X"17082781",
X"8e387533",
X"5574822e",
X"89387483",
X"2eb33880",
X"fe397454",
X"761083fe",
X"06537688",
X"2a8c1708",
X"0552893d",
X"fc055199",
X"c33f83c0",
X"800880df",
X"38029d05",
X"33893d33",
X"71882b07",
X"565680d1",
X"39845476",
X"822b83fc",
X"06537687",
X"2a8c1708",
X"0552893d",
X"fc055199",
X"933f83c0",
X"8008b038",
X"029f0533",
X"0284059e",
X"05337198",
X"2b71902b",
X"07028c05",
X"9d053370",
X"882b7207",
X"8d3d3371",
X"80fffffe",
X"80060751",
X"52535758",
X"56833981",
X"557483c0",
X"800c893d",
X"0d04fb3d",
X"0d83c098",
X"08fe1988",
X"1208fe05",
X"55565480",
X"56747327",
X"8d388214",
X"33757129",
X"94160805",
X"57537583",
X"c0800c87",
X"3d0d04fc",
X"3d0d7652",
X"800b83c0",
X"98087033",
X"51525370",
X"832e0981",
X"06913895",
X"12339413",
X"3371982b",
X"71902b07",
X"5555519b",
X"12339a13",
X"3371882b",
X"07740783",
X"c0800c55",
X"863d0d04",
X"fc3d0d76",
X"83c09808",
X"55558075",
X"23881508",
X"5372812e",
X"88388814",
X"08732685",
X"388152b2",
X"39729038",
X"73335271",
X"832e0981",
X"06853890",
X"14085372",
X"8c160c72",
X"802e8d38",
X"7251fed6",
X"3f83c080",
X"08528539",
X"90140852",
X"7190160c",
X"80527183",
X"c0800c86",
X"3d0d04fa",
X"3d0d7883",
X"c0980871",
X"22810570",
X"83ffff06",
X"57545755",
X"73802e88",
X"38901508",
X"53728638",
X"835280e7",
X"39738f06",
X"527180da",
X"38811390",
X"160c8c15",
X"08537290",
X"38830b84",
X"17225752",
X"73762780",
X"c638bf39",
X"821633ff",
X"0574842a",
X"065271b2",
X"387251fc",
X"b13f8152",
X"7183c080",
X"0827a838",
X"835283c0",
X"80088817",
X"08279c38",
X"83c08008",
X"8c160c83",
X"c0800851",
X"fdbc3f83",
X"c0800890",
X"160c7375",
X"23805271",
X"83c0800c",
X"883d0d04",
X"f23d0d60",
X"6264585e",
X"5b753355",
X"74a02e09",
X"81068838",
X"81167044",
X"56ef3962",
X"70335656",
X"74af2e09",
X"81068438",
X"81164380",
X"0b881c0c",
X"62703351",
X"55749f26",
X"91387a51",
X"fdd23f83",
X"c0800856",
X"807d3483",
X"8139933d",
X"841c0870",
X"58595f8a",
X"55a07670",
X"81055834",
X"ff155574",
X"ff2e0981",
X"06ef3880",
X"705a5c88",
X"7f085f5a",
X"7b811d70",
X"81ff0660",
X"13703370",
X"af327030",
X"a0732771",
X"80250751",
X"51525b53",
X"5e575574",
X"80e73876",
X"ae2e0981",
X"06833881",
X"55787a27",
X"75075574",
X"802e9f38",
X"79883270",
X"3078ae32",
X"70307073",
X"079f2a53",
X"51575156",
X"75bb3888",
X"598b5aff",
X"ab397698",
X"2b557480",
X"25873881",
X"c9e01733",
X"57ff9f17",
X"55749926",
X"8938e017",
X"7081ff06",
X"58557881",
X"1a7081ff",
X"06721b53",
X"5b575576",
X"7534fef8",
X"397b1e7f",
X"0c805576",
X"a0268338",
X"8155748b",
X"19347a51",
X"fc823f83",
X"c0800880",
X"f538a054",
X"7a227085",
X"2b83e006",
X"5455901b",
X"08527c51",
X"93ce3f83",
X"c0800857",
X"83c08008",
X"8181387c",
X"33557480",
X"2e80f438",
X"8b1d3370",
X"832a7081",
X"06515656",
X"74b4388b",
X"7d841d08",
X"83c08008",
X"595b5b58",
X"ff185877",
X"ff2e9a38",
X"79708105",
X"5b337970",
X"81055b33",
X"71713152",
X"56567580",
X"2ee23886",
X"3975802e",
X"96387a51",
X"fbe53fff",
X"863983c0",
X"80085683",
X"c08008b6",
X"38833976",
X"56841b08",
X"8b113351",
X"5574a738",
X"8b1d3370",
X"842a7081",
X"06515656",
X"74893883",
X"56943981",
X"5690397c",
X"51fa943f",
X"83c08008",
X"881c0cfd",
X"81397583",
X"c0800c90",
X"3d0d04f8",
X"3d0d7a7c",
X"59578254",
X"83fe5377",
X"52765192",
X"933f8356",
X"83c08008",
X"80ec3881",
X"17337733",
X"71882b07",
X"56568256",
X"7482d4d5",
X"2e098106",
X"80d43875",
X"54b65377",
X"52765191",
X"e73f83c0",
X"80089838",
X"81173377",
X"3371882b",
X"0783c080",
X"08525656",
X"748182c6",
X"2eac3882",
X"5480d253",
X"77527651",
X"91be3f83",
X"c0800898",
X"38811733",
X"77337188",
X"2b0783c0",
X"80085256",
X"56748182",
X"c62e8338",
X"81567583",
X"c0800c8a",
X"3d0d04eb",
X"3d0d675a",
X"800b83c0",
X"980c90e0",
X"3f83c080",
X"08810655",
X"82567483",
X"ef387475",
X"538f3d70",
X"535759fe",
X"ca3f83c0",
X"800881ff",
X"06577681",
X"2e098106",
X"80d43890",
X"5483be53",
X"74527551",
X"90d23f83",
X"c0800880",
X"c9388f3d",
X"33557480",
X"2e80c938",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"0770587b",
X"575e525e",
X"575957fd",
X"ee3f83c0",
X"800881ff",
X"06577683",
X"2e098106",
X"86388156",
X"82f23976",
X"802e8638",
X"865682e8",
X"39a4548d",
X"53785275",
X"518fe93f",
X"815683c0",
X"800882d4",
X"3802be05",
X"33028405",
X"bd053371",
X"882b0759",
X"5d77ab38",
X"0280ce05",
X"33028405",
X"80cd0533",
X"71982b71",
X"902b0797",
X"3d337088",
X"2b720702",
X"940580cb",
X"05337107",
X"54525e57",
X"595602b7",
X"05337871",
X"29028805",
X"b6053302",
X"8c05b505",
X"3371882b",
X"07701d70",
X"7f8c050c",
X"5f595759",
X"5d8e3d33",
X"821b3402",
X"b9053390",
X"3d337188",
X"2b075a5c",
X"78841b23",
X"02bb0533",
X"028405ba",
X"05337188",
X"2b07565c",
X"74ab3802",
X"80ca0533",
X"02840580",
X"c9053371",
X"982b7190",
X"2b07963d",
X"3370882b",
X"72070294",
X"0580c705",
X"33710751",
X"5253575e",
X"5c747631",
X"78317984",
X"2a903d33",
X"54717131",
X"53565681",
X"91cf3f83",
X"c0800882",
X"0570881c",
X"0c83c080",
X"08e08a05",
X"56567483",
X"dffe2683",
X"38825783",
X"fff67627",
X"85388357",
X"89398656",
X"76802e80",
X"db38767a",
X"3476832e",
X"098106b0",
X"380280d6",
X"05330284",
X"0580d505",
X"3371982b",
X"71902b07",
X"993d3370",
X"882b7207",
X"02940580",
X"d3053371",
X"077f9005",
X"0c525e57",
X"58568639",
X"771b901b",
X"0c841a22",
X"8c1b0819",
X"71842a05",
X"941c0c5d",
X"800b811b",
X"347983c0",
X"980c8056",
X"7583c080",
X"0c973d0d",
X"04e93d0d",
X"83c09808",
X"56855475",
X"802e8182",
X"38800b81",
X"1734993d",
X"e011466a",
X"548a3d70",
X"5458ec05",
X"51f6e53f",
X"83c08008",
X"5483c080",
X"0880df38",
X"893d3354",
X"73802e91",
X"3802ab05",
X"3370842a",
X"81065155",
X"74802e86",
X"38835480",
X"c1397651",
X"f4893f83",
X"c08008a0",
X"170c02bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"3371079c",
X"1c0c5278",
X"981b0c53",
X"56595781",
X"0b811734",
X"74547383",
X"c0800c99",
X"3d0d04f5",
X"3d0d7d7f",
X"617283c0",
X"98085a5d",
X"5d595c80",
X"7b0c8557",
X"75802e81",
X"e0388116",
X"33810655",
X"84577480",
X"2e81d238",
X"91397481",
X"17348639",
X"800b8117",
X"34815781",
X"c0399c16",
X"08981708",
X"31557478",
X"27833874",
X"5877802e",
X"81a93898",
X"16087083",
X"ff065657",
X"7480cf38",
X"821633ff",
X"0577892a",
X"067081ff",
X"065a5578",
X"a0387687",
X"38a01608",
X"558d39a4",
X"160851f0",
X"e93f83c0",
X"80085581",
X"7527ffa8",
X"3874a417",
X"0ca41608",
X"51f2833f",
X"83c08008",
X"5583c080",
X"08802eff",
X"893883c0",
X"800819a8",
X"170c9816",
X"0883ff06",
X"84807131",
X"51557775",
X"27833877",
X"557483ff",
X"ff065498",
X"160883ff",
X"0653a816",
X"08527957",
X"7b83387b",
X"5776518a",
X"8f3f83c0",
X"8008fed0",
X"38981608",
X"1598170c",
X"741a7876",
X"317c0817",
X"7d0c595a",
X"fed33980",
X"577683c0",
X"800c8d3d",
X"0d04fa3d",
X"0d7883c0",
X"98085556",
X"85557380",
X"2e81e338",
X"81143381",
X"06538455",
X"72802e81",
X"d5389c14",
X"08537276",
X"27833872",
X"56981408",
X"57800b98",
X"150c7580",
X"2e81b938",
X"82143370",
X"892b5653",
X"76802eb7",
X"387452ff",
X"1651818c",
X"d03f83c0",
X"8008ff18",
X"76547053",
X"5853818c",
X"c03f83c0",
X"80087326",
X"96387430",
X"70780670",
X"98170c77",
X"7131a417",
X"08525851",
X"538939a0",
X"140870a4",
X"160c5374",
X"7627b938",
X"7251eed6",
X"3f83c080",
X"0853810b",
X"83c08008",
X"278b3888",
X"140883c0",
X"80082688",
X"38800b81",
X"1534b039",
X"83c08008",
X"a4150c98",
X"14081598",
X"150c7575",
X"3156c439",
X"98140816",
X"7098160c",
X"735256ef",
X"c53f83c0",
X"80088c38",
X"83c08008",
X"81153481",
X"55943982",
X"1433ff05",
X"76892a06",
X"83c08008",
X"05a8150c",
X"80557483",
X"c0800c88",
X"3d0d04ef",
X"3d0d6356",
X"855583c0",
X"9808802e",
X"80d23893",
X"3df40584",
X"170c6453",
X"883d7053",
X"765257f1",
X"cf3f83c0",
X"80085583",
X"c08008b4",
X"38883d33",
X"5473802e",
X"a13802a7",
X"05337084",
X"2a708106",
X"51555583",
X"5573802e",
X"97387651",
X"eef53f83",
X"c0800888",
X"170c7551",
X"efa63f83",
X"c0800855",
X"7483c080",
X"0c933d0d",
X"04e43d0d",
X"6ea13d08",
X"405e8556",
X"83c09808",
X"802e8485",
X"389e3df4",
X"05841f0c",
X"7e98387d",
X"51eef53f",
X"83c08008",
X"5683ee39",
X"814181f6",
X"39834181",
X"f139933d",
X"7f960541",
X"59807f82",
X"95055e56",
X"756081ff",
X"05348341",
X"901e0876",
X"2e81d338",
X"a0547d22",
X"70852b83",
X"e0065458",
X"901e0852",
X"78518698",
X"3f83c080",
X"084183c0",
X"8008ffb8",
X"3878335c",
X"7b802eff",
X"b4388b19",
X"3370bf06",
X"71810652",
X"43557480",
X"2e80de38",
X"7b81bf06",
X"55748f24",
X"80d3389a",
X"19335574",
X"80cb38f3",
X"1d70585d",
X"8156758b",
X"2e098106",
X"85388e56",
X"8b39759a",
X"2e098106",
X"83389c56",
X"75197070",
X"81055233",
X"7133811a",
X"821a5f5b",
X"525b5574",
X"86387977",
X"34853980",
X"df773477",
X"7b57577a",
X"a02e0981",
X"06c03881",
X"567b81e5",
X"32703070",
X"9f2a5151",
X"557bae2e",
X"93387480",
X"2e8e3861",
X"832a7081",
X"06515574",
X"802e9738",
X"7d51eddf",
X"3f83c080",
X"084183c0",
X"80088738",
X"901e08fe",
X"af388060",
X"3475802e",
X"88387c52",
X"7f5183a5",
X"3f60802e",
X"8638800b",
X"901f0c60",
X"5660832e",
X"85386081",
X"d038891f",
X"57901e08",
X"802e81a8",
X"38805675",
X"19703351",
X"5574a02e",
X"a0387485",
X"2e098106",
X"843881e5",
X"55747770",
X"81055934",
X"81167081",
X"ff065755",
X"877627d7",
X"38881933",
X"5574a02e",
X"a938ae77",
X"70810559",
X"34885675",
X"19703351",
X"5574a02e",
X"95387477",
X"70810559",
X"34811670",
X"81ff0657",
X"558a7627",
X"e2388b19",
X"337f8805",
X"349f1933",
X"9e1a3371",
X"982b7190",
X"2b079d1c",
X"3370882b",
X"72079c1e",
X"33710764",
X"0c52991d",
X"33981e33",
X"71882b07",
X"53515357",
X"5956747f",
X"84052397",
X"1933961a",
X"3371882b",
X"07565674",
X"7f860523",
X"8077347d",
X"51ebf03f",
X"83c08008",
X"83327030",
X"7072079f",
X"2c83c080",
X"08065256",
X"56961f33",
X"55748a38",
X"891f5296",
X"1f5181b1",
X"3f7583c0",
X"800c9e3d",
X"0d04fd3d",
X"0d757753",
X"54733351",
X"70893871",
X"33517080",
X"2ea13873",
X"33723352",
X"53727127",
X"8538ff51",
X"94397073",
X"27853881",
X"518b3981",
X"14811353",
X"54d33980",
X"517083c0",
X"800c853d",
X"0d04fd3d",
X"0d757754",
X"54723370",
X"81ff0652",
X"5270802e",
X"a3387181",
X"ff068114",
X"ffbf1253",
X"54527099",
X"268938a0",
X"127081ff",
X"06535171",
X"74708105",
X"5634d239",
X"80743485",
X"3d0d04ff",
X"bd3d0d80",
X"c63d0852",
X"a53d7052",
X"54ffb33f",
X"80c73d08",
X"52853d70",
X"5253ffa6",
X"3f725273",
X"51fedf3f",
X"80c53d0d",
X"04fe3d0d",
X"74765353",
X"71708105",
X"53335170",
X"73708105",
X"553470f0",
X"38843d0d",
X"04fe3d0d",
X"74528072",
X"33525370",
X"732e8d38",
X"81128114",
X"71335354",
X"5270f538",
X"7283c080",
X"0c843d0d",
X"04fc3d0d",
X"76557483",
X"c3a8082e",
X"af388053",
X"745187c1",
X"3f83c080",
X"0881ff06",
X"ff147081",
X"ff067230",
X"709f2a51",
X"52555354",
X"72802e84",
X"3871dd38",
X"73fe3874",
X"83c3a80c",
X"863d0d04",
X"ff3d0dff",
X"0b83c3a8",
X"0c84a53f",
X"81518785",
X"3f83c080",
X"0881ff06",
X"5271ee38",
X"81d33f71",
X"83c0800c",
X"833d0d04",
X"fc3d0d76",
X"028405a2",
X"05220288",
X"05a60522",
X"7a545555",
X"55ff823f",
X"72802ea0",
X"3883c3bc",
X"14337570",
X"81055734",
X"81147083",
X"ffff06ff",
X"157083ff",
X"ff065652",
X"5552dd39",
X"800b83c0",
X"800c863d",
X"0d04fc3d",
X"0d76787a",
X"11565355",
X"80537174",
X"2e933872",
X"15517033",
X"83c3bc13",
X"34811281",
X"145452ea",
X"39800b83",
X"c0800c86",
X"3d0d04fd",
X"3d0d9054",
X"83c3a808",
X"5186f43f",
X"83c08008",
X"81ff06ff",
X"15713071",
X"30707307",
X"9f2a729f",
X"2a065255",
X"52555372",
X"db38853d",
X"0d04803d",
X"0d83c3b4",
X"081083c3",
X"ac080790",
X"80a80c82",
X"3d0d0480",
X"0b83c3b4",
X"0ce43f04",
X"810b83c3",
X"b40cdb3f",
X"04ed3f04",
X"7183c3b0",
X"0c04803d",
X"0d8051f4",
X"3f810b83",
X"c3b40c81",
X"0b83c3ac",
X"0cffbb3f",
X"823d0d04",
X"803d0d72",
X"30707407",
X"802583c3",
X"ac0c51ff",
X"a53f823d",
X"0d04803d",
X"0d028b05",
X"339080a4",
X"0c9080a8",
X"08708106",
X"515170f5",
X"389080a4",
X"087081ff",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d81ff51",
X"d13f83c0",
X"800881ff",
X"0683c080",
X"0c823d0d",
X"04803d0d",
X"73902b73",
X"079080b4",
X"0c823d0d",
X"0404fb3d",
X"0d780284",
X"059f0533",
X"70982b55",
X"57557280",
X"259b3875",
X"80ff0656",
X"805280f7",
X"51e03f83",
X"c0800881",
X"ff065473",
X"812680ff",
X"388051fe",
X"e73fffa2",
X"3f8151fe",
X"df3fff9a",
X"3f7551fe",
X"ed3f7498",
X"2a51fee6",
X"3f74902a",
X"7081ff06",
X"5253feda",
X"3f74882a",
X"7081ff06",
X"5253fece",
X"3f7481ff",
X"0651fec6",
X"3f815575",
X"80c02e09",
X"81068638",
X"8195558d",
X"397580c8",
X"2e098106",
X"84388187",
X"557451fe",
X"a53f8a55",
X"fec83f83",
X"c0800881",
X"ff067098",
X"2b545472",
X"80258c38",
X"ff157081",
X"ff065653",
X"74e23873",
X"83c0800c",
X"873d0d04",
X"fa3d0dfd",
X"c53f8051",
X"fdda3f8a",
X"54fe933f",
X"ff147081",
X"ff065553",
X"73f33873",
X"74535580",
X"c051fea6",
X"3f83c080",
X"0881ff06",
X"5473812e",
X"09810682",
X"9f3883aa",
X"5280c851",
X"fe8c3f83",
X"c0800881",
X"ff065372",
X"812e0981",
X"0681a838",
X"7454873d",
X"74115456",
X"fdc83f83",
X"c0800873",
X"34811470",
X"81ff0655",
X"53837427",
X"e538029a",
X"05335372",
X"812e0981",
X"0681d938",
X"029b0533",
X"5380ce90",
X"547281aa",
X"2e8d3881",
X"c73980e4",
X"518ad63f",
X"ff145473",
X"802e81b8",
X"38820a52",
X"81e951fd",
X"a53f83c0",
X"800881ff",
X"065372de",
X"38725280",
X"fa51fd92",
X"3f83c080",
X"0881ff06",
X"53728190",
X"38725473",
X"1653fcd6",
X"3f83c080",
X"08733481",
X"147081ff",
X"06555383",
X"7427e838",
X"873d3370",
X"862a7081",
X"06515454",
X"8c557280",
X"e3388455",
X"80de3974",
X"5281e951",
X"fccc3f83",
X"c0800881",
X"ff065382",
X"5581e956",
X"81732786",
X"38735580",
X"c15680ce",
X"90548a39",
X"80e45189",
X"c83fff14",
X"5473802e",
X"a9388052",
X"7551fc9a",
X"3f83c080",
X"0881ff06",
X"5372e138",
X"84805280",
X"d051fc86",
X"3f83c080",
X"0881ff06",
X"5372802e",
X"83388055",
X"7483c3b8",
X"348051fb",
X"873ffbc2",
X"3f883d0d",
X"04fb3d0d",
X"7754800b",
X"83c3b833",
X"70832a70",
X"81065155",
X"57557275",
X"2e098106",
X"85387389",
X"2b547352",
X"80d151fb",
X"bd3f83c0",
X"800881ff",
X"065372bd",
X"3882b8c0",
X"54fb833f",
X"83c08008",
X"81ff0653",
X"7281ff2e",
X"09810689",
X"38ff1454",
X"73e7389f",
X"397281fe",
X"2e098106",
X"963883c7",
X"bc5283c3",
X"bc51faed",
X"3ffad33f",
X"fad03f83",
X"39815580",
X"51fa893f",
X"fac43f74",
X"81ff0683",
X"c0800c87",
X"3d0d04fb",
X"3d0d7783",
X"c3bc5654",
X"8151f9ec",
X"3f83c3b8",
X"3370832a",
X"70810651",
X"54567285",
X"3873892b",
X"54735280",
X"d851fab6",
X"3f83c080",
X"0881ff06",
X"537280e4",
X"3881ff51",
X"f9d43f81",
X"fe51f9ce",
X"3f848053",
X"74708105",
X"563351f9",
X"c13fff13",
X"7083ffff",
X"06515372",
X"eb387251",
X"f9b03f72",
X"51f9ab3f",
X"f9d03f83",
X"c080089f",
X"0653a788",
X"5472852e",
X"8c389939",
X"80e45187",
X"803fff14",
X"54f9b33f",
X"83c08008",
X"81ff2e84",
X"3873e938",
X"8051f8e4",
X"3ff99f3f",
X"800b83c0",
X"800c873d",
X"0d047183",
X"c7c00c88",
X"80800b83",
X"c7bc0c84",
X"80800b83",
X"c7c40c04",
X"f03d0d83",
X"80805683",
X"c7c00816",
X"83c7bc08",
X"17565474",
X"33743483",
X"c7c40816",
X"54807434",
X"81165675",
X"8380a02e",
X"098106db",
X"3883d080",
X"5683c7c0",
X"081683c7",
X"bc081756",
X"54743374",
X"3483c7c4",
X"08165480",
X"74348116",
X"567583d0",
X"902e0981",
X"06db3883",
X"a8805683",
X"c7c00816",
X"83c7bc08",
X"17565474",
X"33743483",
X"c7c40816",
X"54807434",
X"81165675",
X"83a8902e",
X"098106db",
X"38805683",
X"c7c00816",
X"83c7c408",
X"17555573",
X"33753481",
X"16567581",
X"80802e09",
X"8106e438",
X"87943f89",
X"3d58a253",
X"81cbe052",
X"775180ff",
X"e33f8057",
X"8c805683",
X"c7c40816",
X"77195555",
X"73337534",
X"81168118",
X"585676a2",
X"2e098106",
X"e638860b",
X"87a88334",
X"800b87a8",
X"8234800b",
X"87809a34",
X"af0b8780",
X"9634bf0b",
X"87809734",
X"800b8780",
X"98349f0b",
X"87809934",
X"800b8780",
X"9b34f80b",
X"87a88934",
X"7687a880",
X"34820b87",
X"d08f3482",
X"0b87a881",
X"34923d0d",
X"04fe3d0d",
X"805383c7",
X"c4081383",
X"c7c00814",
X"52527033",
X"72348113",
X"53728180",
X"802e0981",
X"06e43883",
X"80805383",
X"c7c40813",
X"83c7c008",
X"14525270",
X"33723481",
X"13537283",
X"80a02e09",
X"8106e438",
X"83d08053",
X"83c7c408",
X"1383c7c0",
X"08145252",
X"70337234",
X"81135372",
X"83d0902e",
X"098106e4",
X"3883a880",
X"5383c7c4",
X"081383c7",
X"c0081452",
X"52703372",
X"34811353",
X"7283a890",
X"2e098106",
X"e438843d",
X"0d04803d",
X"0d908090",
X"08810683",
X"c0800c82",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe067607",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"812c8106",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fd06",
X"76100772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087082",
X"2cbf0683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fe8306",
X"76822b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"882c8706",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f1ff",
X"0676882b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"708b2cbf",
X"0683c080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870f8",
X"8fff0676",
X"8b2b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087091",
X"2cbf0683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fc87ff",
X"ff067691",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870992c",
X"810683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"ffbf0a06",
X"76992b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80800870",
X"882c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"70892c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708a2c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708b",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8c2cbf06",
X"83c0800c",
X"51823d0d",
X"04fe3d0d",
X"7481e629",
X"872a9080",
X"a00c843d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"81055434",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727084",
X"05540cff",
X"1151f039",
X"843d0d04",
X"fe3d0d81",
X"80805380",
X"5288800a",
X"51ffb33f",
X"a0805380",
X"5282800a",
X"51c73f84",
X"3d0d0480",
X"3d0d8151",
X"fbfd3f72",
X"802e9038",
X"8051fdff",
X"3fce3f81",
X"d2dc3351",
X"fdf53f81",
X"51fc8e3f",
X"8051fc89",
X"3f8051fb",
X"da3f823d",
X"0d04fd3d",
X"0d755280",
X"5480ff72",
X"25883881",
X"0bff8013",
X"5354ffbf",
X"12517099",
X"268638e0",
X"12529e39",
X"ff9f1251",
X"99712795",
X"38d012e0",
X"13705454",
X"51897127",
X"88388f73",
X"27833880",
X"5273802e",
X"85388180",
X"12527181",
X"ff0683c0",
X"800c853d",
X"0d04803d",
X"0d84d8c0",
X"51807170",
X"81055334",
X"7084e0c0",
X"2e098106",
X"f038823d",
X"0d04fe3d",
X"0d029705",
X"3351ff86",
X"3f83c080",
X"0881ff06",
X"83c7cc08",
X"54528073",
X"249b3883",
X"c88c0813",
X"7283c890",
X"08075353",
X"71733483",
X"c7cc0881",
X"0583c7cc",
X"0c843d0d",
X"04fa3d0d",
X"82800a1b",
X"55805788",
X"3dfc0554",
X"79537452",
X"7851cbc8",
X"3f883d0d",
X"04fe3d0d",
X"83c7e408",
X"527451d2",
X"ac3f83c0",
X"80088c38",
X"76537552",
X"83c7e408",
X"51c73f84",
X"3d0d04fe",
X"3d0d83c7",
X"e4085375",
X"527451cc",
X"eb3f83c0",
X"80088d38",
X"77537652",
X"83c7e408",
X"51ffa23f",
X"843d0d04",
X"fd3d0d83",
X"c7e40851",
X"cbdf3f83",
X"c0800890",
X"802e0981",
X"06ad3880",
X"5483c180",
X"805383c0",
X"80085283",
X"c7e40851",
X"fef33f87",
X"c1808014",
X"3387c190",
X"80153481",
X"14547390",
X"802e0981",
X"06e93885",
X"3d0d0481",
X"d0ac0b83",
X"c0800c04",
X"fc3d0d76",
X"5473902e",
X"80ff3873",
X"90248e38",
X"73842e98",
X"3873862e",
X"a63882b9",
X"3973932e",
X"81953873",
X"942e81cf",
X"3882aa39",
X"81808053",
X"82808052",
X"83c7e008",
X"51fe923f",
X"82b53980",
X"54818080",
X"5380c080",
X"5283c7e0",
X"0851fdfd",
X"3f828080",
X"5380c080",
X"5283c7e0",
X"0851fded",
X"3f848180",
X"80143384",
X"81c08015",
X"34848280",
X"80143384",
X"82c08015",
X"34811454",
X"7380c080",
X"2e098106",
X"dc3881eb",
X"39828080",
X"53818080",
X"5283c7e0",
X"0851fdb5",
X"3f805484",
X"82808014",
X"33848180",
X"80153481",
X"14547381",
X"80802e09",
X"8106e838",
X"81bd3981",
X"80805380",
X"c0805283",
X"c7e00851",
X"fd873f80",
X"55848180",
X"80155473",
X"338481c0",
X"80163473",
X"33848280",
X"80163473",
X"338482c0",
X"80163481",
X"15557480",
X"c0802e09",
X"8106d638",
X"80fd3981",
X"808053a0",
X"805283c7",
X"e00851fc",
X"c83f8055",
X"84818080",
X"15547333",
X"8481a080",
X"16347333",
X"8481c080",
X"16347333",
X"8481e080",
X"16347333",
X"84828080",
X"16347333",
X"8482a080",
X"16347333",
X"8482c080",
X"16347333",
X"8482e080",
X"16348115",
X"5574a080",
X"2e098106",
X"ffb6389f",
X"39fb9f3f",
X"800b83c7",
X"cc0c800b",
X"83c8900c",
X"81d0b051",
X"c3fc3f81",
X"b78dc051",
X"f9933f86",
X"3d0d04fc",
X"3d0d7670",
X"5255cf81",
X"3f83c080",
X"08548153",
X"83c08008",
X"80c43874",
X"51cec43f",
X"83c08008",
X"81d0cc53",
X"83c08008",
X"5253ffb4",
X"b13f83c0",
X"8008a338",
X"81d0d052",
X"7251ffb4",
X"a13f83c0",
X"80089338",
X"81d0d452",
X"7251ffb4",
X"913f83c0",
X"8008802e",
X"83388154",
X"73537283",
X"c0800c86",
X"3d0d04f1",
X"3d0d80d5",
X"d70b83c0",
X"b80c83c7",
X"e00851ff",
X"b5c33f83",
X"c7e00851",
X"c4ad3fff",
X"0b81d0d0",
X"5383c080",
X"085256ff",
X"b3d03f83",
X"c0800880",
X"2e9e3880",
X"58913ddc",
X"11555590",
X"53f01552",
X"83c7e008",
X"51c6893f",
X"02b70533",
X"5681a239",
X"83c7e008",
X"51c6e63f",
X"83c08008",
X"5783c080",
X"08828080",
X"2e098106",
X"83388456",
X"83c08008",
X"8180802e",
X"09810680",
X"df38805b",
X"805a8059",
X"f9983f80",
X"0b83c7cc",
X"0c800b83",
X"c8900c81",
X"d0d851c1",
X"f53f80d0",
X"0b83c7cc",
X"0c81d0e8",
X"51c1e73f",
X"80f80b83",
X"c7cc0c81",
X"d0fc51c1",
X"d93f7580",
X"25a23880",
X"52893d70",
X"52558a8d",
X"3f835274",
X"518a863f",
X"78557480",
X"25833890",
X"56807525",
X"dd388656",
X"7680c080",
X"2e098106",
X"85389356",
X"8c3976a0",
X"802e0981",
X"06833894",
X"567551fa",
X"af3f913d",
X"0d04f73d",
X"0d805980",
X"58805780",
X"705656f8",
X"913f800b",
X"83c7cc0c",
X"800b83c8",
X"900c81d1",
X"9051c0ee",
X"3f81800b",
X"83c8900c",
X"81d19451",
X"c0e03f80",
X"d00b83c7",
X"cc0c7430",
X"70760780",
X"2570872b",
X"83c8900c",
X"5153f397",
X"3f83c080",
X"085281d1",
X"9c51c0ba",
X"3f80f80b",
X"83c7cc0c",
X"74813270",
X"30707207",
X"80257087",
X"2b83c890",
X"0c515454",
X"f9ad3f83",
X"c0800852",
X"81d1a851",
X"c0903f81",
X"a00b83c7",
X"cc0c7482",
X"32703070",
X"72078025",
X"70872b83",
X"c8900c51",
X"5483c7e4",
X"085254c1",
X"aa3f83c0",
X"80085281",
X"d1b051ff",
X"bfe03f81",
X"c80b83c7",
X"cc0c7483",
X"32703070",
X"72078025",
X"70872b83",
X"c8900c51",
X"5483c7e0",
X"085254c0",
X"fa3f81d1",
X"b85383c0",
X"8008802e",
X"8e3883c7",
X"e00851c0",
X"e63f83c0",
X"80085372",
X"5281d1c0",
X"51ffbf9a",
X"3f81f00b",
X"83c7cc0c",
X"74843270",
X"30707207",
X"80257087",
X"2b83c890",
X"0c515581",
X"d1c85253",
X"ffbef73f",
X"868da051",
X"f48f3f80",
X"52873d70",
X"525387a9",
X"3f835272",
X"5187a23f",
X"77155574",
X"80258538",
X"80559039",
X"84752585",
X"38845587",
X"39748426",
X"81a13874",
X"842981cc",
X"84055372",
X"0804f187",
X"3f83c080",
X"08775553",
X"73812e09",
X"81068938",
X"83c08008",
X"10539039",
X"73ff2e09",
X"81068838",
X"83c08008",
X"812c5390",
X"73258538",
X"90538839",
X"72802483",
X"38815372",
X"51f0e13f",
X"80d539f0",
X"f33f83c0",
X"80081753",
X"72802585",
X"38805388",
X"39877325",
X"83388753",
X"7251f0ed",
X"3fb53976",
X"86387880",
X"2ead3883",
X"c0b40883",
X"c0b00c8b",
X"df0b83c0",
X"b80c83c7",
X"e40851ff",
X"b0833ff5",
X"ff3f9039",
X"78802e8b",
X"38faa03f",
X"81538c39",
X"78873875",
X"802efc9b",
X"38805372",
X"83c0800c",
X"8b3d0d04",
X"ff3d0d83",
X"c7fc5180",
X"df813f83",
X"c7ec5180",
X"def93ff1",
X"b33f83c0",
X"8008802e",
X"86388051",
X"80da39f1",
X"b83f83c0",
X"800880ce",
X"38f1d83f",
X"83c08008",
X"802eaa38",
X"8151eee7",
X"3febad3f",
X"800b83c7",
X"cc0cfbba",
X"3f83c080",
X"0852ff0b",
X"83c7cc0c",
X"edb33f71",
X"a1387151",
X"eec53f9f",
X"39f18f3f",
X"83c08008",
X"802e9438",
X"8151eeb3",
X"3feaf93f",
X"f9913fed",
X"903f8151",
X"f2a13f83",
X"3d0d04fe",
X"3d0d8052",
X"83c7fc51",
X"80ceb83f",
X"815283c7",
X"ec5180ce",
X"ae3f8280",
X"80538052",
X"81818080",
X"51f19b3f",
X"80c08053",
X"80528481",
X"808051f1",
X"ac3f9080",
X"80528684",
X"808051c1",
X"ad3f83c0",
X"8008a238",
X"81d2ec51",
X"c5f13f83",
X"c7e40853",
X"81d1d052",
X"83c08008",
X"51c0d13f",
X"83c08008",
X"8438f3f4",
X"3f8151f1",
X"b23ffe90",
X"3ffc3983",
X"c08c0802",
X"83c08c0c",
X"fb3d0d02",
X"81d1dc0b",
X"83c0b40c",
X"81d0d40b",
X"83c0ac0c",
X"81d0d00b",
X"83c0bc0c",
X"83c08c08",
X"fc050c80",
X"0b83c7d0",
X"0b83c08c",
X"08f8050c",
X"83c08c08",
X"f4050cff",
X"bfb03f83",
X"c0800886",
X"05fc0683",
X"c08c08f0",
X"050c0283",
X"c08c08f0",
X"0508310d",
X"833d7083",
X"c08c08f8",
X"05087084",
X"0583c08c",
X"08f8050c",
X"0c51ffbb",
X"f83f83c0",
X"8c08f405",
X"08810583",
X"c08c08f4",
X"050c83c0",
X"8c08f405",
X"08872e09",
X"8106ffab",
X"38869480",
X"8051e8c6",
X"3fff0b83",
X"c7cc0c80",
X"0b83c890",
X"0c84d8c0",
X"0b83c88c",
X"0c8151eb",
X"fa3f8151",
X"ec9f3f80",
X"51ec9a3f",
X"8151ecc0",
X"3f8151ed",
X"953f8251",
X"ece33f80",
X"51edb93f",
X"8051ede3",
X"3f80d0f2",
X"528051ff",
X"b9b13ffd",
X"aa3f83c0",
X"8c08fc05",
X"080d800b",
X"83c0800c",
X"873d0d83",
X"c08c0c04",
X"fc3d0d76",
X"5580750c",
X"800b8416",
X"0c800b88",
X"160c83c7",
X"fc5180db",
X"823f83c7",
X"ec5180da",
X"fa3f87d0",
X"893387d0",
X"8f337082",
X"2a708106",
X"70307072",
X"07700970",
X"9f2c7706",
X"9e065451",
X"51565151",
X"5454ede4",
X"3f807398",
X"06535471",
X"882e0981",
X"06833881",
X"54719832",
X"70307080",
X"25767131",
X"84190c51",
X"51528073",
X"86065354",
X"71822e09",
X"81068338",
X"81547186",
X"32703070",
X"80257671",
X"31780c51",
X"51527294",
X"32703070",
X"80258818",
X"0c515283",
X"c0800880",
X"2e80c238",
X"83c08008",
X"812a7081",
X"0683c080",
X"08810631",
X"84170c52",
X"83c08008",
X"832a83c0",
X"8008822a",
X"71810671",
X"81063177",
X"0c535383",
X"c0800884",
X"2a810688",
X"160c83c0",
X"8008852a",
X"81068c16",
X"0c863d0d",
X"04fe3d0d",
X"74765452",
X"7151fe90",
X"3f72812e",
X"a2388173",
X"268d3872",
X"822eab38",
X"72832e9f",
X"38e63971",
X"08e23884",
X"1208dd38",
X"881208d8",
X"38a03988",
X"1208812e",
X"098106cc",
X"38943988",
X"1208812e",
X"8d387108",
X"89388412",
X"08802eff",
X"b738843d",
X"0d04fb3d",
X"0d780284",
X"059f0533",
X"5556800b",
X"81ce8456",
X"5381732b",
X"74065271",
X"802e8338",
X"81527470",
X"82055622",
X"7073902b",
X"0790809c",
X"0c518113",
X"5372882e",
X"098106d9",
X"38805383",
X"c8981333",
X"517081ff",
X"2eb23870",
X"1081cca4",
X"05702255",
X"51807317",
X"70337010",
X"81cca405",
X"70225151",
X"51525273",
X"712e9138",
X"81125271",
X"862e0981",
X"06f13873",
X"90809c0c",
X"81135372",
X"862e0981",
X"06ffb838",
X"80537216",
X"70335151",
X"7081ff2e",
X"94387010",
X"81cca405",
X"70227084",
X"80800790",
X"809c0c51",
X"51811353",
X"72862e09",
X"8106d738",
X"80537216",
X"51703383",
X"c8981434",
X"81135372",
X"862e0981",
X"06ec3887",
X"3d0d0404",
X"ff3d0d74",
X"0284058f",
X"05335252",
X"70883871",
X"9080940c",
X"8e397081",
X"2e098106",
X"86387190",
X"80980c83",
X"3d0d04fb",
X"3d0d029f",
X"05337998",
X"2b70982c",
X"7c982b70",
X"982c83c8",
X"b4157033",
X"70982b70",
X"982c5158",
X"5c5a5155",
X"51545470",
X"732e0981",
X"06943883",
X"c8941433",
X"70982b70",
X"982c5152",
X"5670722e",
X"b1387275",
X"347183c8",
X"94153483",
X"c8953383",
X"c8b53371",
X"982b7190",
X"2b0783c8",
X"94337088",
X"2b720783",
X"c8b43371",
X"079080b8",
X"0c525953",
X"5452873d",
X"0d04fe3d",
X"0d748111",
X"33713371",
X"882b0783",
X"c0800c53",
X"51843d0d",
X"0483c8a0",
X"3383c080",
X"0c04f53d",
X"0d02bb05",
X"33028405",
X"bf053302",
X"880580c3",
X"0533028c",
X"0580c605",
X"22665c5a",
X"5e5c567a",
X"557b5489",
X"53a1527d",
X"5180d0c0",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8d3d0d04",
X"83c08c08",
X"0283c08c",
X"0cf53d0d",
X"83c08c08",
X"88050883",
X"c08c088f",
X"053383c0",
X"8c089205",
X"22028c05",
X"73900583",
X"c08c08e8",
X"050c83c0",
X"8c08f805",
X"0c83c08c",
X"08f0050c",
X"83c08c08",
X"ec050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"f0050883",
X"c08c08e0",
X"050c83c0",
X"8c08fc05",
X"0c83c08c",
X"08f00508",
X"89278a38",
X"890b83c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"860587ff",
X"fc0683c0",
X"8c08e005",
X"0c0283c0",
X"8c08e005",
X"08310d85",
X"3d705583",
X"c08c08ec",
X"05085483",
X"c08c08f0",
X"05085383",
X"c08c08f4",
X"05085283",
X"c08c08e4",
X"050c80d9",
X"f23f83c0",
X"800881ff",
X"0683c08c",
X"08e40508",
X"83c08c08",
X"ec050c83",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08802e8c",
X"3883c08c",
X"08f80508",
X"0d89c839",
X"83c08c08",
X"f0050880",
X"2e89a638",
X"83c08c08",
X"ec050881",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"842ea938",
X"840b83c0",
X"8c08e005",
X"082588c7",
X"3883c08c",
X"08e00508",
X"852e859b",
X"3883c08c",
X"08e00508",
X"a12e87ad",
X"3888ac39",
X"800b83c0",
X"8c08ec05",
X"08850533",
X"83c08c08",
X"e0050c83",
X"c08c08fc",
X"050c83c0",
X"8c08e005",
X"08832e09",
X"81068883",
X"3883c08c",
X"08e80508",
X"81053383",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08812687",
X"e638810b",
X"83c08c08",
X"e0050880",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08fc050c",
X"83c08c08",
X"ec050882",
X"053383c0",
X"8c08e005",
X"08870534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088b0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08e005",
X"088c0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088d0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08e005",
X"088e0523",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088a0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"08057094",
X"0508fcff",
X"ff067194",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08ec0508",
X"86053383",
X"c08c08e0",
X"050c83c0",
X"8c08f405",
X"0c83c08c",
X"08e00508",
X"83c08c08",
X"fc05082e",
X"098106b6",
X"3883c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08fc0508",
X"83c08c08",
X"e005088b",
X"053483c0",
X"8c08ec05",
X"08870533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508812e",
X"8f3883c0",
X"8c08e005",
X"08822eb7",
X"38848c39",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"820b83c0",
X"8c08e005",
X"088a0534",
X"83d93983",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c83",
X"c08c08fc",
X"050883c0",
X"8c08e005",
X"088a0534",
X"83a13983",
X"c08c08fc",
X"0508802e",
X"83953883",
X"c08c08ec",
X"05088305",
X"33830683",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08832e09",
X"810682f3",
X"3883c08c",
X"08ec0508",
X"82053370",
X"982b83c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"83c08c08",
X"e0050880",
X"2582cc38",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"83c08c08",
X"ec050886",
X"053383c0",
X"8c08e005",
X"0880d605",
X"3483c08c",
X"08e00508",
X"840583c0",
X"8c08ec05",
X"08820533",
X"8f0683c0",
X"8c08e405",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"e4050883",
X"c08c08e0",
X"05083483",
X"c08c08ec",
X"05088405",
X"3383c08c",
X"08e00508",
X"81053480",
X"0b83c08c",
X"08e00508",
X"82053483",
X"c08c08e0",
X"050808ff",
X"83ff0682",
X"800783c0",
X"8c08e005",
X"080c83c0",
X"8c08e805",
X"08810533",
X"810583c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"83c08c08",
X"e8050881",
X"05348183",
X"3983c08c",
X"08fc0508",
X"802e80f7",
X"3883c08c",
X"08ec0508",
X"86053383",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08a22e09",
X"810680d7",
X"3883c08c",
X"08ec0508",
X"88053383",
X"c08c08ec",
X"05088705",
X"33718280",
X"290583c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c52",
X"83c08c08",
X"e4050c83",
X"c08c08f4",
X"050c83c0",
X"8c08e405",
X"0883c08c",
X"08e00508",
X"88052383",
X"c08c08ec",
X"05083383",
X"c08c08f0",
X"05087131",
X"7083ffff",
X"0683c08c",
X"08f0050c",
X"83c08c08",
X"e0050c83",
X"c08c08ec",
X"05080583",
X"c08c08ec",
X"050cf6d0",
X"3983c08c",
X"08f80508",
X"0d83c08c",
X"08f00508",
X"83c08c08",
X"e0050c83",
X"c08c08f8",
X"05080d83",
X"c08c08e0",
X"050883c0",
X"800c8d3d",
X"0d83c08c",
X"0c0483c0",
X"8c080283",
X"c08c0ce6",
X"3d0d83c0",
X"8c088805",
X"08028405",
X"83c08c08",
X"e8050c83",
X"c08c08d4",
X"050c800b",
X"83c8bc34",
X"83c08c08",
X"d4050890",
X"0583c08c",
X"08c0050c",
X"800b83c0",
X"8c08c005",
X"0834800b",
X"83c08c08",
X"c0050881",
X"0534800b",
X"83c08c08",
X"c4050c83",
X"c08c08c4",
X"050880d8",
X"2983c08c",
X"08c00508",
X"0583c08c",
X"08ffb405",
X"0c800b83",
X"c08c08ff",
X"b4050880",
X"d8050c83",
X"c08c08ff",
X"b4050884",
X"0583c08c",
X"08ffb405",
X"0c83c08c",
X"08c40508",
X"83c08c08",
X"ffb40508",
X"34880b83",
X"c08c08ff",
X"b4050881",
X"0534800b",
X"83c08c08",
X"ffb40508",
X"82053483",
X"c08c08ff",
X"b4050808",
X"ffa1ff06",
X"a0800783",
X"c08c08ff",
X"b405080c",
X"83c08c08",
X"c4050881",
X"057081ff",
X"0683c08c",
X"08c4050c",
X"83c08c08",
X"ffb4050c",
X"810b83c0",
X"8c08c405",
X"0827fedb",
X"3883c08c",
X"08ec0570",
X"5483c08c",
X"08c8050c",
X"925283c0",
X"8c08d405",
X"085180cd",
X"993f83c0",
X"800881ff",
X"067083c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"05088dea",
X"3883c08c",
X"08f40551",
X"f18c3f83",
X"c0800883",
X"ffff0683",
X"c08c08f6",
X"055283c0",
X"8c08e405",
X"0cf0f33f",
X"83c08008",
X"83ffff06",
X"83c08c08",
X"fd053383",
X"c08c08ff",
X"b8050883",
X"c08c08c4",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08c40508",
X"83c08c08",
X"ffbc0508",
X"2780fe38",
X"83c08c08",
X"c8050854",
X"83c08c08",
X"c4050853",
X"895283c0",
X"8c08d405",
X"085180cc",
X"9e3f83c0",
X"800881ff",
X"0683c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"0880f238",
X"83c08c08",
X"ee0551ef",
X"f13f83c0",
X"800883ff",
X"ff065383",
X"c08c08c4",
X"05085283",
X"c08c08d4",
X"050851f0",
X"b33f83c0",
X"8c08c405",
X"08810570",
X"81ff0683",
X"c08c08c4",
X"050c83c0",
X"8c08ffb4",
X"050cfef1",
X"3983c08c",
X"08c00508",
X"81053383",
X"c08c08ff",
X"b4050c81",
X"db0b83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb4",
X"0508802e",
X"8be03894",
X"3983c08c",
X"08ffb805",
X"0883c08c",
X"08ffbc05",
X"0c8bcb39",
X"83c08c08",
X"f1053352",
X"83c08c08",
X"d4050851",
X"80cb9c3f",
X"800b83c0",
X"8c08c005",
X"08810533",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"c4050c83",
X"c08c08c4",
X"050883c0",
X"8c08ffb4",
X"05082789",
X"e63883c0",
X"8c08c405",
X"0880d829",
X"7083c08c",
X"08c00508",
X"05708805",
X"70830533",
X"83c08c08",
X"cc050c83",
X"c08c08c8",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08d805",
X"0c83c08c",
X"08cc0508",
X"87a63883",
X"c08c08c8",
X"05082202",
X"84057186",
X"0587fffc",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08dc050c",
X"83c08c08",
X"ffb8050c",
X"0283c08c",
X"08ffb405",
X"08310d89",
X"3d705983",
X"c08c08ff",
X"b8050858",
X"83c08c08",
X"ffbc0508",
X"87053357",
X"83c08c08",
X"ffb4050c",
X"a25583c0",
X"8c08cc05",
X"08548653",
X"81815283",
X"c08c08d4",
X"050851be",
X"933f83c0",
X"800881ff",
X"0683c08c",
X"08d0050c",
X"83c08c08",
X"d0050881",
X"c13883c0",
X"8c08ffbc",
X"05089605",
X"5383c08c",
X"08ffb805",
X"085283c0",
X"8c08ffb4",
X"050851a1",
X"c63f83c0",
X"800881ff",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb405",
X"08802e81",
X"853883c0",
X"8c08ffbc",
X"05089405",
X"83c08c08",
X"ffbc0508",
X"96053370",
X"862a83c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08cc05",
X"0c83c08c",
X"08ffb405",
X"08832e09",
X"810680c6",
X"3883c08c",
X"08ffb405",
X"0883c08c",
X"08c80508",
X"82053483",
X"c8a03370",
X"810583c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb4",
X"050883c8",
X"a03483c0",
X"8c08ffb8",
X"050883c0",
X"8c08cc05",
X"083483c0",
X"8c08dc05",
X"080d83c0",
X"8c08d005",
X"0881ff06",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"fbff3883",
X"c08c08d8",
X"050883c0",
X"8c08c005",
X"08058805",
X"70820533",
X"5183c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb405",
X"08832e09",
X"810680e3",
X"3883c08c",
X"08ffb805",
X"0883c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb405",
X"08810570",
X"81ff0651",
X"83c08c08",
X"ffb4050c",
X"810b83c0",
X"8c08ffb4",
X"050827dd",
X"38800b83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b4050881",
X"057081ff",
X"065183c0",
X"8c08ffb4",
X"050c970b",
X"83c08c08",
X"ffb40508",
X"27dd3883",
X"c08c08e4",
X"050880f9",
X"32703070",
X"80255151",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"e0050891",
X"2e098106",
X"80f93883",
X"c08c08ff",
X"b4050880",
X"2e80ec38",
X"83c08c08",
X"c4050880",
X"e238850b",
X"83c08c08",
X"c00508a6",
X"0534a00b",
X"83c08c08",
X"c00508a7",
X"0534850b",
X"83c08c08",
X"c00508a8",
X"053480c0",
X"0b83c08c",
X"08c00508",
X"a9053486",
X"0b83c08c",
X"08c00508",
X"aa053490",
X"0b83c08c",
X"08c00508",
X"ab053486",
X"0b83c08c",
X"08c00508",
X"ac0534a0",
X"0b83c08c",
X"08c00508",
X"ad053483",
X"c08c08e4",
X"050889d8",
X"32703070",
X"80255151",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"e0050883",
X"edec2e09",
X"810680f6",
X"38817083",
X"c08c08ff",
X"b4050806",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb40508",
X"802e80ce",
X"3883c08c",
X"08c40508",
X"80c43884",
X"0b83c08c",
X"08c00508",
X"aa053480",
X"c00b83c0",
X"8c08c005",
X"08ab0534",
X"840b83c0",
X"8c08c005",
X"08ac0534",
X"900b83c0",
X"8c08c005",
X"08ad0534",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"c005088c",
X"053483c0",
X"8c08e405",
X"0880f932",
X"70307080",
X"25515183",
X"c08c08ff",
X"b4050c83",
X"c08c08e0",
X"0508862e",
X"09810680",
X"c3388170",
X"83c08c08",
X"ffb40508",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb405",
X"08802e9c",
X"3883c08c",
X"08c40508",
X"933883c0",
X"8c08ffb8",
X"050883c0",
X"8c08c005",
X"088d0534",
X"83c08c08",
X"c4050880",
X"d82983c0",
X"8c08c005",
X"08057084",
X"05708305",
X"3383c08c",
X"08ffb405",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"ffbc050c",
X"80588057",
X"83c08c08",
X"ffb40508",
X"56805580",
X"548a53a1",
X"5283c08c",
X"08d40508",
X"51b78d3f",
X"83c08008",
X"81ff0670",
X"30709f2a",
X"5183c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"08a02e8c",
X"3883c08c",
X"08ffb405",
X"08f6c238",
X"83c08c08",
X"ffbc0508",
X"8b053383",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b4050880",
X"2eb33883",
X"c08c08c8",
X"05088305",
X"3383c08c",
X"08ffb405",
X"0c805880",
X"5783c08c",
X"08ffb405",
X"08568055",
X"80548b53",
X"a15283c0",
X"8c08d405",
X"0851b688",
X"3f83c08c",
X"08c40508",
X"81057081",
X"ff0683c0",
X"8c08c005",
X"08810533",
X"5283c08c",
X"08c4050c",
X"83c08c08",
X"ffb4050c",
X"f6893980",
X"0b83c08c",
X"08c4050c",
X"83c08c08",
X"c4050880",
X"d82983c0",
X"8c08d405",
X"0805709a",
X"053383c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb4",
X"0508822e",
X"098106a9",
X"3883c8bc",
X"56815580",
X"5483c08c",
X"08ffb405",
X"085383c0",
X"8c08ffb8",
X"05089705",
X"335283c0",
X"8c08d405",
X"0851e48a",
X"3f83c08c",
X"08c40508",
X"81057081",
X"ff0683c0",
X"8c08c405",
X"0c83c08c",
X"08ffb405",
X"0c810b83",
X"c08c08c4",
X"050827fe",
X"fb38810b",
X"83c08c08",
X"c0050834",
X"800b83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08e805",
X"080d83c0",
X"8c08ffbc",
X"050883c0",
X"800c9c3d",
X"0d83c08c",
X"0c04f53d",
X"0d901e57",
X"800b8118",
X"33545978",
X"7327819d",
X"387880d8",
X"29178a11",
X"33545472",
X"832e0981",
X"0680f838",
X"9414335b",
X"a98c3f83",
X"c080085a",
X"80567581",
X"c4291a87",
X"11335454",
X"72802e80",
X"c0387308",
X"81cc982e",
X"098106b5",
X"38807459",
X"557480d8",
X"29189a11",
X"33545472",
X"832e0981",
X"069238a4",
X"14703354",
X"547a7327",
X"8738ff13",
X"53727434",
X"81157081",
X"ff065653",
X"817527d1",
X"38811670",
X"81ff0657",
X"538f7627",
X"ffa43883",
X"c8a033ff",
X"05537283",
X"c8a03481",
X"197081ff",
X"06811933",
X"5e5a537b",
X"7926fee5",
X"38800b83",
X"c0800c8d",
X"3d0d0483",
X"c08c0802",
X"83c08c0c",
X"e63d0d83",
X"c08c0888",
X"05080284",
X"05719005",
X"70337083",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08c8",
X"050c83c0",
X"8c08dc05",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"ffa40508",
X"802e94b5",
X"38800b83",
X"c08c08c8",
X"05088105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08d4050c",
X"83c08c08",
X"d4050883",
X"c08c08ff",
X"a4050825",
X"93fd3883",
X"c08c08d4",
X"050880d8",
X"2983c08c",
X"08c80508",
X"05840570",
X"86053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"a4050880",
X"2e938938",
X"a6b23f83",
X"c08c08ff",
X"b8050880",
X"d4050883",
X"c0800826",
X"92f23802",
X"83c08c08",
X"ffb80508",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08d8",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08fc05",
X"2383c08c",
X"08ffa405",
X"08860583",
X"fc0683c0",
X"8c08ffa4",
X"050c0283",
X"c08c08ff",
X"a4050831",
X"0d853d70",
X"5583c08c",
X"08fc0554",
X"83c08c08",
X"ffb80508",
X"5383c08c",
X"08e00508",
X"5283c08c",
X"08c0050c",
X"ae8a3f83",
X"c0800881",
X"ff0683c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"050891bb",
X"3883c08c",
X"08ffb805",
X"08870533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e80d5",
X"3883c08c",
X"08ffb805",
X"08860533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"822e0981",
X"06b33883",
X"c08c08fc",
X"052283c0",
X"8c08ffa4",
X"050c870b",
X"83c08c08",
X"ffa40508",
X"27973883",
X"c08c08c0",
X"05088205",
X"5283c08c",
X"08c00508",
X"3351dba6",
X"3f83c08c",
X"08ffb805",
X"08860533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"832e0981",
X"0690a438",
X"83c08c08",
X"ffb80508",
X"92057082",
X"053383c0",
X"8c08fc05",
X"2283c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08c4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffa80508",
X"268fe438",
X"800b83c0",
X"8c08e405",
X"0c800b83",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"b0050810",
X"83c08c08",
X"05f80583",
X"c08c08ff",
X"b0050884",
X"2983c08c",
X"08ffb005",
X"08100583",
X"c08c08c4",
X"05080570",
X"84057033",
X"83c08c08",
X"c0050805",
X"703383c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffbc",
X"05082383",
X"c08c08ff",
X"a8050881",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508902e",
X"098106be",
X"3883c08c",
X"08ffa805",
X"083383c0",
X"8c08c005",
X"08058105",
X"70337082",
X"802983c0",
X"8c08ffb4",
X"05080551",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffbc05",
X"082383c0",
X"8c08ffac",
X"05088605",
X"2283c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa805",
X"08a23883",
X"c08c08ff",
X"ac050888",
X"052283c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"050881ff",
X"2e80e538",
X"83c08c08",
X"ffbc0508",
X"227083c0",
X"8c08ffa8",
X"05083170",
X"82802971",
X"3183c08c",
X"08ffac05",
X"08880522",
X"7083c08c",
X"08ffa805",
X"08317073",
X"355383c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c5183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"bc050823",
X"83c08c08",
X"ffb00508",
X"81057081",
X"ff0683c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa4",
X"050c810b",
X"83c08c08",
X"ffb00508",
X"27fce038",
X"83c08c08",
X"f8052283",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a40508bf",
X"26913883",
X"c08c08e4",
X"05088207",
X"83c08c08",
X"e4050c81",
X"c00b83c0",
X"8c08ffa4",
X"05082791",
X"3883c08c",
X"08e40508",
X"810783c0",
X"8c08e405",
X"0c83c08c",
X"08fa0522",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"bf269138",
X"83c08c08",
X"e4050888",
X"0783c08c",
X"08e4050c",
X"81c00b83",
X"c08c08ff",
X"a4050827",
X"913883c0",
X"8c08e405",
X"08840783",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffb00508",
X"1083c08c",
X"08c40508",
X"05709005",
X"703383c0",
X"8c08c005",
X"08057033",
X"72810533",
X"70720651",
X"535183c0",
X"8c08ffa8",
X"050c5183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e9b3890",
X"0b83c08c",
X"08ffb005",
X"082b83c0",
X"8c08e405",
X"080783c0",
X"8c08e405",
X"0c83c08c",
X"08ffb005",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a4050c97",
X"0b83c08c",
X"08ffb005",
X"0827fef4",
X"3883c08c",
X"08ffb805",
X"08900533",
X"83c08c08",
X"e4050883",
X"c08c08ff",
X"b4050c83",
X"c08c08c4",
X"050c83c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffb8",
X"05088c05",
X"082e83ff",
X"3883c08c",
X"08ffb405",
X"0883c08c",
X"08ffb805",
X"088c050c",
X"83c08c08",
X"ffb80508",
X"89053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e83b938",
X"83c08c08",
X"e40583c0",
X"8c08ffb4",
X"05088f06",
X"83c08c08",
X"e4050c83",
X"c08c08cc",
X"050c800b",
X"83c08c08",
X"f0050c80",
X"0b83c08c",
X"08f40523",
X"800b81ce",
X"943383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffbc",
X"05082e82",
X"d33883c0",
X"8c08f005",
X"81ce940b",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"d0050c83",
X"c08c08ff",
X"ac050833",
X"83c08c08",
X"ffac0508",
X"81053381",
X"722b8172",
X"2b077083",
X"c08c08ff",
X"b4050806",
X"5283c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffa805",
X"082e0981",
X"0681be38",
X"83c08c08",
X"ffbc0508",
X"852680f6",
X"3883c08c",
X"08ffac05",
X"08820533",
X"7081ff06",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa40508",
X"802e80ca",
X"3883c08c",
X"08ffbc05",
X"0883c08c",
X"08ffbc05",
X"08810570",
X"81ff0683",
X"c08c08d0",
X"05087305",
X"5383c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb005",
X"0883c08c",
X"08ffa405",
X"083483c0",
X"8c08ffac",
X"05088305",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e9d",
X"38810b83",
X"c08c08ff",
X"a405082b",
X"83c08c08",
X"cc050808",
X"0783c08c",
X"08cc0508",
X"0c83c08c",
X"08ffac05",
X"08840570",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa405",
X"08fdc838",
X"83c08c08",
X"f0055280",
X"51d0c33f",
X"83c08c08",
X"e4050852",
X"83c08c08",
X"c4050851",
X"d1fe3f83",
X"c08c08fb",
X"05337081",
X"800a2981",
X"0a057098",
X"2c5583c0",
X"8c08ffa4",
X"050c83c0",
X"8c08f905",
X"33708180",
X"0a29810a",
X"0570982c",
X"5583c08c",
X"08ffa405",
X"0c83c08c",
X"08c40508",
X"5383c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa805",
X"0cd1d43f",
X"83c08c08",
X"ffb80508",
X"88053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e84e038",
X"83c08c08",
X"ffb80508",
X"90053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050881",
X"2684c038",
X"807081ce",
X"c80b81ce",
X"c80b8105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffb405",
X"082e81ae",
X"3883c08c",
X"08ffac05",
X"08842983",
X"c08c08ff",
X"a8050805",
X"703383c0",
X"8c08c005",
X"08057033",
X"72810533",
X"70720651",
X"535183c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"aa38810b",
X"83c08c08",
X"ffac0508",
X"2b83c08c",
X"08ffb405",
X"08077083",
X"ffff0683",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"ac050881",
X"057081ff",
X"0681cec8",
X"71842971",
X"05708105",
X"33515383",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a40508fe",
X"d43883c0",
X"8c08ffb8",
X"05088a05",
X"2283c08c",
X"08c0050c",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"c005082e",
X"82ad3880",
X"0b83c08c",
X"08e8050c",
X"800b83c0",
X"8c08ec05",
X"23807083",
X"c08c08e8",
X"0583c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffb005",
X"0c81af39",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffac0508",
X"2c708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e80",
X"e73883c0",
X"8c08ffb0",
X"050883c0",
X"8c08ffb0",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ffbc0508",
X"730583c0",
X"8c08ffb8",
X"05089005",
X"3383c08c",
X"08ffac05",
X"08842905",
X"535383c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050881ce",
X"ca053383",
X"c08c08ff",
X"a4050834",
X"83c08c08",
X"ffac0508",
X"81057081",
X"ff0683c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa4",
X"050c8f0b",
X"83c08c08",
X"ffac0508",
X"2783c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb005",
X"0885268c",
X"3883c08c",
X"08ffa405",
X"08fea938",
X"83c08c08",
X"e8055280",
X"51caf33f",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffb80508",
X"8a052383",
X"c08c08ff",
X"b8050880",
X"d2053383",
X"c08c08ff",
X"b8050880",
X"d4050805",
X"83c08c08",
X"ffb80508",
X"80d4050c",
X"83c08c08",
X"d805080d",
X"83c08c08",
X"d4050881",
X"800a2981",
X"800a0570",
X"982c83c0",
X"8c08c805",
X"08810533",
X"83c08c08",
X"ffa8050c",
X"5183c08c",
X"08d4050c",
X"83c08c08",
X"ffa80508",
X"83c08c08",
X"d4050824",
X"ec853880",
X"0b83c08c",
X"08ffa805",
X"0c83c08c",
X"08dc0508",
X"0d83c08c",
X"08ffa805",
X"0883c080",
X"0c9c3d0d",
X"83c08c0c",
X"04f33d0d",
X"02bf0533",
X"02840580",
X"c3053383",
X"c8bc335a",
X"5b597980",
X"2e8d3878",
X"78065776",
X"802e8e38",
X"81893978",
X"78065776",
X"802e80ff",
X"3883c8bc",
X"33707a07",
X"58587988",
X"38780970",
X"79065157",
X"7683c8bc",
X"3492973f",
X"83c08008",
X"5e805c8f",
X"5d7d1c87",
X"11335858",
X"76802e80",
X"c1387708",
X"81cc982e",
X"098106b6",
X"38805b81",
X"5a7d1c70",
X"1c9a1133",
X"59595976",
X"822e0981",
X"06943883",
X"c8bc5681",
X"55805476",
X"53971833",
X"527851cb",
X"c53fff1a",
X"80d81c5c",
X"5a798025",
X"d038ff1d",
X"81c41d5d",
X"5d7c8025",
X"ffa7388f",
X"3d0d04e9",
X"3d0d696c",
X"02880580",
X"ea05225c",
X"5a5b8070",
X"71415e58",
X"ff78797a",
X"7b7c7d46",
X"4c4a4540",
X"5d436299",
X"3d346202",
X"840580dd",
X"05347779",
X"2280ffff",
X"06544572",
X"79237978",
X"2e888738",
X"7a708105",
X"5c337084",
X"2a718c06",
X"70822a5a",
X"56568306",
X"ff1b7083",
X"ffff065c",
X"54568054",
X"75742e91",
X"387a7081",
X"055c33ff",
X"1b7083ff",
X"ff065c54",
X"54817627",
X"9b387381",
X"ff067b70",
X"81055d33",
X"55748280",
X"2905ff1b",
X"7083ffff",
X"065c5454",
X"827627aa",
X"387383ff",
X"ff067b70",
X"81055d33",
X"70902b72",
X"077d7081",
X"055f3370",
X"982b7207",
X"fe1f7083",
X"ffff0640",
X"52525252",
X"54547e80",
X"2e80c438",
X"7686f738",
X"748a2e09",
X"81069438",
X"811f7081",
X"ff06811e",
X"7081ff06",
X"5f524053",
X"86dc3974",
X"8c2e0981",
X"0686d338",
X"ff1f7081",
X"ff06ff1e",
X"7081ff06",
X"5f524053",
X"7b632586",
X"bd38ff43",
X"86b83976",
X"812e83bb",
X"38768124",
X"89387680",
X"2e8d3886",
X"a5397682",
X"2e84a638",
X"869c39f8",
X"15537284",
X"26849538",
X"72842981",
X"cf880553",
X"72080464",
X"802e80cd",
X"38782283",
X"80800653",
X"72838080",
X"2e098106",
X"bc388056",
X"756427a4",
X"38751e70",
X"83ffff06",
X"77101b90",
X"1172832a",
X"58515751",
X"53737534",
X"72870681",
X"712b5153",
X"72811634",
X"81167081",
X"ff065753",
X"977627cc",
X"387f8407",
X"40800b99",
X"3d435661",
X"16703370",
X"982b7098",
X"2c515151",
X"53807324",
X"80fb3860",
X"73291e70",
X"83ffff06",
X"7a228380",
X"80065258",
X"53728380",
X"802e0981",
X"0680de38",
X"60883270",
X"30707207",
X"80256390",
X"32703070",
X"72078025",
X"73075354",
X"58515553",
X"73802ebd",
X"38768706",
X"5372b638",
X"75842976",
X"10057911",
X"84117983",
X"2a575751",
X"53737534",
X"60811634",
X"65861423",
X"66881423",
X"7587387f",
X"8107408d",
X"3975812e",
X"09810685",
X"387f8207",
X"40811670",
X"81ff0657",
X"53817627",
X"fee53863",
X"61291e70",
X"83ffff06",
X"5f538070",
X"4642ff02",
X"840580dd",
X"0534ff0b",
X"993d3483",
X"f539811c",
X"7081ff06",
X"5d538042",
X"73812e09",
X"81068e38",
X"7781800a",
X"2981800a",
X"055880d3",
X"3973802e",
X"89387382",
X"2e098106",
X"8d387c81",
X"800a2981",
X"800a055d",
X"a439815f",
X"83b839ff",
X"1c7081ff",
X"065d537b",
X"63258338",
X"ff437c80",
X"2e92387c",
X"81800a29",
X"81ff0a05",
X"5d7c982c",
X"5d839339",
X"77802e92",
X"38778180",
X"0a2981ff",
X"0a055877",
X"982c5882",
X"fd397753",
X"839e3974",
X"892680f4",
X"38748429",
X"81cf9c05",
X"53720804",
X"73872e82",
X"e1387385",
X"2e82db38",
X"73882e82",
X"d538738c",
X"2e82cf38",
X"73892e09",
X"81068638",
X"814582c2",
X"3973812e",
X"09810682",
X"b9386280",
X"2582b338",
X"7b982b70",
X"982c5143",
X"82a83973",
X"83ffff06",
X"46829f39",
X"7383ffff",
X"06478296",
X"397381ff",
X"0641828e",
X"3973811a",
X"34828739",
X"7381ff06",
X"4481ff39",
X"7e5382a0",
X"3974812e",
X"81e33874",
X"81248938",
X"74802e8d",
X"3881e739",
X"74822e81",
X"d83881de",
X"3974567b",
X"83388156",
X"74537386",
X"2e098106",
X"97387581",
X"06537280",
X"2e8e3878",
X"2282ffff",
X"06fe8080",
X"0753b639",
X"7b833881",
X"5373822e",
X"09810697",
X"38728106",
X"5372802e",
X"8e387822",
X"81ffff06",
X"81808007",
X"5393397b",
X"9638fc14",
X"53728126",
X"8e387822",
X"ff808007",
X"53727923",
X"80e53980",
X"5573812e",
X"09810683",
X"38735577",
X"5377802e",
X"89387481",
X"06537280",
X"ca3872d0",
X"15545572",
X"81268338",
X"81557780",
X"2eb93874",
X"81065372",
X"802eb038",
X"78228380",
X"80065372",
X"8380802e",
X"0981069f",
X"3873b02e",
X"09810687",
X"3861993d",
X"34913973",
X"b12e0981",
X"06893861",
X"02840580",
X"dd053461",
X"8105538c",
X"39617431",
X"81055384",
X"39611453",
X"7283ffff",
X"064279f7",
X"fb387d83",
X"2a537282",
X"1a347822",
X"83808006",
X"53728380",
X"802e0981",
X"06883881",
X"537f872e",
X"83388053",
X"7283c080",
X"0c993d0d",
X"04fd3d0d",
X"75831133",
X"82123371",
X"982b7190",
X"2b078114",
X"3370882b",
X"72077533",
X"710783c0",
X"800c5253",
X"54565452",
X"853d0d04",
X"f63d0d02",
X"b7053302",
X"8405bb05",
X"33028805",
X"bf05335b",
X"5b5b8058",
X"80577888",
X"2b7a0756",
X"80557a54",
X"8153a352",
X"7c5192cc",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8c3d0d04",
X"f63d0d02",
X"b7053302",
X"8405bb05",
X"33028805",
X"bf05335b",
X"5b5b8058",
X"80577888",
X"2b7a0756",
X"80557a54",
X"8353a352",
X"7c519290",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8c3d0d04",
X"f73d0d02",
X"b3053302",
X"8405b605",
X"22605a58",
X"56805580",
X"54805381",
X"a3527b51",
X"91e23f83",
X"c0800881",
X"ff0683c0",
X"800c8b3d",
X"0d04ee3d",
X"0d649011",
X"5c5c807b",
X"34800b84",
X"1c0c800b",
X"881c3481",
X"0b891c34",
X"880b8a1c",
X"34800b8b",
X"1c34881b",
X"08c10681",
X"07881c0c",
X"8f3d7054",
X"5d88527b",
X"519beb3f",
X"83c08008",
X"81ff0670",
X"5b597881",
X"a938903d",
X"335e81db",
X"5a7d892e",
X"09810681",
X"99387c53",
X"92527b51",
X"9bc43f83",
X"c0800881",
X"ff06705b",
X"59788182",
X"387c5888",
X"577856a9",
X"55785486",
X"5381a052",
X"7b5190d0",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"80e03802",
X"ba05337b",
X"347c5478",
X"537d527b",
X"519bac3f",
X"83c08008",
X"81ff0670",
X"5b597880",
X"c13802bd",
X"0533527b",
X"519bc43f",
X"83c08008",
X"81ff0670",
X"5b5978aa",
X"38817b33",
X"5a5a7979",
X"26993880",
X"54795388",
X"527b51fd",
X"bb3f811a",
X"7081ff06",
X"7c33525b",
X"59e43981",
X"0b881c34",
X"805a7983",
X"c0800c94",
X"3d0d0480",
X"0b83c080",
X"0c04f93d",
X"0d790284",
X"05ab0533",
X"8e3d7054",
X"585858ff",
X"beb03f8a",
X"3d8a0551",
X"ffbea73f",
X"7551fc8d",
X"3f83c080",
X"08848681",
X"2ebe3883",
X"c0800884",
X"86812699",
X"3883c080",
X"08848280",
X"2e80e638",
X"83c08008",
X"8482812e",
X"9f3881b4",
X"3983c080",
X"0880c082",
X"832e80f4",
X"3883c080",
X"0880c086",
X"832e80e8",
X"38819939",
X"83c09c33",
X"55805674",
X"762e0981",
X"06818b38",
X"74547653",
X"91527751",
X"fbd63f74",
X"54765390",
X"527751fb",
X"cb3f7454",
X"76538452",
X"7751fbfc",
X"3f810b83",
X"c09c3481",
X"b15680de",
X"39805476",
X"53915277",
X"51fba93f",
X"80547653",
X"90527751",
X"fb9e3f80",
X"0b83c09c",
X"34765287",
X"18335197",
X"963fb539",
X"80547653",
X"94527751",
X"fb823f80",
X"54765390",
X"527751fa",
X"f73f7551",
X"ffbcdb3f",
X"83c08008",
X"892a8106",
X"53765287",
X"18335190",
X"cd3f800b",
X"83c09c34",
X"80567583",
X"c0800c89",
X"3d0d04f2",
X"3d0d6090",
X"115a5880",
X"0b881a33",
X"71595656",
X"74762e82",
X"a53882ac",
X"3f841908",
X"83c08008",
X"26829538",
X"78335a81",
X"0b8e3d23",
X"903df811",
X"55f40553",
X"99185277",
X"518ae53f",
X"83c08008",
X"81ff0670",
X"57557477",
X"2e098106",
X"81d93886",
X"39745681",
X"d2398156",
X"82578e3d",
X"33770655",
X"74802ebb",
X"38800b8d",
X"3d34903d",
X"f0055484",
X"53755277",
X"51facd3f",
X"83c08008",
X"81ff0655",
X"749d387b",
X"53755277",
X"51fce73f",
X"83c08008",
X"81ff0655",
X"7481b12e",
X"818b3874",
X"ffb33876",
X"1081fc06",
X"81177081",
X"ff065856",
X"57877627",
X"ffa83881",
X"56757a26",
X"80eb3880",
X"0b8d3d34",
X"8c3d7055",
X"57845375",
X"527751f9",
X"f73f83c0",
X"800881ff",
X"06557480",
X"c1387651",
X"ffbad73f",
X"83c08008",
X"82870655",
X"7482812e",
X"098106aa",
X"3802ae05",
X"33810755",
X"74028405",
X"ae05347b",
X"53755277",
X"51fbeb3f",
X"83c08008",
X"81ff0655",
X"7481b12e",
X"903874fe",
X"b8388116",
X"7081ff06",
X"5755ff91",
X"39805675",
X"81ff0656",
X"973f83c0",
X"80088fd0",
X"05841a0c",
X"75577683",
X"c0800c90",
X"3d0d0404",
X"9080a008",
X"83c0800c",
X"04ff3d0d",
X"7387e829",
X"51ffa2f9",
X"3f833d0d",
X"040483c8",
X"c00b83c0",
X"800c04fd",
X"3d0d7577",
X"5454800b",
X"83c8a034",
X"728a3890",
X"90800b84",
X"150c9039",
X"72812e09",
X"81068838",
X"9098800b",
X"84150c84",
X"140883c8",
X"b80c800b",
X"88150c80",
X"0b8c150c",
X"83c8b808",
X"53820b87",
X"80143481",
X"51ff9e3f",
X"83c8b808",
X"53800b88",
X"143483c8",
X"b8085381",
X"0b878014",
X"3483c8b8",
X"0853800b",
X"8c143483",
X"c8b80853",
X"800ba414",
X"34917434",
X"800b83c0",
X"a034800b",
X"83c0a434",
X"800b83c0",
X"a8348054",
X"7381c429",
X"83c8c405",
X"53800b83",
X"14348114",
X"7081ff06",
X"55538f74",
X"27e63885",
X"3d0d04fe",
X"3d0d7476",
X"82113370",
X"bf068171",
X"2bff0556",
X"51515253",
X"90712783",
X"38ff5276",
X"51717123",
X"83c8b808",
X"51871333",
X"90123480",
X"0b83c0a4",
X"34800b83",
X"c0a83488",
X"13338a14",
X"33525271",
X"802eaa38",
X"7081ff06",
X"51845270",
X"83387052",
X"7183c0a4",
X"348a1333",
X"70307080",
X"25842b70",
X"88075151",
X"52537083",
X"c0a83490",
X"397081ff",
X"06517083",
X"38985271",
X"83c0a834",
X"800b83c0",
X"800c843d",
X"0d04f13d",
X"0d616568",
X"028c0580",
X"cb053302",
X"900580ce",
X"05220294",
X"0580d605",
X"22424041",
X"5a4040fd",
X"8b3f83c0",
X"8008a788",
X"055b8070",
X"715b5b52",
X"83943983",
X"c8b80851",
X"7d941234",
X"83c0a433",
X"81075580",
X"7054567f",
X"862680ea",
X"387f8429",
X"81cfd005",
X"83c8b808",
X"53517008",
X"04800b84",
X"1334a139",
X"77337030",
X"70802583",
X"71315151",
X"52537084",
X"13348d39",
X"810b8413",
X"34b83983",
X"0b841334",
X"81705456",
X"ad39810b",
X"841334a2",
X"39773370",
X"30708025",
X"83713151",
X"51525370",
X"84133480",
X"78335252",
X"70833881",
X"52717834",
X"81537488",
X"075583c0",
X"a83383c8",
X"b8085257",
X"810b81d0",
X"123483c8",
X"b8085181",
X"0b819012",
X"347e802e",
X"ae387280",
X"2ea9387e",
X"ff1e5254",
X"7083ffff",
X"06537283",
X"ffff2e97",
X"38737081",
X"05553383",
X"c8b80853",
X"517081c0",
X"1334ff13",
X"51de3983",
X"c8b808a8",
X"11335351",
X"76881234",
X"83c8b808",
X"51747134",
X"81ff5291",
X"3983c8b8",
X"08a01133",
X"70810651",
X"5253708f",
X"38fafd3f",
X"7a83c080",
X"0826e638",
X"81883981",
X"0ba01434",
X"83c8b808",
X"a8113380",
X"ff067078",
X"07525351",
X"70802e80",
X"ed387186",
X"2a708106",
X"51517080",
X"2e913880",
X"78335253",
X"70833881",
X"53727834",
X"80e03971",
X"842a7081",
X"06515170",
X"802e9b38",
X"81197083",
X"ffff067d",
X"30709f2a",
X"51525a51",
X"787c2e09",
X"8106af38",
X"a4397183",
X"2a708106",
X"51517080",
X"2e933881",
X"1a7081ff",
X"065b5179",
X"832e0981",
X"0690388a",
X"3971a306",
X"5170802e",
X"85387151",
X"9239f9e4",
X"3f7a83c0",
X"800826fc",
X"e2387181",
X"bf065170",
X"83c0800c",
X"913d0d04",
X"f63d0d02",
X"b3053302",
X"8405b705",
X"33028805",
X"ba052259",
X"5959800b",
X"8c3d348c",
X"3dfc0556",
X"80558054",
X"76537752",
X"7851fbf2",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8c3d0d04",
X"f33d0d7f",
X"6264028c",
X"0580c205",
X"22722281",
X"1533425f",
X"415e5959",
X"8078237d",
X"53783352",
X"8151ffa0",
X"3f83c080",
X"0881ff06",
X"5675802e",
X"86387554",
X"81ad3983",
X"c8b808a8",
X"1133821b",
X"3370862a",
X"70810673",
X"982b5351",
X"575c5657",
X"79802583",
X"38815673",
X"762e8738",
X"81f05481",
X"8239818c",
X"17337081",
X"ff067922",
X"7d713190",
X"2b70902c",
X"7009709f",
X"2c720670",
X"52525351",
X"53575754",
X"75742483",
X"38755574",
X"84808029",
X"fc808005",
X"70902c51",
X"5574ff2e",
X"943883c8",
X"b8088180",
X"11335154",
X"737c7081",
X"055e34db",
X"39772276",
X"05547378",
X"23790970",
X"9f2a7081",
X"06821c33",
X"81bf0671",
X"862b0751",
X"51515473",
X"821a347c",
X"76268a38",
X"7722547a",
X"7426febb",
X"38805473",
X"83c0800c",
X"8f3d0d04",
X"f93d0d7a",
X"57800b89",
X"3d23893d",
X"fc055376",
X"527951f8",
X"da3f83c0",
X"800881ff",
X"06705755",
X"7496387c",
X"547b5388",
X"3d225276",
X"51fde53f",
X"83c08008",
X"81ff0656",
X"7583c080",
X"0c893d0d",
X"04f03d0d",
X"62660288",
X"0580ce05",
X"22415d5e",
X"80028405",
X"80d20522",
X"7f810533",
X"ff115a5d",
X"5a5d81da",
X"5876bf26",
X"80e93878",
X"802e80e1",
X"387a5878",
X"7b278338",
X"7858821e",
X"3370872a",
X"585a7692",
X"3d34923d",
X"fc055677",
X"557b547e",
X"537d3352",
X"8251f8de",
X"3f83c080",
X"0881ff06",
X"5d800b92",
X"3d33585a",
X"76802e83",
X"38815a82",
X"1e3380ff",
X"067a872b",
X"07577682",
X"1f347c91",
X"38787831",
X"7083ffff",
X"06791e5e",
X"5a57ff9b",
X"397c5877",
X"83c0800c",
X"923d0d04",
X"f83d0d7b",
X"028405b2",
X"05225858",
X"800b8a3d",
X"238a3dfc",
X"05537752",
X"7a51f6f7",
X"3f83c080",
X"0881ff06",
X"70575574",
X"96387d54",
X"7653893d",
X"22527751",
X"feaf3f83",
X"c0800881",
X"ff065675",
X"83c0800c",
X"8a3d0d04",
X"ec3d0d66",
X"6e028805",
X"80df0533",
X"028c0580",
X"e3053302",
X"900580e7",
X"05330294",
X"0580eb05",
X"33029805",
X"80ee0522",
X"4143415f",
X"5c405702",
X"80f20522",
X"963d2396",
X"3df00553",
X"84177053",
X"775259f6",
X"863f83c0",
X"800881ff",
X"06587781",
X"e538777a",
X"81800658",
X"40807725",
X"83388140",
X"79943d34",
X"7b028405",
X"80c90534",
X"7c028405",
X"80ca0534",
X"7d028405",
X"80cb0534",
X"7a953d34",
X"7a882a57",
X"76028405",
X"80cd0534",
X"953d2257",
X"76028405",
X"80ce0534",
X"76882a57",
X"76028405",
X"80cf0534",
X"77923d34",
X"963dec11",
X"57578855",
X"f4175492",
X"3d225377",
X"527751f6",
X"953f83c0",
X"800881ff",
X"06587780",
X"ed387e80",
X"2e80cb38",
X"923d2279",
X"0858587f",
X"802e9c38",
X"76818080",
X"07790c7e",
X"54963dfc",
X"05537783",
X"ffff0652",
X"7851f9fc",
X"3f993976",
X"82808007",
X"790c7e54",
X"953d2253",
X"7783ffff",
X"06527851",
X"fc8f3f83",
X"c0800881",
X"ff065877",
X"9d38923d",
X"22538052",
X"7f307080",
X"25847131",
X"535157f9",
X"873f83c0",
X"800881ff",
X"06587783",
X"c0800c96",
X"3d0d04f6",
X"3d0d7c02",
X"8405b705",
X"335b5b80",
X"58805780",
X"56805579",
X"54855380",
X"527a51fd",
X"a33f83c0",
X"800881ff",
X"06597885",
X"3879871c",
X"347883c0",
X"800c8c3d",
X"0d04f93d",
X"0d02a705",
X"33028405",
X"ab053302",
X"8805af05",
X"33585957",
X"800b83c8",
X"c7335454",
X"72742e9f",
X"38811470",
X"81ff0655",
X"53738f26",
X"81b63873",
X"81c42983",
X"c8c40583",
X"11335153",
X"72e33873",
X"81c42983",
X"c8c00555",
X"800b8716",
X"34768816",
X"34758a16",
X"34778916",
X"3480750c",
X"83c8b808",
X"8c160c80",
X"0b841634",
X"880b8516",
X"34800b86",
X"16348415",
X"08ffa1ff",
X"06a08007",
X"84160c81",
X"147081ff",
X"06535374",
X"51febc3f",
X"83c08008",
X"81ff0670",
X"55537280",
X"cd388a39",
X"7308750c",
X"725480c2",
X"397281d2",
X"e0555681",
X"d2e00880",
X"2eb23875",
X"84291470",
X"08765370",
X"08515454",
X"722d83c0",
X"800881ff",
X"06537280",
X"2ece3881",
X"167081ff",
X"0681d2e0",
X"71842911",
X"53565753",
X"7208d038",
X"80547383",
X"c0800c89",
X"3d0d04f9",
X"3d0d7957",
X"800b8418",
X"0883c8b8",
X"0c58f088",
X"3f881708",
X"83c08008",
X"2783ed38",
X"effa3f83",
X"c0800881",
X"0588180c",
X"83c8b808",
X"b8113370",
X"81ff0651",
X"51547381",
X"2ea43873",
X"81248838",
X"73782e8a",
X"38b83973",
X"822e9538",
X"b1397633",
X"81f00654",
X"73902ea6",
X"38917734",
X"a1397358",
X"763381f0",
X"06547390",
X"2e098106",
X"9138efa8",
X"3f83c080",
X"0881c805",
X"8c180ca0",
X"77348056",
X"7581c429",
X"83c8c711",
X"33555573",
X"802eaa38",
X"83c8c015",
X"70085654",
X"74802e9d",
X"38881508",
X"802e9638",
X"8c140883",
X"c8b8082e",
X"09810689",
X"38735188",
X"15085473",
X"2d811670",
X"81ff0657",
X"548f7627",
X"ffba3876",
X"335473b0",
X"2e819938",
X"73b0248f",
X"3873912e",
X"ab3873a0",
X"2e80f538",
X"82a63973",
X"80d02e81",
X"e4387380",
X"d0248b38",
X"7380c02e",
X"81993882",
X"8f397381",
X"802e81fb",
X"38828539",
X"80567581",
X"c42983c8",
X"c4118311",
X"33565955",
X"73802ea8",
X"3883c8c0",
X"15700856",
X"5474802e",
X"9b388c14",
X"0883c8b8",
X"082e0981",
X"068e3873",
X"51841508",
X"54732d80",
X"0b831934",
X"81167081",
X"ff065754",
X"8f7627ff",
X"b9389277",
X"3481b539",
X"edc23f8c",
X"170883c0",
X"80082781",
X"a738b077",
X"3481a139",
X"83c8b808",
X"54800b8c",
X"153483c8",
X"b8085484",
X"0b881534",
X"80c07734",
X"ed963f83",
X"c08008b2",
X"058c180c",
X"80fa39ed",
X"873f8c17",
X"0883c080",
X"082780ec",
X"3883c8b8",
X"0854810b",
X"8c153483",
X"c8b80854",
X"800b8815",
X"3483c8b8",
X"0854880b",
X"a01534ec",
X"db3f83c0",
X"80089405",
X"8c180c80",
X"d07734bc",
X"3983c8b8",
X"08a01133",
X"70832a70",
X"81065151",
X"55557380",
X"2ea63888",
X"0ba01634",
X"ecae3f8c",
X"170883c0",
X"80082794",
X"38ff8077",
X"348e3977",
X"53805280",
X"51fa8b3f",
X"ff907734",
X"83c8b808",
X"a0113370",
X"832a7081",
X"06515155",
X"5573802e",
X"8638880b",
X"a0163489",
X"3d0d04f6",
X"3d0d02b3",
X"05330284",
X"05b70533",
X"5b5b800b",
X"83c8c470",
X"84127274",
X"5d59575b",
X"58568315",
X"33537280",
X"2e80f338",
X"7333537a",
X"732e0981",
X"0680e738",
X"81143353",
X"79732e09",
X"810680da",
X"38805574",
X"81c42983",
X"c8c80570",
X"33831b33",
X"58555373",
X"762e0981",
X"068a3881",
X"13335273",
X"51ff9c3f",
X"81157081",
X"ff065653",
X"8f7527d3",
X"38800b83",
X"c8c01970",
X"08565455",
X"73752e91",
X"38725184",
X"14085372",
X"2d83c080",
X"0881ff06",
X"55800b83",
X"18347453",
X"a0398116",
X"81c41981",
X"c41781c4",
X"1781c41d",
X"81c41c5c",
X"5d575759",
X"568f7625",
X"fee83880",
X"537283c0",
X"800c8c3d",
X"0d04f83d",
X"0d02ae05",
X"227d5957",
X"80568155",
X"80548653",
X"8180527a",
X"51f5953f",
X"83c08008",
X"81ff0683",
X"c0800c8a",
X"3d0d04f7",
X"3d0d02b2",
X"05220284",
X"05b70533",
X"605a5b57",
X"80568255",
X"79548653",
X"8180527b",
X"51f4e53f",
X"83c08008",
X"81ff0683",
X"c0800c8b",
X"3d0d04f8",
X"3d0d02af",
X"05335980",
X"58805780",
X"56805578",
X"54895380",
X"527a51f4",
X"bb3f83c0",
X"800881ff",
X"0683c080",
X"0c8a3d0d",
X"0483c08c",
X"080283c0",
X"8c0cfd3d",
X"0d805383",
X"c08c088c",
X"05085283",
X"c08c0888",
X"05085183",
X"d43f83c0",
X"80087083",
X"c0800c54",
X"853d0d83",
X"c08c0c04",
X"83c08c08",
X"0283c08c",
X"0cfd3d0d",
X"815383c0",
X"8c088c05",
X"085283c0",
X"8c088805",
X"085183a1",
X"3f83c080",
X"087083c0",
X"800c5485",
X"3d0d83c0",
X"8c0c0483",
X"c08c0802",
X"83c08c0c",
X"f93d0d80",
X"0b83c08c",
X"08fc050c",
X"83c08c08",
X"88050880",
X"25b93883",
X"c08c0888",
X"05083083",
X"c08c0888",
X"050c800b",
X"83c08c08",
X"f4050c83",
X"c08c08fc",
X"05088a38",
X"810b83c0",
X"8c08f405",
X"0c83c08c",
X"08f40508",
X"83c08c08",
X"fc050c83",
X"c08c088c",
X"05088025",
X"b93883c0",
X"8c088c05",
X"083083c0",
X"8c088c05",
X"0c800b83",
X"c08c08f0",
X"050c83c0",
X"8c08fc05",
X"088a3881",
X"0b83c08c",
X"08f0050c",
X"83c08c08",
X"f0050883",
X"c08c08fc",
X"050c8053",
X"83c08c08",
X"8c050852",
X"83c08c08",
X"88050851",
X"81df3f83",
X"c0800870",
X"83c08c08",
X"f8050c54",
X"83c08c08",
X"fc050880",
X"2e903883",
X"c08c08f8",
X"05083083",
X"c08c08f8",
X"050c83c0",
X"8c08f805",
X"087083c0",
X"800c5489",
X"3d0d83c0",
X"8c0c0483",
X"c08c0802",
X"83c08c0c",
X"fb3d0d80",
X"0b83c08c",
X"08fc050c",
X"83c08c08",
X"88050880",
X"25993883",
X"c08c0888",
X"05083083",
X"c08c0888",
X"050c810b",
X"83c08c08",
X"fc050c83",
X"c08c088c",
X"05088025",
X"903883c0",
X"8c088c05",
X"083083c0",
X"8c088c05",
X"0c815383",
X"c08c088c",
X"05085283",
X"c08c0888",
X"050851bd",
X"3f83c080",
X"087083c0",
X"8c08f805",
X"0c5483c0",
X"8c08fc05",
X"08802e90",
X"3883c08c",
X"08f80508",
X"3083c08c",
X"08f8050c",
X"83c08c08",
X"f8050870",
X"83c0800c",
X"54873d0d",
X"83c08c0c",
X"0483c08c",
X"080283c0",
X"8c0cfd3d",
X"0d810b83",
X"c08c08fc",
X"050c800b",
X"83c08c08",
X"f8050c83",
X"c08c088c",
X"050883c0",
X"8c088805",
X"0827b938",
X"83c08c08",
X"fc050880",
X"2eae3880",
X"0b83c08c",
X"088c0508",
X"24a23883",
X"c08c088c",
X"05081083",
X"c08c088c",
X"050c83c0",
X"8c08fc05",
X"081083c0",
X"8c08fc05",
X"0cffb839",
X"83c08c08",
X"fc050880",
X"2e80e138",
X"83c08c08",
X"8c050883",
X"c08c0888",
X"050826ad",
X"3883c08c",
X"08880508",
X"83c08c08",
X"8c050831",
X"83c08c08",
X"88050c83",
X"c08c08f8",
X"050883c0",
X"8c08fc05",
X"080783c0",
X"8c08f805",
X"0c83c08c",
X"08fc0508",
X"812a83c0",
X"8c08fc05",
X"0c83c08c",
X"088c0508",
X"812a83c0",
X"8c088c05",
X"0cff9539",
X"83c08c08",
X"90050880",
X"2e933883",
X"c08c0888",
X"05087083",
X"c08c08f4",
X"050c5191",
X"3983c08c",
X"08f80508",
X"7083c08c",
X"08f4050c",
X"5183c08c",
X"08f40508",
X"83c0800c",
X"853d0d83",
X"c08c0c04",
X"83c08c08",
X"0283c08c",
X"0cff3d0d",
X"800b83c0",
X"8c08fc05",
X"0c83c08c",
X"08880508",
X"8106ff11",
X"70097083",
X"c08c088c",
X"05080683",
X"c08c08fc",
X"05081183",
X"c08c08fc",
X"050c83c0",
X"8c088805",
X"08812a83",
X"c08c0888",
X"050c83c0",
X"8c088c05",
X"081083c0",
X"8c088c05",
X"0c515151",
X"5183c08c",
X"08880508",
X"802e8438",
X"ffab3983",
X"c08c08fc",
X"05087083",
X"c0800c51",
X"833d0d83",
X"c08c0c04",
X"fc3d0d76",
X"70797b55",
X"5555558f",
X"72278c38",
X"72750783",
X"06517080",
X"2ea938ff",
X"125271ff",
X"2e983872",
X"70810554",
X"33747081",
X"055634ff",
X"125271ff",
X"2e098106",
X"ea387483",
X"c0800c86",
X"3d0d0474",
X"51727084",
X"05540871",
X"70840553",
X"0c727084",
X"05540871",
X"70840553",
X"0c727084",
X"05540871",
X"70840553",
X"0c727084",
X"05540871",
X"70840553",
X"0cf01252",
X"718f26c9",
X"38837227",
X"95387270",
X"84055408",
X"71708405",
X"530cfc12",
X"52718326",
X"ed387054",
X"ff813900",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00002d8e",
X"00002dcf",
X"00002def",
X"00002e14",
X"00002e20",
X"000038f6",
X"0000413a",
X"000041f3",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3a00",
X"0c0c3b00",
X"0a0a0008",
X"0b0b0008",
X"07070008",
X"0a0b4300",
X"080b4200",
X"04044500",
X"05054400",
X"06060004",
X"08080004",
X"09090004",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"00004e7f",
X"00005186",
X"00004f92",
X"00005186",
X"00004fcf",
X"00005020",
X"0000505f",
X"00005068",
X"00005186",
X"00005186",
X"00005186",
X"00005186",
X"00005071",
X"00005079",
X"00005080",
X"00005286",
X"0000537f",
X"00005493",
X"00005789",
X"000057a4",
X"00005790",
X"000057a4",
X"000057ab",
X"000057b6",
X"000057bd",
X"25732025",
X"73000000",
X"20000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"31364b00",
X"556e6b6e",
X"6f776e20",
X"74797065",
X"206f6620",
X"63617274",
X"72696467",
X"65210000",
X"41353200",
X"43415200",
X"42494e00",
X"31366b20",
X"63617274",
X"20747970",
X"65000000",
X"4c656674",
X"20666f72",
X"206f6e65",
X"20636869",
X"70000000",
X"52696768",
X"7420666f",
X"72207477",
X"6f206368",
X"69700000",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a257300",
X"45786974",
X"00000000",
X"35323030",
X"2e726f6d",
X"00000000",
X"524f4d00",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"00000000",
X"000067c4",
X"00006618",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"35323030",
X"00000000",
X"2f617461",
X"72353230",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
