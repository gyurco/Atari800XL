
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f1",
X"b0738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80f4",
X"e80c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f0",
X"f12d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580f0b0",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80da8604",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"775193b0",
X"3f83e080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3380f4f0",
X"0b80f4f0",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"52775192",
X"df3f83e0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583e0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"55b3933f",
X"83e08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"811451b2",
X"ab3f83e0",
X"80083070",
X"83e08008",
X"07802583",
X"e0800c53",
X"863d0d04",
X"fc3d0d76",
X"70525599",
X"cc3f83e0",
X"80085481",
X"5383e080",
X"0880c738",
X"7451998f",
X"3f83e080",
X"080b0b80",
X"f2f05383",
X"e0800852",
X"53ff8f3f",
X"83e08008",
X"a5380b0b",
X"80f2f452",
X"7251fefe",
X"3f83e080",
X"0894380b",
X"0b80f2f8",
X"527251fe",
X"ed3f83e0",
X"8008802e",
X"83388154",
X"73537283",
X"e0800c86",
X"3d0d04fd",
X"3d0d7570",
X"525498e5",
X"3f815383",
X"e0800898",
X"38735198",
X"ae3f83e0",
X"a0085283",
X"e0800851",
X"feb43f83",
X"e0800853",
X"7283e080",
X"0c853d0d",
X"04e03d0d",
X"a33d0870",
X"525e8ed3",
X"3f83e080",
X"0833943d",
X"56547394",
X"3880f7ec",
X"52745184",
X"c7397d52",
X"785191d6",
X"3f84d139",
X"7d518ebb",
X"3f83e080",
X"08527451",
X"8deb3f83",
X"e0a80852",
X"933d7052",
X"5d94c63f",
X"83e08008",
X"59800b83",
X"e0800855",
X"5b83e080",
X"087b2e94",
X"38811b74",
X"525b97c8",
X"3f83e080",
X"085483e0",
X"8008ee38",
X"805aff7a",
X"437a427a",
X"415f7909",
X"709f2c7b",
X"065b547a",
X"7a248438",
X"ff1b5af6",
X"1a700970",
X"9f2c7206",
X"7bff125a",
X"5a525555",
X"80752595",
X"38765197",
X"873f83e0",
X"800876ff",
X"18585557",
X"738024ed",
X"38747f2e",
X"873880c2",
X"993f745f",
X"78ff1b70",
X"585d5880",
X"7a259538",
X"775196dc",
X"3f83e080",
X"0876ff18",
X"58555873",
X"8024ed38",
X"800b83e7",
X"bc0c800b",
X"83e7dc0c",
X"0b0b80f2",
X"fc518bae",
X"3f81800b",
X"83e7dc0c",
X"0b0b80f3",
X"84518b9e",
X"3fa80b83",
X"e7bc0c76",
X"802e80e8",
X"3883e7bc",
X"08777932",
X"70307072",
X"07802570",
X"872b83e7",
X"dc0c5156",
X"78535656",
X"968f3f83",
X"e0800880",
X"2e8a380b",
X"0b80f38c",
X"518ae33f",
X"765195cf",
X"3f83e080",
X"08520b0b",
X"80f49851",
X"8ad03f76",
X"5195d53f",
X"83e08008",
X"83e7bc08",
X"55577574",
X"258638a8",
X"1656f739",
X"7583e7bc",
X"0c86f076",
X"24ff9438",
X"87980b83",
X"e7bc0c77",
X"802eb738",
X"7751958b",
X"3f83e080",
X"08785255",
X"95ab3f0b",
X"0b80f394",
X"5483e080",
X"088f3887",
X"39807634",
X"fd95390b",
X"0b80f390",
X"54745373",
X"520b0b80",
X"f2e45189",
X"e93f8054",
X"0b0b80f4",
X"e45189de",
X"3f811454",
X"73a82e09",
X"8106ed38",
X"868da051",
X"be9b3f80",
X"52903d70",
X"525480de",
X"f83f8352",
X"735180de",
X"f03f6180",
X"2e80ff38",
X"7b5473ff",
X"2e963878",
X"802e8180",
X"38785194",
X"ab3f83e0",
X"8008ff15",
X"5559e739",
X"78802e80",
X"eb387851",
X"94a73f83",
X"e0800880",
X"2efc8338",
X"785193ef",
X"3f83e080",
X"08520b0b",
X"80f2ec51",
X"abcd3f83",
X"e08008a4",
X"387c51ad",
X"853f83e0",
X"80085574",
X"ff165654",
X"807425fb",
X"ee38741d",
X"70335556",
X"73af2efe",
X"c838e839",
X"785193ad",
X"3f83e080",
X"08527c51",
X"acbc3ffb",
X"ce397f88",
X"29601005",
X"7a056105",
X"5afbff39",
X"a23d0d04",
X"803d0d90",
X"80f83370",
X"81ff0670",
X"842a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"a80b9080",
X"f834b80b",
X"9080f834",
X"7083e080",
X"0c823d0d",
X"04803d0d",
X"9080f833",
X"7081ff06",
X"70852a81",
X"32708106",
X"51515151",
X"70802e8d",
X"38980b90",
X"80f834b8",
X"0b9080f8",
X"347083e0",
X"800c823d",
X"0d04930b",
X"9080fc34",
X"ff0b9080",
X"e83404ff",
X"3d0d028f",
X"05335280",
X"0b9080fc",
X"348a51bb",
X"f03fdf3f",
X"80f80b90",
X"80e03480",
X"0b9080c8",
X"34fa1252",
X"719080c0",
X"34800b90",
X"80d83471",
X"9080d034",
X"9080f852",
X"807234b8",
X"7234833d",
X"0d04803d",
X"0d028b05",
X"33517090",
X"80f434fe",
X"bf3f83e0",
X"8008802e",
X"f638823d",
X"0d04803d",
X"0d853980",
X"c5ae3ffe",
X"d83f83e0",
X"8008802e",
X"f2389080",
X"f4337081",
X"ff0683e0",
X"800c5182",
X"3d0d0480",
X"3d0da30b",
X"9080fc34",
X"ff0b9080",
X"e8349080",
X"f851a871",
X"34b87134",
X"823d0d04",
X"803d0d90",
X"80fc3370",
X"81c00670",
X"30708025",
X"83e0800c",
X"51515182",
X"3d0d0480",
X"3d0d9080",
X"f8337081",
X"ff067083",
X"2a813270",
X"81065151",
X"51517080",
X"2ee838b0",
X"0b9080f8",
X"34b80b90",
X"80f83482",
X"3d0d0480",
X"3d0d9080",
X"ac088106",
X"83e0800c",
X"823d0d04",
X"fd3d0d75",
X"77545480",
X"73259438",
X"73708105",
X"55335280",
X"f3985185",
X"a13fff13",
X"53e93985",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"80dbd93f",
X"83e08008",
X"7a27ed38",
X"74802e80",
X"e0387452",
X"755180db",
X"c33f83e0",
X"80087553",
X"76525480",
X"dbc63f83",
X"e080087a",
X"53755256",
X"80dba93f",
X"83e08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"e08008c2",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9c",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fbfd3f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd13f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbad3f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83e0900c",
X"7183e094",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383e090",
X"085283e0",
X"940851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"99d25351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fd3d",
X"0d757052",
X"54a3c33f",
X"83e08008",
X"14537274",
X"2e9238ff",
X"13703353",
X"5371af2e",
X"098106ee",
X"38811353",
X"7283e080",
X"0c853d0d",
X"04fd3d0d",
X"75777053",
X"5454c73f",
X"83e08008",
X"732ea138",
X"83e08008",
X"733152ff",
X"125271ff",
X"2e8f3872",
X"70810554",
X"33747081",
X"055634eb",
X"39ff1454",
X"80743485",
X"3d0d0480",
X"3d0d7251",
X"ff903f82",
X"3d0d0471",
X"83e0800c",
X"04803d0d",
X"72518071",
X"34810bbc",
X"120c800b",
X"80c0120c",
X"823d0d04",
X"800b83e2",
X"d408248a",
X"38a4ad3f",
X"ff0b83e2",
X"d40c800b",
X"83e0800c",
X"04ff3d0d",
X"735283e0",
X"b008722e",
X"8d38d93f",
X"71519698",
X"3f7183e0",
X"b00c833d",
X"0d04f43d",
X"0d7e6062",
X"5c5a5581",
X"54bc1508",
X"81913874",
X"51cf3f79",
X"58807a25",
X"80f73883",
X"e3840870",
X"892a5783",
X"ff067884",
X"80723156",
X"56577378",
X"25833873",
X"557583e2",
X"d4082e84",
X"38ff893f",
X"83e2d408",
X"8025a638",
X"75892b51",
X"98db3f83",
X"e384088f",
X"3dfc1155",
X"5c548152",
X"f81b5196",
X"c53f7614",
X"83e3840c",
X"7583e2d4",
X"0c745376",
X"527851a2",
X"de3f83e0",
X"800883e3",
X"84081683",
X"e3840c78",
X"7631761b",
X"5b595677",
X"8024ff8b",
X"38617a71",
X"0c547554",
X"75802e83",
X"38815473",
X"83e0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"9b3f7651",
X"feaf3f86",
X"3dfc0553",
X"78527751",
X"95e83f79",
X"75710c54",
X"83e08008",
X"5483e080",
X"08802e83",
X"38815473",
X"83e0800c",
X"863d0d04",
X"fe3d0d75",
X"83e2d408",
X"53538072",
X"24893871",
X"732e8438",
X"fdd63f74",
X"51fdea3f",
X"725197ad",
X"3f83e080",
X"085283e0",
X"8008802e",
X"83388152",
X"7183e080",
X"0c843d0d",
X"04803d0d",
X"7280c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d72bc11",
X"0883e080",
X"0c51823d",
X"0d0480c4",
X"0b83e080",
X"0c04fd3d",
X"0d757771",
X"54705355",
X"539f9b3f",
X"82c81308",
X"bc150c82",
X"c0130880",
X"c0150cfc",
X"eb3f7351",
X"93aa3f73",
X"83e0b00c",
X"83e08008",
X"5383e080",
X"08802e83",
X"38815372",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"775553fc",
X"bf3f7280",
X"2ea538bc",
X"13085273",
X"519ea53f",
X"83e08008",
X"8f387752",
X"7251ff9a",
X"3f83e080",
X"08538a39",
X"82cc1308",
X"53d83981",
X"537283e0",
X"800c853d",
X"0d04fe3d",
X"0dff0b83",
X"e2d40c74",
X"83e0b40c",
X"7583e2d0",
X"0c9f923f",
X"83e08008",
X"81ff0652",
X"81537199",
X"3883e2ec",
X"518e943f",
X"83e08008",
X"5283e080",
X"08802e83",
X"38725271",
X"537283e0",
X"800c843d",
X"0d04fa3d",
X"0d787a82",
X"c4120882",
X"c4120870",
X"72245956",
X"56575773",
X"732e0981",
X"06913880",
X"c0165280",
X"c017519c",
X"963f83e0",
X"80085574",
X"83e0800c",
X"883d0d04",
X"f63d0d7c",
X"5b807b71",
X"5c54577a",
X"772e8c38",
X"811a82cc",
X"1408545a",
X"72f63880",
X"5980d939",
X"7a548157",
X"80707b7b",
X"315a5755",
X"ff185374",
X"732580c1",
X"3882cc14",
X"08527351",
X"ff8c3f80",
X"0b83e080",
X"0825a138",
X"82cc1408",
X"82cc1108",
X"82cc160c",
X"7482cc12",
X"0c537580",
X"2e863872",
X"82cc170c",
X"72548057",
X"7382cc15",
X"08811757",
X"5556ffb8",
X"39811959",
X"800bff1b",
X"54547873",
X"25833881",
X"54768132",
X"70750651",
X"5372ff90",
X"388c3d0d",
X"04f73d0d",
X"7b7d5a5a",
X"82d05283",
X"e2d00851",
X"80cee13f",
X"83e08008",
X"57f9e13f",
X"795283e2",
X"d85195b4",
X"3f83e080",
X"08548053",
X"83e08008",
X"732e0981",
X"06828338",
X"83e0b408",
X"0b0b80f2",
X"ec537052",
X"569bd33f",
X"0b0b80f2",
X"ec5280c0",
X"16519bc6",
X"3f75bc17",
X"0c7382c0",
X"170c810b",
X"82c4170c",
X"810b82c8",
X"170c7382",
X"cc170cff",
X"1782d017",
X"55578191",
X"3983e0c0",
X"3370822a",
X"70810651",
X"54557281",
X"80387481",
X"2a810658",
X"7780f638",
X"74842a81",
X"0682c415",
X"0c83e0c0",
X"33810682",
X"c8150c79",
X"5273519a",
X"ed3f7351",
X"9b843f83",
X"e0800814",
X"53af7370",
X"81055534",
X"72bc150c",
X"83e0c152",
X"72519ace",
X"3f83e0b8",
X"0882c015",
X"0c83e0ce",
X"5280c014",
X"519abb3f",
X"78802e8d",
X"38735178",
X"2d83e080",
X"08802e99",
X"387782cc",
X"150c7580",
X"2e863873",
X"82cc170c",
X"7382d015",
X"ff195955",
X"5676802e",
X"9b3883e0",
X"b85283e2",
X"d85194aa",
X"3f83e080",
X"088a3883",
X"e0c13353",
X"72fed238",
X"78802e89",
X"3883e0b4",
X"0851fcb8",
X"3f83e0b4",
X"08537283",
X"e0800c8b",
X"3d0d04ff",
X"3d0d8052",
X"7351fdb5",
X"3f833d0d",
X"04f03d0d",
X"62705254",
X"f6903f83",
X"e0800874",
X"53873d70",
X"535555f6",
X"b03ff790",
X"3f7351d3",
X"3f635374",
X"5283e080",
X"0851fab8",
X"3f923d0d",
X"047183e0",
X"800c0480",
X"c01283e0",
X"800c0480",
X"3d0d7282",
X"c0110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"82cc1108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"7282c411",
X"0883e080",
X"0c51823d",
X"0d04f93d",
X"0d7983e0",
X"98085757",
X"81772781",
X"96387688",
X"17082781",
X"8e387533",
X"5574822e",
X"89387483",
X"2eb33880",
X"fe397454",
X"761083fe",
X"06537688",
X"2a8c1708",
X"0552893d",
X"fc055199",
X"c03f83e0",
X"800880df",
X"38029d05",
X"33893d33",
X"71882b07",
X"565680d1",
X"39845476",
X"822b83fc",
X"06537687",
X"2a8c1708",
X"0552893d",
X"fc055199",
X"903f83e0",
X"8008b038",
X"029f0533",
X"0284059e",
X"05337198",
X"2b71902b",
X"07028c05",
X"9d053370",
X"882b7207",
X"8d3d3371",
X"80fffffe",
X"80060751",
X"52535758",
X"56833981",
X"557483e0",
X"800c893d",
X"0d04fb3d",
X"0d83e098",
X"08fe1988",
X"1208fe05",
X"55565480",
X"56747327",
X"8d388214",
X"33757129",
X"94160805",
X"57537583",
X"e0800c87",
X"3d0d04fc",
X"3d0d7652",
X"800b83e0",
X"98087033",
X"51525370",
X"832e0981",
X"06913895",
X"12339413",
X"3371982b",
X"71902b07",
X"5555519b",
X"12339a13",
X"3371882b",
X"07740783",
X"e0800c55",
X"863d0d04",
X"fc3d0d76",
X"83e09808",
X"55558075",
X"23881508",
X"5372812e",
X"88388814",
X"08732685",
X"388152b2",
X"39729038",
X"73335271",
X"832e0981",
X"06853890",
X"14085372",
X"8c160c72",
X"802e8d38",
X"7251fed6",
X"3f83e080",
X"08528539",
X"90140852",
X"7190160c",
X"80527183",
X"e0800c86",
X"3d0d04fa",
X"3d0d7883",
X"e0980871",
X"22810570",
X"83ffff06",
X"57545755",
X"73802e88",
X"38901508",
X"53728638",
X"835280e7",
X"39738f06",
X"527180da",
X"38811390",
X"160c8c15",
X"08537290",
X"38830b84",
X"17225752",
X"73762780",
X"c638bf39",
X"821633ff",
X"0574842a",
X"065271b2",
X"387251fc",
X"b13f8152",
X"7183e080",
X"0827a838",
X"835283e0",
X"80088817",
X"08279c38",
X"83e08008",
X"8c160c83",
X"e0800851",
X"fdbc3f83",
X"e0800890",
X"160c7375",
X"23805271",
X"83e0800c",
X"883d0d04",
X"f23d0d60",
X"6264585e",
X"5b753355",
X"74a02e09",
X"81068838",
X"81167044",
X"56ef3962",
X"70335656",
X"74af2e09",
X"81068438",
X"81164380",
X"0b881c0c",
X"62703351",
X"55749f26",
X"91387a51",
X"fdd23f83",
X"e0800856",
X"807d3483",
X"8139933d",
X"841c0870",
X"58595f8a",
X"55a07670",
X"81055834",
X"ff155574",
X"ff2e0981",
X"06ef3880",
X"705a5c88",
X"7f085f5a",
X"7b811d70",
X"81ff0660",
X"13703370",
X"af327030",
X"a0732771",
X"80250751",
X"51525b53",
X"5e575574",
X"80e73876",
X"ae2e0981",
X"06833881",
X"55787a27",
X"75075574",
X"802e9f38",
X"79883270",
X"3078ae32",
X"70307073",
X"079f2a53",
X"51575156",
X"75bb3888",
X"598b5aff",
X"ab397698",
X"2b557480",
X"25873880",
X"f0c01733",
X"57ff9f17",
X"55749926",
X"8938e017",
X"7081ff06",
X"58557881",
X"1a7081ff",
X"06721b53",
X"5b575576",
X"7534fef8",
X"397b1e7f",
X"0c805576",
X"a0268338",
X"8155748b",
X"19347a51",
X"fc823f83",
X"e0800880",
X"f538a054",
X"7a227085",
X"2b83e006",
X"5455901b",
X"08527c51",
X"93cb3f83",
X"e0800857",
X"83e08008",
X"8181387c",
X"33557480",
X"2e80f438",
X"8b1d3370",
X"832a7081",
X"06515656",
X"74b4388b",
X"7d841d08",
X"83e08008",
X"595b5b58",
X"ff185877",
X"ff2e9a38",
X"79708105",
X"5b337970",
X"81055b33",
X"71713152",
X"56567580",
X"2ee23886",
X"3975802e",
X"96387a51",
X"fbe53fff",
X"863983e0",
X"80085683",
X"e08008b6",
X"38833976",
X"56841b08",
X"8b113351",
X"5574a738",
X"8b1d3370",
X"842a7081",
X"06515656",
X"74893883",
X"56943981",
X"5690397c",
X"51fa943f",
X"83e08008",
X"881c0cfd",
X"81397583",
X"e0800c90",
X"3d0d04f8",
X"3d0d7a7c",
X"59578254",
X"83fe5377",
X"52765192",
X"903f8356",
X"83e08008",
X"80ec3881",
X"17337733",
X"71882b07",
X"56568256",
X"7482d4d5",
X"2e098106",
X"80d43875",
X"54b65377",
X"52765191",
X"e43f83e0",
X"80089838",
X"81173377",
X"3371882b",
X"0783e080",
X"08525656",
X"748182c6",
X"2eac3882",
X"5480d253",
X"77527651",
X"91bb3f83",
X"e0800898",
X"38811733",
X"77337188",
X"2b0783e0",
X"80085256",
X"56748182",
X"c62e8338",
X"81567583",
X"e0800c8a",
X"3d0d04eb",
X"3d0d675a",
X"800b83e0",
X"980c90dd",
X"3f83e080",
X"08810655",
X"82567483",
X"ee387475",
X"538f3d70",
X"535759fe",
X"ca3f83e0",
X"800881ff",
X"06577681",
X"2e098106",
X"80d43890",
X"5483be53",
X"74527551",
X"90cf3f83",
X"e0800880",
X"c9388f3d",
X"33557480",
X"2e80c938",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"0770587b",
X"575e525e",
X"575957fd",
X"ee3f83e0",
X"800881ff",
X"06577683",
X"2e098106",
X"86388156",
X"82f13976",
X"802e8638",
X"865682e7",
X"39a4548d",
X"53785275",
X"518fe63f",
X"815683e0",
X"800882d3",
X"3802be05",
X"33028405",
X"bd053371",
X"882b0759",
X"5d77ab38",
X"0280ce05",
X"33028405",
X"80cd0533",
X"71982b71",
X"902b0797",
X"3d337088",
X"2b720702",
X"940580cb",
X"05337107",
X"54525e57",
X"595602b7",
X"05337871",
X"29028805",
X"b6053302",
X"8c05b505",
X"3371882b",
X"07701d70",
X"7f8c050c",
X"5f595759",
X"5d8e3d33",
X"821b3402",
X"b9053390",
X"3d337188",
X"2b075a5c",
X"78841b23",
X"02bb0533",
X"028405ba",
X"05337188",
X"2b07565c",
X"74ab3802",
X"80ca0533",
X"02840580",
X"c9053371",
X"982b7190",
X"2b07963d",
X"3370882b",
X"72070294",
X"0580c705",
X"33710751",
X"5253575e",
X"5c747631",
X"78317984",
X"2a903d33",
X"54717131",
X"535656bf",
X"c73f83e0",
X"80088205",
X"70881c0c",
X"83e08008",
X"e08a0556",
X"567483df",
X"fe268338",
X"825783ff",
X"f6762785",
X"38835789",
X"39865676",
X"802e80db",
X"38767a34",
X"76832e09",
X"8106b038",
X"0280d605",
X"33028405",
X"80d50533",
X"71982b71",
X"902b0799",
X"3d337088",
X"2b720702",
X"940580d3",
X"05337107",
X"7f90050c",
X"525e5758",
X"56863977",
X"1b901b0c",
X"841a228c",
X"1b081971",
X"842a0594",
X"1c0c5d80",
X"0b811b34",
X"7983e098",
X"0c805675",
X"83e0800c",
X"973d0d04",
X"e93d0d83",
X"e0980856",
X"85547580",
X"2e818238",
X"800b8117",
X"34993de0",
X"11466a54",
X"8a3d7054",
X"58ec0551",
X"f6e63f83",
X"e0800854",
X"83e08008",
X"80df3889",
X"3d335473",
X"802e9138",
X"02ab0533",
X"70842a81",
X"06515574",
X"802e8638",
X"835480c1",
X"397651f4",
X"8a3f83e0",
X"8008a017",
X"0c02bf05",
X"33028405",
X"be053371",
X"982b7190",
X"2b07028c",
X"05bd0533",
X"70882b72",
X"07953d33",
X"71079c1c",
X"0c527898",
X"1b0c5356",
X"5957810b",
X"81173474",
X"547383e0",
X"800c993d",
X"0d04f53d",
X"0d7d7f61",
X"7283e098",
X"085a5d5d",
X"595c807b",
X"0c855775",
X"802e81e0",
X"38811633",
X"81065584",
X"5774802e",
X"81d23891",
X"39748117",
X"34863980",
X"0b811734",
X"815781c0",
X"399c1608",
X"98170831",
X"55747827",
X"83387458",
X"77802e81",
X"a9389816",
X"087083ff",
X"06565774",
X"80cf3882",
X"1633ff05",
X"77892a06",
X"7081ff06",
X"5a5578a0",
X"38768738",
X"a0160855",
X"8d39a416",
X"0851f0ea",
X"3f83e080",
X"08558175",
X"27ffa838",
X"74a4170c",
X"a4160851",
X"f2843f83",
X"e0800855",
X"83e08008",
X"802eff89",
X"3883e080",
X"0819a817",
X"0c981608",
X"83ff0684",
X"80713151",
X"55777527",
X"83387755",
X"7483ffff",
X"06549816",
X"0883ff06",
X"53a81608",
X"5279577b",
X"83387b57",
X"76518a8d",
X"3f83e080",
X"08fed038",
X"98160815",
X"98170c74",
X"1a787631",
X"7c08177d",
X"0c595afe",
X"d3398057",
X"7683e080",
X"0c8d3d0d",
X"04fa3d0d",
X"7883e098",
X"08555685",
X"5573802e",
X"81e13881",
X"14338106",
X"53845572",
X"802e81d3",
X"389c1408",
X"53727627",
X"83387256",
X"98140857",
X"800b9815",
X"0c75802e",
X"81b73882",
X"14337089",
X"2b565376",
X"802eb538",
X"7452ff16",
X"51bac93f",
X"83e08008",
X"ff187654",
X"70535853",
X"baba3f83",
X"e0800873",
X"26963874",
X"30707806",
X"7098170c",
X"777131a4",
X"17085258",
X"51538939",
X"a0140870",
X"a4160c53",
X"747627b9",
X"387251ee",
X"d93f83e0",
X"80085381",
X"0b83e080",
X"08278b38",
X"88140883",
X"e0800826",
X"8838800b",
X"811534b0",
X"3983e080",
X"08a4150c",
X"98140815",
X"98150c75",
X"753156c4",
X"39981408",
X"16709816",
X"0c735256",
X"efc83f83",
X"e080088c",
X"3883e080",
X"08811534",
X"81559439",
X"821433ff",
X"0576892a",
X"0683e080",
X"0805a815",
X"0c805574",
X"83e0800c",
X"883d0d04",
X"ef3d0d63",
X"56855583",
X"e0980880",
X"2e80d238",
X"933df405",
X"84170c64",
X"53883d70",
X"53765257",
X"f1d23f83",
X"e0800855",
X"83e08008",
X"b438883d",
X"33547380",
X"2ea13802",
X"a7053370",
X"842a7081",
X"06515555",
X"83557380",
X"2e973876",
X"51eef83f",
X"83e08008",
X"88170c75",
X"51efa93f",
X"83e08008",
X"557483e0",
X"800c933d",
X"0d04e43d",
X"0d6ea13d",
X"08405e85",
X"5683e098",
X"08802e84",
X"85389e3d",
X"f405841f",
X"0c7e9838",
X"7d51eef8",
X"3f83e080",
X"085683ee",
X"39814181",
X"f6398341",
X"81f13993",
X"3d7f9605",
X"4159807f",
X"8295055e",
X"56756081",
X"ff053483",
X"41901e08",
X"762e81d3",
X"38a0547d",
X"2270852b",
X"83e00654",
X"58901e08",
X"52785186",
X"983f83e0",
X"80084183",
X"e08008ff",
X"b8387833",
X"5c7b802e",
X"ffb4388b",
X"193370bf",
X"06718106",
X"52435574",
X"802e80de",
X"387b81bf",
X"0655748f",
X"2480d338",
X"9a193355",
X"7480cb38",
X"f31d7058",
X"5d815675",
X"8b2e0981",
X"0685388e",
X"568b3975",
X"9a2e0981",
X"0683389c",
X"56751970",
X"70810552",
X"33713381",
X"1a821a5f",
X"5b525b55",
X"74863879",
X"77348539",
X"80df7734",
X"777b5757",
X"7aa02e09",
X"8106c038",
X"81567b81",
X"e5327030",
X"709f2a51",
X"51557bae",
X"2e933874",
X"802e8e38",
X"61832a70",
X"81065155",
X"74802e97",
X"387d51ed",
X"e23f83e0",
X"80084183",
X"e0800887",
X"38901e08",
X"feaf3880",
X"60347580",
X"2e88387c",
X"527f5183",
X"a53f6080",
X"2e863880",
X"0b901f0c",
X"60566083",
X"2e853860",
X"81d03889",
X"1f57901e",
X"08802e81",
X"a8388056",
X"75197033",
X"515574a0",
X"2ea03874",
X"852e0981",
X"06843881",
X"e5557477",
X"70810559",
X"34811670",
X"81ff0657",
X"55877627",
X"d7388819",
X"335574a0",
X"2ea938ae",
X"77708105",
X"59348856",
X"75197033",
X"515574a0",
X"2e953874",
X"77708105",
X"59348116",
X"7081ff06",
X"57558a76",
X"27e2388b",
X"19337f88",
X"05349f19",
X"339e1a33",
X"71982b71",
X"902b079d",
X"1c337088",
X"2b72079c",
X"1e337107",
X"640c5299",
X"1d33981e",
X"3371882b",
X"07535153",
X"57595674",
X"7f840523",
X"97193396",
X"1a337188",
X"2b075656",
X"747f8605",
X"23807734",
X"7d51ebf3",
X"3f83e080",
X"08833270",
X"30707207",
X"9f2c83e0",
X"80080652",
X"5656961f",
X"3355748a",
X"38891f52",
X"961f5181",
X"b13f7583",
X"e0800c9e",
X"3d0d04fd",
X"3d0d7577",
X"53547333",
X"51708938",
X"71335170",
X"802ea138",
X"73337233",
X"52537271",
X"278538ff",
X"51943970",
X"73278538",
X"81518b39",
X"81148113",
X"5354d339",
X"80517083",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"54547233",
X"7081ff06",
X"52527080",
X"2ea33871",
X"81ff0681",
X"14ffbf12",
X"53545270",
X"99268938",
X"a0127081",
X"ff065351",
X"71747081",
X"055634d2",
X"39807434",
X"853d0d04",
X"ffbd3d0d",
X"80c63d08",
X"52a53d70",
X"5254ffb3",
X"3f80c73d",
X"0852853d",
X"705253ff",
X"a63f7252",
X"7351fedf",
X"3f80c53d",
X"0d04fe3d",
X"0d747653",
X"53717081",
X"05533351",
X"70737081",
X"05553470",
X"f038843d",
X"0d04fe3d",
X"0d745280",
X"72335253",
X"70732e8d",
X"38811281",
X"14713353",
X"545270f5",
X"387283e0",
X"800c843d",
X"0d04fc3d",
X"0d765574",
X"83e39808",
X"2eaf3880",
X"53745187",
X"c13f83e0",
X"800881ff",
X"06ff1470",
X"81ff0672",
X"30709f2a",
X"51525553",
X"5472802e",
X"843871dd",
X"3873fe38",
X"7483e398",
X"0c863d0d",
X"04ff3d0d",
X"ff0b83e3",
X"980c84a5",
X"3f815187",
X"853f83e0",
X"800881ff",
X"065271ee",
X"3881d33f",
X"7183e080",
X"0c833d0d",
X"04fc3d0d",
X"76028405",
X"a2052202",
X"8805a605",
X"227a5455",
X"5555ff82",
X"3f72802e",
X"a03883e3",
X"ac143375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552dd",
X"39800b83",
X"e0800c86",
X"3d0d04fc",
X"3d0d7678",
X"7a115653",
X"55805371",
X"742e9338",
X"72155170",
X"3383e3ac",
X"13348112",
X"81145452",
X"ea39800b",
X"83e0800c",
X"863d0d04",
X"fd3d0d90",
X"5483e398",
X"085186f4",
X"3f83e080",
X"0881ff06",
X"ff157130",
X"71307073",
X"079f2a72",
X"9f2a0652",
X"55525553",
X"72db3885",
X"3d0d0480",
X"3d0d83e3",
X"a4081083",
X"e39c0807",
X"9080a80c",
X"823d0d04",
X"800b83e3",
X"a40ce43f",
X"04810b83",
X"e3a40cdb",
X"3f04ed3f",
X"047183e3",
X"a00c0480",
X"3d0d8051",
X"f43f810b",
X"83e3a40c",
X"810b83e3",
X"9c0cffbb",
X"3f823d0d",
X"04803d0d",
X"72307074",
X"07802583",
X"e39c0c51",
X"ffa53f82",
X"3d0d0480",
X"3d0d028b",
X"05339080",
X"a40c9080",
X"a8087081",
X"06515170",
X"f5389080",
X"a4087081",
X"ff0683e0",
X"800c5182",
X"3d0d0480",
X"3d0d81ff",
X"51d13f83",
X"e0800881",
X"ff0683e0",
X"800c823d",
X"0d04803d",
X"0d73902b",
X"73079080",
X"b40c823d",
X"0d0404fb",
X"3d0d7802",
X"84059f05",
X"3370982b",
X"55575572",
X"80259b38",
X"7580ff06",
X"56805280",
X"f751e03f",
X"83e08008",
X"81ff0654",
X"73812680",
X"ff388051",
X"fee73fff",
X"a23f8151",
X"fedf3fff",
X"9a3f7551",
X"feed3f74",
X"982a51fe",
X"e63f7490",
X"2a7081ff",
X"065253fe",
X"da3f7488",
X"2a7081ff",
X"065253fe",
X"ce3f7481",
X"ff0651fe",
X"c63f8155",
X"7580c02e",
X"09810686",
X"38819555",
X"8d397580",
X"c82e0981",
X"06843881",
X"87557451",
X"fea53f8a",
X"55fec83f",
X"83e08008",
X"81ff0670",
X"982b5454",
X"7280258c",
X"38ff1570",
X"81ff0656",
X"5374e238",
X"7383e080",
X"0c873d0d",
X"04fa3d0d",
X"fdc53f80",
X"51fdda3f",
X"8a54fe93",
X"3fff1470",
X"81ff0655",
X"5373f338",
X"73745355",
X"80c051fe",
X"a63f83e0",
X"800881ff",
X"06547381",
X"2e098106",
X"829f3883",
X"aa5280c8",
X"51fe8c3f",
X"83e08008",
X"81ff0653",
X"72812e09",
X"810681a8",
X"38745487",
X"3d741154",
X"56fdc83f",
X"83e08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e53802",
X"9a053353",
X"72812e09",
X"810681d9",
X"38029b05",
X"335380ce",
X"90547281",
X"aa2e8d38",
X"81c73980",
X"e4518a89",
X"3fff1454",
X"73802e81",
X"b838820a",
X"5281e951",
X"fda53f83",
X"e0800881",
X"ff065372",
X"de387252",
X"80fa51fd",
X"923f83e0",
X"800881ff",
X"06537281",
X"90387254",
X"731653fc",
X"d63f83e0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e8",
X"38873d33",
X"70862a70",
X"81065154",
X"548c5572",
X"80e33884",
X"5580de39",
X"745281e9",
X"51fccc3f",
X"83e08008",
X"81ff0653",
X"825581e9",
X"56817327",
X"86387355",
X"80c15680",
X"ce90548a",
X"3980e451",
X"88fb3fff",
X"14547380",
X"2ea93880",
X"527551fc",
X"9a3f83e0",
X"800881ff",
X"065372e1",
X"38848052",
X"80d051fc",
X"863f83e0",
X"800881ff",
X"06537280",
X"2e833880",
X"557483e3",
X"a8348051",
X"fb873ffb",
X"c23f883d",
X"0d04fb3d",
X"0d775480",
X"0b83e3a8",
X"3370832a",
X"70810651",
X"55575572",
X"752e0981",
X"06853873",
X"892b5473",
X"5280d151",
X"fbbd3f83",
X"e0800881",
X"ff065372",
X"bd3882b8",
X"c054fb83",
X"3f83e080",
X"0881ff06",
X"537281ff",
X"2e098106",
X"8938ff14",
X"5473e738",
X"9f397281",
X"fe2e0981",
X"06963883",
X"e7ac5283",
X"e3ac51fa",
X"ed3ffad3",
X"3ffad03f",
X"83398155",
X"8051fa89",
X"3ffac43f",
X"7481ff06",
X"83e0800c",
X"873d0d04",
X"fb3d0d77",
X"83e3ac56",
X"548151f9",
X"ec3f83e3",
X"a8337083",
X"2a708106",
X"51545672",
X"85387389",
X"2b547352",
X"80d851fa",
X"b63f83e0",
X"800881ff",
X"06537280",
X"e43881ff",
X"51f9d43f",
X"81fe51f9",
X"ce3f8480",
X"53747081",
X"05563351",
X"f9c13fff",
X"137083ff",
X"ff065153",
X"72eb3872",
X"51f9b03f",
X"7251f9ab",
X"3ff9d03f",
X"83e08008",
X"9f0653a7",
X"88547285",
X"2e8c3899",
X"3980e451",
X"86b33fff",
X"1454f9b3",
X"3f83e080",
X"0881ff2e",
X"843873e9",
X"388051f8",
X"e43ff99f",
X"3f800b83",
X"e0800c87",
X"3d0d0471",
X"83e7b00c",
X"8880800b",
X"83e7ac0c",
X"8480800b",
X"83e7b40c",
X"04fd3d0d",
X"77701755",
X"7705ff1a",
X"535371ff",
X"2e943873",
X"70810555",
X"33517073",
X"70810555",
X"34ff1252",
X"e939853d",
X"0d04fc3d",
X"0d87a681",
X"55743383",
X"e7b834a0",
X"5483a080",
X"5383e7b0",
X"085283e7",
X"ac0851ff",
X"b83fa054",
X"83a48053",
X"83e7b008",
X"5283e7ac",
X"0851ffa5",
X"3f905483",
X"a8805383",
X"e7b00852",
X"83e7ac08",
X"51ff923f",
X"a0538052",
X"83e7b408",
X"83a08005",
X"51858b3f",
X"a0538052",
X"83e7b408",
X"83a48005",
X"5184fb3f",
X"90538052",
X"83e7b408",
X"83a88005",
X"5184eb3f",
X"ff753483",
X"a0805480",
X"5383e7b0",
X"085283e7",
X"b40851fe",
X"cc3f80d0",
X"805483b0",
X"805383e7",
X"b0085283",
X"e7b40851",
X"feb73f86",
X"913fa254",
X"805383e7",
X"b4088c80",
X"055280f5",
X"e451fea1",
X"3f860b87",
X"a8833480",
X"0b87a882",
X"34800b87",
X"a09a34af",
X"0b87a096",
X"34bf0b87",
X"a0973480",
X"0b87a098",
X"349f0b87",
X"a0993480",
X"0b87a09b",
X"34e00b87",
X"a88934a2",
X"0b87a880",
X"34830b87",
X"a48f3482",
X"0b87a881",
X"34863d0d",
X"04fd3d0d",
X"83a08054",
X"805383e7",
X"b4085283",
X"e7b00851",
X"fdbf3f80",
X"d0805483",
X"b0805383",
X"e7b40852",
X"83e7b008",
X"51fdaa3f",
X"a05483a0",
X"805383e7",
X"b4085283",
X"e7b00851",
X"fd973fa0",
X"5483a480",
X"5383e7b4",
X"085283e7",
X"b00851fd",
X"843f9054",
X"83a88053",
X"83e7b408",
X"5283e7b0",
X"0851fcf1",
X"3f83e7b8",
X"3387a681",
X"34853d0d",
X"04803d0d",
X"90809008",
X"810683e0",
X"800c823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087081",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fd0676",
X"1007720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870822c",
X"bf0683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe830676",
X"822b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087088",
X"2c870683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f1ff06",
X"76882b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"8b2cbf06",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f88f",
X"ff06768b",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870912c",
X"bf0683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fc87ffff",
X"0676912b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90808008",
X"70882c81",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"0870892c",
X"810683e0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708a",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8b2c8106",
X"83e0800c",
X"51823d0d",
X"04fe3d0d",
X"7481e629",
X"872a9080",
X"a00c843d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"81055434",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727084",
X"05540cff",
X"1151f039",
X"843d0d04",
X"fe3d0d84",
X"80805380",
X"5288800a",
X"51ffb33f",
X"81808053",
X"80528280",
X"0a51c63f",
X"843d0d04",
X"803d0d81",
X"51fcbf3f",
X"72802e83",
X"38d23f81",
X"51fcdd3f",
X"8051fcd8",
X"3f8051fc",
X"a93f823d",
X"0d04fd3d",
X"0d755280",
X"5480ff72",
X"25883881",
X"0bff8013",
X"5354ffbf",
X"12517099",
X"268638e0",
X"12529e39",
X"ff9f1251",
X"99712795",
X"38d012e0",
X"13705454",
X"51897127",
X"88388f73",
X"27833880",
X"5273802e",
X"85388180",
X"12527181",
X"ff0683e0",
X"800c853d",
X"0d04803d",
X"0d84d8c0",
X"51807170",
X"81055334",
X"7084e0c0",
X"2e098106",
X"f038823d",
X"0d04fe3d",
X"0d029705",
X"3351ff86",
X"3f83e080",
X"0881ff06",
X"83e7bc08",
X"54528073",
X"249b3883",
X"e7d80813",
X"7283e7dc",
X"08075353",
X"71733483",
X"e7bc0881",
X"0583e7bc",
X"0c843d0d",
X"04fa3d0d",
X"82800a1b",
X"55805788",
X"3dfc0554",
X"79537452",
X"7851cca4",
X"3f883d0d",
X"04fe3d0d",
X"83e7d408",
X"527451d3",
X"883f83e0",
X"80088c38",
X"76537552",
X"83e7d408",
X"51c73f84",
X"3d0d04fe",
X"3d0d83e7",
X"d4085375",
X"527451cd",
X"c73f83e0",
X"80088d38",
X"77537652",
X"83e7d408",
X"51ffa23f",
X"843d0d04",
X"fe3d0d83",
X"e7d40851",
X"ccbb3f83",
X"e0800881",
X"80802e09",
X"81068838",
X"83c18080",
X"539b3983",
X"e7d40851",
X"cc9f3f83",
X"e0800880",
X"d0802e09",
X"81069338",
X"83c1b080",
X"5383e080",
X"085283e7",
X"d40851fe",
X"d83f843d",
X"0d04803d",
X"0dfab43f",
X"83e08008",
X"842980f6",
X"88057008",
X"83e0800c",
X"51823d0d",
X"04ee3d0d",
X"80438042",
X"80418070",
X"5a5bfdd2",
X"3f800b83",
X"e7bc0c80",
X"0b83e7dc",
X"0c80f3e4",
X"51c78b3f",
X"81800b83",
X"e7dc0c80",
X"f3e851c6",
X"fd3f80d0",
X"0b83e7bc",
X"0c783070",
X"7a078025",
X"70872b83",
X"e7dc0c51",
X"55f9a73f",
X"83e08008",
X"5280f3f0",
X"51c6d73f",
X"80f80b83",
X"e7bc0c78",
X"81327030",
X"70720780",
X"2570872b",
X"83e7dc0c",
X"515656fe",
X"f13f83e0",
X"80085280",
X"f3fc51c6",
X"ad3f81a0",
X"0b83e7bc",
X"0c788232",
X"70307072",
X"07802570",
X"872b83e7",
X"dc0c5156",
X"83e7d408",
X"5256c7c7",
X"3f83e080",
X"085280f4",
X"8451c5fe",
X"3f81f00b",
X"83e7bc0c",
X"810b83e7",
X"c05b5883",
X"e7bc0882",
X"197a3270",
X"30707207",
X"80257087",
X"2b83e7dc",
X"0c51578e",
X"3d7055ff",
X"1b545757",
X"5799913f",
X"79708405",
X"5b0851c6",
X"fe3f7454",
X"83e08008",
X"53775280",
X"f48c51c5",
X"b13fa817",
X"83e7bc0c",
X"81185877",
X"852e0981",
X"06ffb038",
X"83900b83",
X"e7bc0c78",
X"87327030",
X"70720780",
X"2570872b",
X"83e7dc0c",
X"515656f8",
X"cd3f80f4",
X"9c5583e0",
X"8008802e",
X"8e3883e7",
X"d00851c6",
X"aa3f83e0",
X"80085574",
X"5280f4a4",
X"51c4df3f",
X"83e00b83",
X"e7bc0c78",
X"88327030",
X"70720780",
X"2570872b",
X"83e7dc0c",
X"515780f4",
X"b05255c4",
X"bd3f868d",
X"a051f985",
X"3f805291",
X"3d705255",
X"99e33f83",
X"52745199",
X"dc3f6119",
X"59788025",
X"85388059",
X"90398879",
X"25853888",
X"59873978",
X"882682db",
X"3878822b",
X"5580f2c0",
X"150804f6",
X"c13f83e0",
X"80086157",
X"5575812e",
X"09810689",
X"3883e080",
X"08105590",
X"3975ff2e",
X"09810688",
X"3883e080",
X"08812c55",
X"90752585",
X"38905588",
X"39748024",
X"83388155",
X"7451f69b",
X"3f829039",
X"f6ad3f83",
X"e0800861",
X"05557480",
X"25853880",
X"55883987",
X"75258338",
X"87557451",
X"f6a63f81",
X"ee396087",
X"3862802e",
X"81e53883",
X"e0a40883",
X"e0a00c8b",
X"df0b83e0",
X"a80c83e7",
X"d40851ff",
X"b5db3ffa",
X"e73f81c7",
X"39605680",
X"76259938",
X"8af80b83",
X"e0a80c83",
X"e7b41570",
X"085255ff",
X"b5bb3f74",
X"08529139",
X"75802591",
X"3883e7b4",
X"150851c4",
X"983f8052",
X"fd1951b8",
X"3962802e",
X"818d3883",
X"e7b41570",
X"0883e7c0",
X"08720c83",
X"e7c00cfd",
X"1a705351",
X"558b813f",
X"83e08008",
X"5680518a",
X"f73f83e0",
X"80085274",
X"51878f3f",
X"75528051",
X"87883f80",
X"d6396055",
X"807525b8",
X"3883e0ac",
X"0883e0a0",
X"0c8bdf0b",
X"83e0a80c",
X"83e7d008",
X"51ffb4c5",
X"3f83e7d0",
X"0851ffb1",
X"df3f83e0",
X"800881ff",
X"06705255",
X"f5b13f74",
X"802e9c38",
X"8155a039",
X"74802593",
X"3883e7d0",
X"0851c389",
X"3f8051f5",
X"963f8439",
X"6287387a",
X"802efa8a",
X"38805574",
X"83e0800c",
X"943d0d04",
X"fe3d0df5",
X"943f83e0",
X"8008802e",
X"86388051",
X"80f739f5",
X"993f83e0",
X"800880eb",
X"38f5b93f",
X"83e08008",
X"802eaa38",
X"8151f2f6",
X"3fefef3f",
X"800b83e7",
X"bc0cf9b9",
X"3f83e080",
X"0853ff0b",
X"83e7bc0c",
X"f1db3f72",
X"be387251",
X"f2d43fbc",
X"39f4f03f",
X"83e08008",
X"802eb138",
X"8151f2c2",
X"3fefbb3f",
X"8af80b83",
X"e0a80c83",
X"e7c00851",
X"ffb38a3f",
X"ff0b83e7",
X"bc0cf1a5",
X"3f83e7c0",
X"08528051",
X"85983f81",
X"51f5d13f",
X"843d0d04",
X"fc3d0d90",
X"80805286",
X"84808051",
X"c5dc3f83",
X"e0800880",
X"c33888e9",
X"3f80f7dc",
X"51ca9c3f",
X"83e08008",
X"559c800a",
X"5480c080",
X"5380f4b8",
X"5283e080",
X"0851f79f",
X"3f83e7d4",
X"085380f4",
X"c8527451",
X"c4e63f83",
X"e0800884",
X"38f7ad3f",
X"8151f4f8",
X"3f92f53f",
X"8151f4f0",
X"3ffe913f",
X"fc3983e0",
X"8c080283",
X"e08c0cfb",
X"3d0d0280",
X"f4d40b83",
X"e0a40c80",
X"f4d80b83",
X"e09c0c80",
X"f4dc0b83",
X"e0ac0c83",
X"e08c08fc",
X"050c800b",
X"83e7c00b",
X"83e08c08",
X"f8050c83",
X"e08c08f4",
X"050cc3be",
X"3f83e080",
X"088605fc",
X"0683e08c",
X"08f0050c",
X"0283e08c",
X"08f00508",
X"310d833d",
X"7083e08c",
X"08f80508",
X"70840583",
X"e08c08f8",
X"050c0c51",
X"c0873f83",
X"e08c08f4",
X"05088105",
X"83e08c08",
X"f4050c83",
X"e08c08f4",
X"0508862e",
X"098106ff",
X"ad388694",
X"808051ec",
X"d23fff0b",
X"83e7bc0c",
X"800b83e7",
X"dc0c84d8",
X"c00b83e7",
X"d80c8151",
X"effc3f81",
X"51f0a13f",
X"8051f09c",
X"3f8151f0",
X"c23f8151",
X"f1973f82",
X"51f0e53f",
X"8051f1bb",
X"3f80d082",
X"528051ff",
X"bdc53ffd",
X"bf3f83e0",
X"8c08fc05",
X"080d800b",
X"83e0800c",
X"873d0d83",
X"e08c0c04",
X"803d0d81",
X"ff51800b",
X"83e7e812",
X"34ff1151",
X"70f43882",
X"3d0d04ff",
X"3d0d7370",
X"33535181",
X"11337134",
X"71811234",
X"833d0d04",
X"fb3d0d77",
X"79565680",
X"70715555",
X"52717525",
X"ac387216",
X"70337014",
X"7081ff06",
X"55515151",
X"71742789",
X"38811270",
X"81ff0653",
X"51718114",
X"7083ffff",
X"06555254",
X"747324d6",
X"387183e0",
X"800c873d",
X"0d04fc3d",
X"0d7655ff",
X"b6f13f83",
X"e0800880",
X"2ef53883",
X"ea840886",
X"057081ff",
X"065253ff",
X"b4f13f84",
X"39fb813f",
X"ffb6d03f",
X"83e08008",
X"812ef238",
X"80547315",
X"53ffb5b6",
X"3f83e080",
X"08733481",
X"14547385",
X"2e098106",
X"e9388439",
X"fad63fff",
X"b6a53f83",
X"e0800880",
X"2ef23874",
X"3383e7e8",
X"34811533",
X"83e7e934",
X"82153383",
X"e7ea3483",
X"153383e7",
X"eb348452",
X"83e7e851",
X"feba3f83",
X"e0800881",
X"ff068416",
X"33565372",
X"752e0981",
X"068d38ff",
X"b59a3f83",
X"e0800880",
X"2e9a3883",
X"ea8408a8",
X"2e098106",
X"8938860b",
X"83ea840c",
X"8739a80b",
X"83ea840c",
X"80e451ef",
X"d43f863d",
X"0d04f43d",
X"0d7e6059",
X"55805d80",
X"75822b71",
X"83ea8812",
X"0c83ea9c",
X"175b5b57",
X"76793477",
X"772e83b8",
X"38765277",
X"51ffbed0",
X"3f8e3dfc",
X"05549053",
X"83e9f052",
X"7751ffbe",
X"8b3f7c56",
X"75902e09",
X"81068394",
X"3883e9f0",
X"51fd943f",
X"83e9f251",
X"fd8d3f83",
X"e9f451fd",
X"863f7683",
X"ea800c77",
X"51ffbbd7",
X"3f80f2f4",
X"5283e080",
X"0851ffab",
X"913f83e0",
X"8008812e",
X"09810680",
X"d4387683",
X"ea980c82",
X"0b83e9f0",
X"34ff960b",
X"83e9f134",
X"7751ffbe",
X"9c3f83e0",
X"80085583",
X"e0800877",
X"25883883",
X"e080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583e9f2",
X"347483e9",
X"f3347683",
X"e9f434ff",
X"800b83e9",
X"f5348190",
X"3983e9f0",
X"3383e9f1",
X"3371882b",
X"07565b74",
X"83ffff2e",
X"09810680",
X"e838fe80",
X"0b83ea98",
X"0c810b83",
X"ea800cff",
X"0b83e9f0",
X"34ff0b83",
X"e9f13477",
X"51ffbda9",
X"3f83e080",
X"0883eaa0",
X"0c83e080",
X"085583e0",
X"80088025",
X"883883e0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83e9f234",
X"7483e9f3",
X"347683e9",
X"f434ff80",
X"0b83e9f5",
X"34810b83",
X"e9ff34a5",
X"39748596",
X"2e098106",
X"80fe3875",
X"83ea980c",
X"7751ffbc",
X"dd3f83e9",
X"ff3383e0",
X"80080755",
X"7483e9ff",
X"3483e9ff",
X"33810655",
X"74802e83",
X"38845783",
X"e9f43383",
X"e9f53371",
X"882b0756",
X"5c748180",
X"2e098106",
X"a13883e9",
X"f23383e9",
X"f3337188",
X"2b07565b",
X"ad807527",
X"87387682",
X"07579c39",
X"76810757",
X"96397482",
X"802e0981",
X"06873876",
X"83075787",
X"397481ff",
X"268a3877",
X"83ea881b",
X"0c767934",
X"8e3d0d04",
X"803d0d72",
X"842983ea",
X"88057008",
X"83e0800c",
X"51823d0d",
X"04fe3d0d",
X"800b83e9",
X"ec0c800b",
X"83e9e80c",
X"ff0b83e7",
X"e40ca80b",
X"83ea840c",
X"ae51ffaf",
X"ba3f800b",
X"83ea8854",
X"52807370",
X"8405550c",
X"81125271",
X"842e0981",
X"06ef3884",
X"3d0d04fe",
X"3d0d7402",
X"84059605",
X"22535371",
X"802e9738",
X"72708105",
X"543351ff",
X"afc43fff",
X"127083ff",
X"ff065152",
X"e639843d",
X"0d04fe3d",
X"0d029205",
X"225382ac",
X"51eae63f",
X"80c351ff",
X"afa03f81",
X"9651ead9",
X"3f725283",
X"e7e851ff",
X"b23f7252",
X"83e7e851",
X"f8ee3f83",
X"e0800881",
X"ff0651ff",
X"aefc3f84",
X"3d0d04ff",
X"b13d0d80",
X"d13df805",
X"51f9973f",
X"83e9ec08",
X"810583e9",
X"ec0c80cf",
X"3d33cf11",
X"7081ff06",
X"51565674",
X"832688ed",
X"38758f06",
X"ff055675",
X"83e7e408",
X"2e9b3875",
X"83269638",
X"7583e7e4",
X"0c758429",
X"83ea8805",
X"70085355",
X"7551fa96",
X"3f807624",
X"88c93875",
X"842983ea",
X"88055574",
X"08802e88",
X"ba3883e7",
X"e4088429",
X"83ea8805",
X"70080288",
X"0582b905",
X"33525b55",
X"7480d22e",
X"84b13874",
X"80d22490",
X"3874bf2e",
X"9c387480",
X"d02e81d7",
X"3887f839",
X"7480d32e",
X"80d23874",
X"80d72e81",
X"c63887e7",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055656",
X"ffadf83f",
X"80c151ff",
X"adb03ff6",
X"e73f860b",
X"83e7e834",
X"815283e7",
X"e851ffae",
X"d33f8151",
X"fde43f74",
X"8938860b",
X"83ea840c",
X"8739a80b",
X"83ea840c",
X"ffadc43f",
X"80c151ff",
X"acfc3ff6",
X"b33f900b",
X"83e9ff33",
X"81065656",
X"74802e83",
X"38985683",
X"e9f43383",
X"e9f53371",
X"882b0756",
X"59748180",
X"2e098106",
X"9c3883e9",
X"f23383e9",
X"f3337188",
X"2b075657",
X"ad807527",
X"8c387581",
X"80075685",
X"3975a007",
X"567583e7",
X"e834ff0b",
X"83e7e934",
X"e00b83e7",
X"ea34800b",
X"83e7eb34",
X"845283e7",
X"e851ffad",
X"c73f8451",
X"869e3902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"5659ffac",
X"b63f7951",
X"ffb7a33f",
X"83e08008",
X"802e8b38",
X"80ce51ff",
X"abe03f85",
X"f23980c1",
X"51ffabd6",
X"3fffaccb",
X"3fffaafe",
X"3f83ea98",
X"08588375",
X"259b3883",
X"e9f43383",
X"e9f53371",
X"882b07fc",
X"1771297a",
X"05838005",
X"5a51578d",
X"39748180",
X"2918ff80",
X"05588180",
X"57805676",
X"762e9338",
X"ffabaf3f",
X"83e08008",
X"83e7e817",
X"34811656",
X"ea39ffab",
X"9d3f83e0",
X"800881ff",
X"06775383",
X"e7e85256",
X"f4d63f83",
X"e0800881",
X"ff065575",
X"752e0981",
X"06818a38",
X"ffab9c3f",
X"80c151ff",
X"aad43fff",
X"abc93f77",
X"527951ff",
X"b5b23f80",
X"5e80d13d",
X"fdf40554",
X"765383e7",
X"e8527951",
X"ffb3bf3f",
X"0282b905",
X"33558158",
X"7480d72e",
X"098106bd",
X"3880d13d",
X"fdf00554",
X"76538f3d",
X"70537a52",
X"59ffb4c4",
X"3f805676",
X"762ea238",
X"751983e7",
X"e8173371",
X"33707232",
X"70307080",
X"2570307e",
X"06811d5d",
X"5e515151",
X"525b55db",
X"3982ac51",
X"e59f3f77",
X"802e8638",
X"80c35184",
X"3980ce51",
X"ffa9cf3f",
X"ffaac43f",
X"ffa8f73f",
X"83dd3902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"59558070",
X"5d59ffa9",
X"ea3f80c1",
X"51ffa9a2",
X"3f83ea80",
X"08792e82",
X"de3883ea",
X"a00880fc",
X"055580fd",
X"52745186",
X"d73f83e0",
X"80085b77",
X"8224b238",
X"ff187087",
X"2b83ffff",
X"800680f6",
X"a80583e7",
X"e8595755",
X"81805575",
X"70810557",
X"33777081",
X"055934ff",
X"157081ff",
X"06515574",
X"ea38828d",
X"397782e8",
X"2e81ab38",
X"7782e92e",
X"09810681",
X"b23880f4",
X"e051ffaf",
X"a53f7858",
X"77873270",
X"30707207",
X"80257a8a",
X"32703070",
X"72078025",
X"73075354",
X"5a515755",
X"75802e97",
X"38787826",
X"9238a00b",
X"83e7e81a",
X"34811970",
X"81ff065a",
X"55eb3981",
X"187081ff",
X"0659558a",
X"7827ffbc",
X"388f5883",
X"e7e31833",
X"83e7e819",
X"34ff1870",
X"81ff0659",
X"55778426",
X"ea389058",
X"800b83e7",
X"e8193481",
X"187081ff",
X"0670982b",
X"52595574",
X"8025e938",
X"80c6557a",
X"858f2484",
X"3880c255",
X"7483e7e8",
X"3480f10b",
X"83e7eb34",
X"810b83e7",
X"ec347a83",
X"e7e9347a",
X"882c5574",
X"83e7ea34",
X"80cb3982",
X"f0782580",
X"c4387780",
X"fd29fd97",
X"d3055279",
X"51ffb1e0",
X"3f80d13d",
X"fdec0554",
X"80fd5383",
X"e7e85279",
X"51ffb198",
X"3f7b8119",
X"59567580",
X"fc248338",
X"78587788",
X"2c557483",
X"e8e53477",
X"83e8e634",
X"7583e8e7",
X"34818059",
X"80cc3983",
X"ea980857",
X"8378259b",
X"3883e9f4",
X"3383e9f5",
X"3371882b",
X"07fc1a71",
X"29790583",
X"80055951",
X"598d3977",
X"81802917",
X"ff800557",
X"81805976",
X"527951ff",
X"b0ee3f80",
X"d13dfdec",
X"05547853",
X"83e7e852",
X"7951ffb0",
X"a73f7851",
X"f6b83fff",
X"a6e13fff",
X"a5943f8b",
X"3983e9e8",
X"08810583",
X"e9e80c80",
X"d13d0d04",
X"f6d93feb",
X"9f3ff939",
X"fc3d0d76",
X"78718429",
X"83ea8805",
X"70085153",
X"5353709e",
X"3880ce72",
X"3480cf0b",
X"81133480",
X"ce0b8213",
X"3480c50b",
X"83133470",
X"84133480",
X"e73983ea",
X"9c133354",
X"80d27234",
X"73822a70",
X"81065151",
X"80cf5370",
X"843880d7",
X"53728113",
X"34a00b82",
X"13347383",
X"06517081",
X"2e9e3870",
X"81248838",
X"70802e8f",
X"389f3970",
X"822e9238",
X"70832e92",
X"38933980",
X"d8558e39",
X"80d35589",
X"3980cd55",
X"843980c4",
X"55748313",
X"3480c40b",
X"84133480",
X"0b851334",
X"863d0d04",
X"fd3d0d75",
X"5380730c",
X"800b8414",
X"0c800b88",
X"140c87a6",
X"80337081",
X"ff067081",
X"2a813271",
X"81327181",
X"06718106",
X"3184180c",
X"55567083",
X"2a813271",
X"822a8132",
X"71810671",
X"81063177",
X"0c525451",
X"5187a090",
X"33700981",
X"0688150c",
X"51853d0d",
X"04fe3d0d",
X"74765452",
X"7151ffa0",
X"3f72812e",
X"a2388173",
X"268d3872",
X"822eab38",
X"72832e9f",
X"38e63971",
X"08e23884",
X"1208dd38",
X"881208d8",
X"38a03988",
X"1208812e",
X"098106cc",
X"38943988",
X"1208812e",
X"8d387108",
X"89388412",
X"08802eff",
X"b738843d",
X"0d04fc3d",
X"0d767853",
X"54815380",
X"55873971",
X"10731054",
X"52737226",
X"5172802e",
X"a7387080",
X"2e863871",
X"8025e838",
X"72802e98",
X"38717426",
X"89387372",
X"31757407",
X"56547281",
X"2a72812a",
X"5353e539",
X"73517883",
X"38745170",
X"83e0800c",
X"863d0d04",
X"fe3d0d80",
X"53755274",
X"51ffa33f",
X"843d0d04",
X"fe3d0d81",
X"53755274",
X"51ff933f",
X"843d0d04",
X"fb3d0d77",
X"79555580",
X"56747625",
X"86387430",
X"55815673",
X"80258838",
X"73307681",
X"32575480",
X"53735274",
X"51fee73f",
X"83e08008",
X"5475802e",
X"873883e0",
X"80083054",
X"7383e080",
X"0c873d0d",
X"04fa3d0d",
X"787a5755",
X"80577477",
X"25863874",
X"30558157",
X"759f2c54",
X"81537574",
X"32743152",
X"7451feaa",
X"3f83e080",
X"08547680",
X"2e873883",
X"e0800830",
X"547383e0",
X"800c883d",
X"0d040000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002ab3",
X"00002af4",
X"00002b16",
X"00002b3d",
X"00002b3d",
X"00002b3d",
X"00002b3d",
X"00002bae",
X"00002c00",
X"25732025",
X"73000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"6e616d65",
X"20000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"000039a0",
X"000039a4",
X"000039ac",
X"000039b8",
X"000039c4",
X"000039d0",
X"000039dc",
X"000039e0",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
