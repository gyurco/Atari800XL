
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80ea",
X"e0738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80ee",
X"a40c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580e8",
X"9a2d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580e7d9",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80d1b104",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"775193b0",
X"3f83e080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3380eeac",
X"0b80eeac",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"52775192",
X"df3f83e0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583e0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"55b3963f",
X"83e08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"811451b2",
X"ae3f83e0",
X"80083070",
X"83e08008",
X"07802583",
X"e0800c53",
X"863d0d04",
X"fc3d0d76",
X"70525599",
X"cd3f83e0",
X"80085481",
X"5383e080",
X"0880c738",
X"74519990",
X"3f83e080",
X"080b0b80",
X"eca05383",
X"e0800852",
X"53ff8f3f",
X"83e08008",
X"a5380b0b",
X"80eca452",
X"7251fefe",
X"3f83e080",
X"0894380b",
X"0b80eca8",
X"527251fe",
X"ed3f83e0",
X"8008802e",
X"83388154",
X"73537283",
X"e0800c86",
X"3d0d04fd",
X"3d0d7570",
X"525498e6",
X"3f815383",
X"e0800898",
X"38735198",
X"af3f83e0",
X"a0085283",
X"e0800851",
X"feb43f83",
X"e0800853",
X"7283e080",
X"0c853d0d",
X"04e03d0d",
X"a33d0870",
X"525e8ed1",
X"3f83e080",
X"0833943d",
X"56547394",
X"3880f1a8",
X"52745184",
X"c6397d52",
X"785191d6",
X"3f84d039",
X"7d518eb9",
X"3f83e080",
X"08527451",
X"8de93f83",
X"e0a80852",
X"933d7052",
X"5d94c73f",
X"83e08008",
X"59800b83",
X"e0800855",
X"5b83e080",
X"087b2e94",
X"38811b74",
X"525b97c9",
X"3f83e080",
X"085483e0",
X"8008ee38",
X"805aff7a",
X"437a427a",
X"415f7909",
X"709f2c7b",
X"065b547a",
X"7a248438",
X"ff1b5af6",
X"1a700970",
X"9f2c7206",
X"7bff125a",
X"5a525555",
X"80752595",
X"38765197",
X"883f83e0",
X"800876ff",
X"18585557",
X"738024ed",
X"38747f2e",
X"8638b8db",
X"3f745f78",
X"ff1b7058",
X"5d58807a",
X"25953877",
X"5196de3f",
X"83e08008",
X"76ff1858",
X"55587380",
X"24ed3880",
X"0b83e3ac",
X"0c800b83",
X"e3d00c0b",
X"0b80ecac",
X"518bad3f",
X"81800b83",
X"e3d00c0b",
X"0b80ecb4",
X"518b9d3f",
X"a80b83e3",
X"ac0c7680",
X"2e80e838",
X"83e3ac08",
X"77793270",
X"30707207",
X"80257087",
X"2b83e3d0",
X"0c515678",
X"53565696",
X"913f83e0",
X"8008802e",
X"8a380b0b",
X"80ecbc51",
X"8ae23f76",
X"5195d13f",
X"83e08008",
X"520b0b80",
X"edc8518a",
X"cf3f7651",
X"95d73f83",
X"e0800883",
X"e3ac0855",
X"57757425",
X"8638a816",
X"56f73975",
X"83e3ac0c",
X"86f07624",
X"ff943887",
X"980b83e3",
X"ac0c7780",
X"2eb73877",
X"51958d3f",
X"83e08008",
X"78525595",
X"ad3f0b0b",
X"80ecc454",
X"83e08008",
X"8f388739",
X"807634fd",
X"96390b0b",
X"80ecc054",
X"74537352",
X"0b0b80ec",
X"945189e8",
X"3f80540b",
X"0b80eea0",
X"5189dd3f",
X"81145473",
X"a82e0981",
X"06ed3886",
X"8da051b4",
X"d03f8052",
X"903d7052",
X"5480d6a2",
X"3f835273",
X"5180d69a",
X"3f61802e",
X"80ff387b",
X"5473ff2e",
X"96387880",
X"2e818038",
X"785194ad",
X"3f83e080",
X"08ff1555",
X"59e73978",
X"802e80eb",
X"38785194",
X"a93f83e0",
X"8008802e",
X"fc843878",
X"5193f13f",
X"83e08008",
X"520b0b80",
X"ec9c51ab",
X"d13f83e0",
X"8008a438",
X"7c51ad89",
X"3f83e080",
X"085574ff",
X"16565480",
X"7425fbef",
X"38741d70",
X"33555673",
X"af2efec8",
X"38e83978",
X"5193af3f",
X"83e08008",
X"527c51ac",
X"c03ffbcf",
X"397f8829",
X"6010057a",
X"0561055a",
X"fc8039a2",
X"3d0d0480",
X"3d0d9080",
X"f8337081",
X"ff067084",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d38a8",
X"0b9080f8",
X"34b80b90",
X"80f83470",
X"83e0800c",
X"823d0d04",
X"803d0d90",
X"80f83370",
X"81ff0670",
X"852a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"980b9080",
X"f834b80b",
X"9080f834",
X"7083e080",
X"0c823d0d",
X"04930b90",
X"80fc34ff",
X"0b9080e8",
X"3404ff3d",
X"0d028f05",
X"3352800b",
X"9080fc34",
X"8a51b2a5",
X"3fdf3f80",
X"f80b9080",
X"e034800b",
X"9080c834",
X"fa125271",
X"9080c034",
X"800b9080",
X"d8347190",
X"80d03490",
X"80f85280",
X"7234b872",
X"34833d0d",
X"04803d0d",
X"028b0533",
X"51709080",
X"f434febf",
X"3f83e080",
X"08802ef6",
X"38823d0d",
X"04803d0d",
X"8439bbf1",
X"3ffed93f",
X"83e08008",
X"802ef338",
X"9080f433",
X"7081ff06",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"a30b9080",
X"fc34ff0b",
X"9080e834",
X"9080f851",
X"a87134b8",
X"7134823d",
X"0d04803d",
X"0d9080fc",
X"337081c0",
X"06703070",
X"802583e0",
X"800c5151",
X"51823d0d",
X"04803d0d",
X"9080f833",
X"7081ff06",
X"70832a81",
X"32708106",
X"51515151",
X"70802ee8",
X"38b00b90",
X"80f834b8",
X"0b9080f8",
X"34823d0d",
X"04803d0d",
X"9080ac08",
X"810683e0",
X"800c823d",
X"0d04fd3d",
X"0d757754",
X"54807325",
X"94387370",
X"81055533",
X"5280ecc8",
X"5185a13f",
X"ff1353e9",
X"39853d0d",
X"04f63d0d",
X"7c7e6062",
X"5a5d5b56",
X"80598155",
X"8539747a",
X"29557452",
X"755180d3",
X"843f83e0",
X"80087a27",
X"ed387480",
X"2e80e038",
X"74527551",
X"80d2ee3f",
X"83e08008",
X"75537652",
X"5480d2f1",
X"3f83e080",
X"087a5375",
X"525680d2",
X"d43f83e0",
X"80087930",
X"707b079f",
X"2a707780",
X"24075151",
X"54557287",
X"3883e080",
X"08c23876",
X"8118b016",
X"55585889",
X"74258b38",
X"b714537a",
X"853880d7",
X"14537278",
X"34811959",
X"ff9c3980",
X"77348c3d",
X"0d04f73d",
X"0d7b7d7f",
X"62029005",
X"bb053357",
X"59565a5a",
X"b0587283",
X"38a05875",
X"70708105",
X"52337159",
X"54559039",
X"8074258e",
X"38ff1477",
X"70810559",
X"33545472",
X"ef3873ff",
X"15555380",
X"73258938",
X"77527951",
X"782def39",
X"75337557",
X"5372802e",
X"90387252",
X"7951782d",
X"75708105",
X"573353ed",
X"398b3d0d",
X"04ee3d0d",
X"64666969",
X"70708105",
X"52335b4a",
X"5c5e5e76",
X"802e82f9",
X"3876a52e",
X"09810682",
X"e0388070",
X"41677070",
X"81055233",
X"714a5957",
X"5f76b02e",
X"0981068c",
X"38757081",
X"05573376",
X"4857815f",
X"d0175675",
X"892680da",
X"3876675c",
X"59805c93",
X"39778a24",
X"80c3387b",
X"8a29187b",
X"7081055d",
X"335a5cd0",
X"197081ff",
X"06585889",
X"7727a438",
X"ff9f1970",
X"81ff06ff",
X"a91b5a51",
X"56857627",
X"9238ffbf",
X"197081ff",
X"06515675",
X"85268a38",
X"c9195877",
X"8025ffb9",
X"387a477b",
X"407881ff",
X"06577680",
X"e42e80e5",
X"387680e4",
X"24a73876",
X"80d82e81",
X"86387680",
X"d8249038",
X"76802e81",
X"cc3876a5",
X"2e81b638",
X"81b93976",
X"80e32e81",
X"8c3881af",
X"397680f5",
X"2e9b3876",
X"80f5248b",
X"387680f3",
X"2e818138",
X"81993976",
X"80f82e80",
X"ca38818f",
X"39913d70",
X"55578053",
X"8a527984",
X"1b710853",
X"5b56fbfd",
X"3f7655ab",
X"3979841b",
X"7108943d",
X"705b5b52",
X"5b567580",
X"258c3875",
X"3056ad78",
X"340280c1",
X"05577654",
X"80538a52",
X"7551fbd1",
X"3f77557e",
X"54b83991",
X"3d705577",
X"80d83270",
X"30708025",
X"56515856",
X"90527984",
X"1b710853",
X"5b57fbad",
X"3f7555db",
X"3979841b",
X"83123354",
X"5b569839",
X"79841b71",
X"08575b56",
X"80547f53",
X"7c527d51",
X"fc9c3f87",
X"3976527d",
X"517c2d66",
X"70335881",
X"0547fd83",
X"39943d0d",
X"047283e0",
X"900c7183",
X"e0940c04",
X"fb3d0d88",
X"3d707084",
X"05520857",
X"54755383",
X"e0900852",
X"83e09408",
X"51fcc63f",
X"873d0d04",
X"ff3d0d73",
X"70085351",
X"02930533",
X"72347008",
X"8105710c",
X"833d0d04",
X"fc3d0d87",
X"3d881155",
X"785499d0",
X"5351fc99",
X"3f805287",
X"3d51d13f",
X"863d0d04",
X"fd3d0d75",
X"705254a3",
X"c83f83e0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83e0",
X"8008732e",
X"a13883e0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183e0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83e2d408",
X"248b3880",
X"cf943fff",
X"0b83e2d4",
X"0c800b83",
X"e0800c04",
X"ff3d0d73",
X"5283e0b0",
X"08722e8d",
X"38d83f71",
X"51969c3f",
X"7183e0b0",
X"0c833d0d",
X"04f43d0d",
X"7e60625c",
X"5a558154",
X"bc150881",
X"92387451",
X"cf3f7958",
X"807a2580",
X"f83883e3",
X"84087089",
X"2a5783ff",
X"06788480",
X"72315656",
X"57737825",
X"83387355",
X"7583e2d4",
X"082e8438",
X"ff883f83",
X"e2d40880",
X"25a63875",
X"892b5198",
X"df3f83e3",
X"84088f3d",
X"fc11555c",
X"548152f8",
X"1b5196c9",
X"3f761483",
X"e3840c75",
X"83e2d40c",
X"74537652",
X"785180cd",
X"a63f83e0",
X"800883e3",
X"84081683",
X"e3840c78",
X"7631761b",
X"5b595677",
X"8024ff8a",
X"38617a71",
X"0c547554",
X"75802e83",
X"38815473",
X"83e0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"993f7651",
X"feae3f86",
X"3dfc0553",
X"78527751",
X"95eb3f79",
X"75710c54",
X"83e08008",
X"5483e080",
X"08802e83",
X"38815473",
X"83e0800c",
X"863d0d04",
X"fe3d0d75",
X"83e2d408",
X"53538072",
X"24893871",
X"732e8438",
X"fdd43f74",
X"51fde93f",
X"725197b0",
X"3f83e080",
X"085283e0",
X"8008802e",
X"83388152",
X"7183e080",
X"0c843d0d",
X"04803d0d",
X"7280c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d72bc11",
X"0883e080",
X"0c51823d",
X"0d0480c4",
X"0b83e080",
X"0c04fd3d",
X"0d757771",
X"54705355",
X"539f9e3f",
X"82c81308",
X"bc150c82",
X"c0130880",
X"c0150cfc",
X"e93f7351",
X"93ad3f73",
X"83e0b00c",
X"83e08008",
X"5383e080",
X"08802e83",
X"38815372",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"775553fc",
X"bd3f7280",
X"2ea538bc",
X"13085273",
X"519ea83f",
X"83e08008",
X"8f387752",
X"7251ff9a",
X"3f83e080",
X"08538a39",
X"82cc1308",
X"53d83981",
X"537283e0",
X"800c853d",
X"0d04fe3d",
X"0dff0b83",
X"e2d40c74",
X"83e0b40c",
X"7583e2d0",
X"0c80c9e9",
X"3f83e080",
X"0881ff06",
X"52815371",
X"993883e2",
X"ec518e96",
X"3f83e080",
X"085283e0",
X"8008802e",
X"83387252",
X"71537283",
X"e0800c84",
X"3d0d04fa",
X"3d0d787a",
X"82c41208",
X"82c41208",
X"70722459",
X"56565757",
X"73732e09",
X"81069138",
X"80c01652",
X"80c01751",
X"9c983f83",
X"e0800855",
X"7483e080",
X"0c883d0d",
X"04f63d0d",
X"7c5b807b",
X"715c5457",
X"7a772e8c",
X"38811a82",
X"cc140854",
X"5a72f638",
X"805980d9",
X"397a5481",
X"5780707b",
X"7b315a57",
X"55ff1853",
X"74732580",
X"c13882cc",
X"14085273",
X"51ff8c3f",
X"800b83e0",
X"800825a1",
X"3882cc14",
X"0882cc11",
X"0882cc16",
X"0c7482cc",
X"120c5375",
X"802e8638",
X"7282cc17",
X"0c725480",
X"577382cc",
X"15088117",
X"575556ff",
X"b8398119",
X"59800bff",
X"1b545478",
X"73258338",
X"81547681",
X"32707506",
X"515372ff",
X"90388c3d",
X"0d04f73d",
X"0d7b7d5a",
X"5a82d052",
X"83e2d008",
X"5180c689",
X"3f83e080",
X"0857f9de",
X"3f795283",
X"e2d85195",
X"b63f83e0",
X"80085480",
X"5383e080",
X"08732e09",
X"81068283",
X"3883e0b4",
X"080b0b80",
X"ec9c5370",
X"52569bd5",
X"3f0b0b80",
X"ec9c5280",
X"c016519b",
X"c83f75bc",
X"170c7382",
X"c0170c81",
X"0b82c417",
X"0c810b82",
X"c8170c73",
X"82cc170c",
X"ff1782d0",
X"17555781",
X"913983e0",
X"c0337082",
X"2a708106",
X"51545572",
X"81803874",
X"812a8106",
X"587780f6",
X"3874842a",
X"810682c4",
X"150c83e0",
X"c0338106",
X"82c8150c",
X"79527351",
X"9aef3f73",
X"519b863f",
X"83e08008",
X"1453af73",
X"70810555",
X"3472bc15",
X"0c83e0c1",
X"5272519a",
X"d03f83e0",
X"b80882c0",
X"150c83e0",
X"ce5280c0",
X"14519abd",
X"3f78802e",
X"8d387351",
X"782d83e0",
X"8008802e",
X"99387782",
X"cc150c75",
X"802e8638",
X"7382cc17",
X"0c7382d0",
X"15ff1959",
X"55567680",
X"2e9b3883",
X"e0b85283",
X"e2d85194",
X"ac3f83e0",
X"80088a38",
X"83e0c133",
X"5372fed2",
X"3878802e",
X"893883e0",
X"b40851fc",
X"b83f83e0",
X"b4085372",
X"83e0800c",
X"8b3d0d04",
X"ff3d0d80",
X"527351fd",
X"b53f833d",
X"0d04f03d",
X"0d627052",
X"54f68d3f",
X"83e08008",
X"7453873d",
X"70535555",
X"f6ad3ff7",
X"8d3f7351",
X"d33f6353",
X"745283e0",
X"800851fa",
X"b73f923d",
X"0d047183",
X"e0800c04",
X"80c01283",
X"e0800c04",
X"803d0d72",
X"82c01108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"7282cc11",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282c4",
X"110883e0",
X"800c5182",
X"3d0d04f9",
X"3d0d7983",
X"e0980857",
X"57817727",
X"81983876",
X"88170827",
X"81903875",
X"33557482",
X"2e893874",
X"832eb438",
X"81803974",
X"54761083",
X"fe065376",
X"882a8c17",
X"08055289",
X"3dfc0551",
X"80c4833f",
X"83e08008",
X"80e03802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d23984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"5180c3d2",
X"3f83e080",
X"08b03802",
X"9f053302",
X"84059e05",
X"3371982b",
X"71902b07",
X"028c059d",
X"05337088",
X"2b72078d",
X"3d337180",
X"fffffe80",
X"06075152",
X"53575856",
X"83398155",
X"7483e080",
X"0c893d0d",
X"04fb3d0d",
X"83e09808",
X"fe198812",
X"08fe0555",
X"56548056",
X"7473278d",
X"38821433",
X"75712994",
X"16080557",
X"537583e0",
X"800c873d",
X"0d04fc3d",
X"0d765280",
X"0b83e098",
X"08703351",
X"52537083",
X"2e098106",
X"91389512",
X"33941333",
X"71982b71",
X"902b0755",
X"55519b12",
X"339a1333",
X"71882b07",
X"740783e0",
X"800c5586",
X"3d0d04fc",
X"3d0d7683",
X"e0980855",
X"55807523",
X"88150853",
X"72812e88",
X"38881408",
X"73268538",
X"8152b239",
X"72903873",
X"33527183",
X"2e098106",
X"85389014",
X"0853728c",
X"160c7280",
X"2e8d3872",
X"51fed63f",
X"83e08008",
X"52853990",
X"14085271",
X"90160c80",
X"527183e0",
X"800c863d",
X"0d04fa3d",
X"0d7883e0",
X"98087122",
X"81057083",
X"ffff0657",
X"54575573",
X"802e8838",
X"90150853",
X"72863883",
X"5280e739",
X"738f0652",
X"7180da38",
X"81139016",
X"0c8c1508",
X"53729038",
X"830b8417",
X"22575273",
X"762780c6",
X"38bf3982",
X"1633ff05",
X"74842a06",
X"5271b238",
X"7251fcaf",
X"3f815271",
X"83e08008",
X"27a83883",
X"5283e080",
X"08881708",
X"279c3883",
X"e080088c",
X"160c83e0",
X"800851fd",
X"bc3f83e0",
X"80089016",
X"0c737523",
X"80527183",
X"e0800c88",
X"3d0d04f2",
X"3d0d6062",
X"64585e5b",
X"75335574",
X"a02e0981",
X"06883881",
X"16704456",
X"ef396270",
X"33565674",
X"af2e0981",
X"06843881",
X"1643800b",
X"881c0c62",
X"70335155",
X"749f2691",
X"387a51fd",
X"d23f83e0",
X"80085680",
X"7d348381",
X"39933d84",
X"1c087058",
X"595f8a55",
X"a0767081",
X"055834ff",
X"155574ff",
X"2e098106",
X"ef388070",
X"5a5c887f",
X"085f5a7b",
X"811d7081",
X"ff066013",
X"703370af",
X"327030a0",
X"73277180",
X"25075151",
X"525b535e",
X"57557480",
X"e73876ae",
X"2e098106",
X"83388155",
X"787a2775",
X"07557480",
X"2e9f3879",
X"88327030",
X"78ae3270",
X"30707307",
X"9f2a5351",
X"57515675",
X"bb388859",
X"8b5affab",
X"3976982b",
X"55748025",
X"873880e9",
X"f0173357",
X"ff9f1755",
X"74992689",
X"38e01770",
X"81ff0658",
X"5578811a",
X"7081ff06",
X"721b535b",
X"57557675",
X"34fef839",
X"7b1e7f0c",
X"805576a0",
X"26833881",
X"55748b19",
X"347a51fc",
X"823f83e0",
X"800880f5",
X"38a0547a",
X"2270852b",
X"83e00654",
X"55901b08",
X"527c51be",
X"8d3f83e0",
X"80085783",
X"e0800881",
X"81387c33",
X"5574802e",
X"80f4388b",
X"1d337083",
X"2a708106",
X"51565674",
X"b4388b7d",
X"841d0883",
X"e0800859",
X"5b5b58ff",
X"185877ff",
X"2e9a3879",
X"7081055b",
X"33797081",
X"055b3371",
X"71315256",
X"5675802e",
X"e2388639",
X"75802e96",
X"387a51fb",
X"e53fff86",
X"3983e080",
X"085683e0",
X"8008b638",
X"83397656",
X"841b088b",
X"11335155",
X"74a7388b",
X"1d337084",
X"2a708106",
X"51565674",
X"89388356",
X"94398156",
X"90397c51",
X"fa943f83",
X"e0800888",
X"1c0cfd81",
X"397583e0",
X"800c903d",
X"0d04f83d",
X"0d7a7c59",
X"57825483",
X"fe537752",
X"7651bcd2",
X"3f835683",
X"e0800880",
X"ec388117",
X"33773371",
X"882b0756",
X"56825674",
X"82d4d52e",
X"09810680",
X"d4387554",
X"b6537752",
X"7651bca6",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"ac388254",
X"80d25377",
X"527651bb",
X"fd3f83e0",
X"80089838",
X"81173377",
X"3371882b",
X"0783e080",
X"08525656",
X"748182c6",
X"2e833881",
X"567583e0",
X"800c8a3d",
X"0d04eb3d",
X"0d675a80",
X"0b83e098",
X"0cbbb23f",
X"83e08008",
X"81065582",
X"567483ee",
X"38747553",
X"8f3d7053",
X"5759feca",
X"3f83e080",
X"0881ff06",
X"5776812e",
X"09810680",
X"d4389054",
X"83be5374",
X"527551bb",
X"913f83e0",
X"800880c9",
X"388f3d33",
X"5574802e",
X"80c93802",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"70587b57",
X"5e525e57",
X"5957fdee",
X"3f83e080",
X"0881ff06",
X"5776832e",
X"09810686",
X"38815682",
X"f1397680",
X"2e863886",
X"5682e739",
X"a4548d53",
X"78527551",
X"baa83f81",
X"5683e080",
X"0882d338",
X"02be0533",
X"028405bd",
X"05337188",
X"2b07595d",
X"77ab3802",
X"80ce0533",
X"02840580",
X"cd053371",
X"982b7190",
X"2b07973d",
X"3370882b",
X"72070294",
X"0580cb05",
X"33710754",
X"525e5759",
X"5602b705",
X"33787129",
X"028805b6",
X"0533028c",
X"05b50533",
X"71882b07",
X"701d707f",
X"8c050c5f",
X"5957595d",
X"8e3d3382",
X"1b3402b9",
X"0533903d",
X"3371882b",
X"075a5c78",
X"841b2302",
X"bb053302",
X"8405ba05",
X"3371882b",
X"07565c74",
X"ab380280",
X"ca053302",
X"840580c9",
X"05337198",
X"2b71902b",
X"07963d33",
X"70882b72",
X"07029405",
X"80c70533",
X"71075152",
X"53575e5c",
X"74763178",
X"3179842a",
X"903d3354",
X"71713153",
X"5656b6ed",
X"3f83e080",
X"08820570",
X"881c0c83",
X"e08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83e0980c",
X"80567583",
X"e0800c97",
X"3d0d04e9",
X"3d0d83e0",
X"98085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e63f83e0",
X"80085483",
X"e0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f48a",
X"3f83e080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383e080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83e09808",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0e83f",
X"83e08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"843f83e0",
X"80085583",
X"e0800880",
X"2eff8938",
X"83e08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"51b4cf3f",
X"83e08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83e0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83e09808",
X"55568555",
X"73802e81",
X"e1388114",
X"33810653",
X"84557280",
X"2e81d338",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b7388214",
X"3370892b",
X"56537680",
X"2eb53874",
X"52ff1651",
X"b1ef3f83",
X"e08008ff",
X"18765470",
X"535853b1",
X"e03f83e0",
X"80087326",
X"96387430",
X"70780670",
X"98170c77",
X"7131a417",
X"08525851",
X"538939a0",
X"140870a4",
X"160c5374",
X"7627b938",
X"7251eed7",
X"3f83e080",
X"0853810b",
X"83e08008",
X"278b3888",
X"140883e0",
X"80082688",
X"38800b81",
X"1534b039",
X"83e08008",
X"a4150c98",
X"14081598",
X"150c7575",
X"3156c439",
X"98140816",
X"7098160c",
X"735256ef",
X"c83f83e0",
X"80088c38",
X"83e08008",
X"81153481",
X"55943982",
X"1433ff05",
X"76892a06",
X"83e08008",
X"05a8150c",
X"80557483",
X"e0800c88",
X"3d0d04ef",
X"3d0d6356",
X"855583e0",
X"9808802e",
X"80d23893",
X"3df40584",
X"170c6453",
X"883d7053",
X"765257f1",
X"d23f83e0",
X"80085583",
X"e08008b4",
X"38883d33",
X"5473802e",
X"a13802a7",
X"05337084",
X"2a708106",
X"51555583",
X"5573802e",
X"97387651",
X"eef83f83",
X"e0800888",
X"170c7551",
X"efa93f83",
X"e0800855",
X"7483e080",
X"0c933d0d",
X"04e43d0d",
X"6ea13d08",
X"405e8556",
X"83e09808",
X"802e8485",
X"389e3df4",
X"05841f0c",
X"7e98387d",
X"51eef83f",
X"83e08008",
X"5683ee39",
X"814181f6",
X"39834181",
X"f139933d",
X"7f960541",
X"59807f82",
X"95055e56",
X"756081ff",
X"05348341",
X"901e0876",
X"2e81d338",
X"a0547d22",
X"70852b83",
X"e0065458",
X"901e0852",
X"7851b0da",
X"3f83e080",
X"084183e0",
X"8008ffb8",
X"3878335c",
X"7b802eff",
X"b4388b19",
X"3370bf06",
X"71810652",
X"43557480",
X"2e80de38",
X"7b81bf06",
X"55748f24",
X"80d3389a",
X"19335574",
X"80cb38f3",
X"1d70585d",
X"8156758b",
X"2e098106",
X"85388e56",
X"8b39759a",
X"2e098106",
X"83389c56",
X"75197070",
X"81055233",
X"7133811a",
X"821a5f5b",
X"525b5574",
X"86387977",
X"34853980",
X"df773477",
X"7b57577a",
X"a02e0981",
X"06c03881",
X"567b81e5",
X"32703070",
X"9f2a5151",
X"557bae2e",
X"93387480",
X"2e8e3861",
X"832a7081",
X"06515574",
X"802e9738",
X"7d51ede2",
X"3f83e080",
X"084183e0",
X"80088738",
X"901e08fe",
X"af388060",
X"3475802e",
X"88387c52",
X"7f5183a5",
X"3f60802e",
X"8638800b",
X"901f0c60",
X"5660832e",
X"85386081",
X"d038891f",
X"57901e08",
X"802e81a8",
X"38805675",
X"19703351",
X"5574a02e",
X"a0387485",
X"2e098106",
X"843881e5",
X"55747770",
X"81055934",
X"81167081",
X"ff065755",
X"877627d7",
X"38881933",
X"5574a02e",
X"a938ae77",
X"70810559",
X"34885675",
X"19703351",
X"5574a02e",
X"95387477",
X"70810559",
X"34811670",
X"81ff0657",
X"558a7627",
X"e2388b19",
X"337f8805",
X"349f1933",
X"9e1a3371",
X"982b7190",
X"2b079d1c",
X"3370882b",
X"72079c1e",
X"33710764",
X"0c52991d",
X"33981e33",
X"71882b07",
X"53515357",
X"5956747f",
X"84052397",
X"1933961a",
X"3371882b",
X"07565674",
X"7f860523",
X"8077347d",
X"51ebf33f",
X"83e08008",
X"83327030",
X"7072079f",
X"2c83e080",
X"08065256",
X"56961f33",
X"55748a38",
X"891f5296",
X"1f5181b1",
X"3f7583e0",
X"800c9e3d",
X"0d04fd3d",
X"0d757753",
X"54733351",
X"70893871",
X"33517080",
X"2ea13873",
X"33723352",
X"53727127",
X"8538ff51",
X"94397073",
X"27853881",
X"518b3981",
X"14811353",
X"54d33980",
X"517083e0",
X"800c853d",
X"0d04fd3d",
X"0d757754",
X"54723370",
X"81ff0652",
X"5270802e",
X"a3387181",
X"ff068114",
X"ffbf1253",
X"54527099",
X"268938a0",
X"127081ff",
X"06535171",
X"74708105",
X"5634d239",
X"80743485",
X"3d0d04ff",
X"bd3d0d80",
X"c63d0852",
X"a53d7052",
X"54ffb33f",
X"80c73d08",
X"52853d70",
X"5253ffa6",
X"3f725273",
X"51fedf3f",
X"80c53d0d",
X"04fe3d0d",
X"74765353",
X"71708105",
X"53335170",
X"73708105",
X"553470f0",
X"38843d0d",
X"04fe3d0d",
X"74528072",
X"33525370",
X"732e8d38",
X"81128114",
X"71335354",
X"5270f538",
X"7283e080",
X"0c843d0d",
X"047183e3",
X"9c0c8880",
X"800b83e3",
X"980c8480",
X"800b83e3",
X"a00c04fd",
X"3d0d7770",
X"17557705",
X"ff1a5353",
X"71ff2e94",
X"38737081",
X"05553351",
X"70737081",
X"055534ff",
X"1252e939",
X"853d0d04",
X"fc3d0d87",
X"a6815574",
X"3383e3a4",
X"34a05483",
X"a0805383",
X"e39c0852",
X"83e39808",
X"51ffb83f",
X"a05483a4",
X"805383e3",
X"9c085283",
X"e3980851",
X"ffa53f90",
X"5483a880",
X"5383e39c",
X"085283e3",
X"980851ff",
X"923fa053",
X"805283e3",
X"a00883a0",
X"80055185",
X"b93fa053",
X"805283e3",
X"a00883a4",
X"80055185",
X"a93f9053",
X"805283e3",
X"a00883a8",
X"80055185",
X"993fff75",
X"3483a080",
X"54805383",
X"e39c0852",
X"83e3a008",
X"51fecc3f",
X"80d08054",
X"83b08053",
X"83e39c08",
X"5283e3a0",
X"0851feb7",
X"3f86cc3f",
X"a2548053",
X"83e3a008",
X"8c800552",
X"80efa051",
X"fea13f86",
X"0b87a883",
X"34800b87",
X"a8823480",
X"0b87a09a",
X"34af0b87",
X"a09634bf",
X"0b87a097",
X"34800b87",
X"a098349f",
X"0b87a099",
X"34800b87",
X"a09b34e0",
X"0b87a889",
X"34a20b87",
X"a8803483",
X"0b87a48f",
X"34820b87",
X"a8813486",
X"3d0d04fd",
X"3d0d83a0",
X"80548053",
X"83e3a008",
X"5283e39c",
X"0851fdbf",
X"3f80d080",
X"5483b080",
X"5383e3a0",
X"085283e3",
X"9c0851fd",
X"aa3fa054",
X"83a08053",
X"83e3a008",
X"5283e39c",
X"0851fd97",
X"3fa05483",
X"a4805383",
X"e3a00852",
X"83e39c08",
X"51fd843f",
X"905483a8",
X"805383e3",
X"a0085283",
X"e39c0851",
X"fcf13f83",
X"e3a43387",
X"a6813485",
X"3d0d0480",
X"3d0d9080",
X"90088106",
X"83e0800c",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fe0676",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70812c81",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870fd",
X"06761007",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"822cbf06",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fe83",
X"0676822b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70882c87",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870f1",
X"ff067688",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"08708b2c",
X"bf0683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"f88fff06",
X"768b2b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"912cbf06",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fc87",
X"ffff0676",
X"912b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087099",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70ffbf0a",
X"0676992b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90808008",
X"70882c81",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"0870892c",
X"810683e0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708a",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8b2c8106",
X"83e0800c",
X"51823d0d",
X"04fe3d0d",
X"7481e629",
X"872a9080",
X"a00c843d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"81055434",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727084",
X"05540cff",
X"1151f039",
X"843d0d04",
X"fe3d0d84",
X"80805380",
X"5288800a",
X"51ffb33f",
X"81808053",
X"80528280",
X"0a51c63f",
X"843d0d04",
X"803d0d81",
X"51fc913f",
X"72802e90",
X"388051fe",
X"933fcd3f",
X"83e3a833",
X"51fe893f",
X"8151fca2",
X"3f8051fc",
X"9d3f8051",
X"fbee3f82",
X"3d0d04fd",
X"3d0d7552",
X"805480ff",
X"72258838",
X"810bff80",
X"135354ff",
X"bf125170",
X"99268638",
X"e012529e",
X"39ff9f12",
X"51997127",
X"9538d012",
X"e0137054",
X"54518971",
X"2788388f",
X"73278338",
X"80527380",
X"2e853881",
X"80125271",
X"81ff0683",
X"e0800c85",
X"3d0d0480",
X"3d0d84d8",
X"c0518071",
X"70810553",
X"347084e0",
X"c02e0981",
X"06f03882",
X"3d0d04fe",
X"3d0d0297",
X"053351ff",
X"863f83e0",
X"800881ff",
X"0683e3ac",
X"08545280",
X"73249b38",
X"83e3cc08",
X"137283e3",
X"d0080753",
X"53717334",
X"83e3ac08",
X"810583e3",
X"ac0c843d",
X"0d04fa3d",
X"0d82800a",
X"1b558057",
X"883dfc05",
X"54795374",
X"527851d5",
X"e33f883d",
X"0d04fe3d",
X"0d83e3c4",
X"08527451",
X"dcc83f83",
X"e080088c",
X"38765375",
X"5283e3c4",
X"0851c73f",
X"843d0d04",
X"fe3d0d83",
X"e3c40853",
X"75527451",
X"d7863f83",
X"e080088d",
X"38775376",
X"5283e3c4",
X"0851ffa2",
X"3f843d0d",
X"04fe3d0d",
X"83e3c408",
X"51d5fa3f",
X"83e08008",
X"8180802e",
X"09810688",
X"3883c180",
X"80539b39",
X"83e3c408",
X"51d5de3f",
X"83e08008",
X"80d0802e",
X"09810693",
X"3883c1b0",
X"805383e0",
X"80085283",
X"e3c40851",
X"fed83f84",
X"3d0d0480",
X"3d0df9f9",
X"3f83e080",
X"08842980",
X"efc40570",
X"0883e080",
X"0c51823d",
X"0d04ee3d",
X"0d804380",
X"42804180",
X"705a5bfd",
X"d23f800b",
X"83e3ac0c",
X"800b83e3",
X"d00c80ed",
X"9451d0c8",
X"3f81800b",
X"83e3d00c",
X"80ed9851",
X"d0ba3f80",
X"d00b83e3",
X"ac0c7830",
X"707a0780",
X"2570872b",
X"83e3d00c",
X"5155f8ec",
X"3f83e080",
X"085280ed",
X"a051d094",
X"3f80f80b",
X"83e3ac0c",
X"78813270",
X"30707207",
X"80257087",
X"2b83e3d0",
X"0c515656",
X"fef13f83",
X"e0800852",
X"80edac51",
X"cfea3f81",
X"a00b83e3",
X"ac0c7882",
X"32703070",
X"72078025",
X"70872b83",
X"e3d00c51",
X"5683e3c4",
X"085256d1",
X"843f83e0",
X"80085280",
X"edb451cf",
X"bb3f81f0",
X"0b83e3ac",
X"0c810b83",
X"e3b05b58",
X"83e3ac08",
X"82197a32",
X"70307072",
X"07802570",
X"872b83e3",
X"d00c5157",
X"8e3d7055",
X"ff1b5457",
X"575799f9",
X"3f797084",
X"055b0851",
X"d0bb3f74",
X"5483e080",
X"08537752",
X"80edbc51",
X"ceee3fa8",
X"1783e3ac",
X"0c811858",
X"77852e09",
X"8106ffb0",
X"3883900b",
X"83e3ac0c",
X"78873270",
X"30707207",
X"80257087",
X"2b83e3d0",
X"0c515656",
X"f8923f80",
X"edcc5583",
X"e0800880",
X"2e8e3883",
X"e3c00851",
X"cfe73f83",
X"e0800855",
X"745280ed",
X"d451ce9c",
X"3f83e00b",
X"83e3ac0c",
X"78883270",
X"30707207",
X"80257087",
X"2b83e3d0",
X"0c515780",
X"ede05255",
X"cdfa3f86",
X"8da051f8",
X"f83f8052",
X"913d7052",
X"559acb3f",
X"83527451",
X"9ac43f61",
X"19597880",
X"25853880",
X"59903988",
X"79258538",
X"88598739",
X"78882682",
X"db387882",
X"2b5580eb",
X"f0150804",
X"f6863f83",
X"e0800861",
X"57557581",
X"2e098106",
X"893883e0",
X"80081055",
X"903975ff",
X"2e098106",
X"883883e0",
X"8008812c",
X"55907525",
X"85389055",
X"88397480",
X"24833881",
X"557451f5",
X"e03f8290",
X"39f5f23f",
X"83e08008",
X"61055574",
X"80258538",
X"80558839",
X"87752583",
X"38875574",
X"51f5eb3f",
X"81ee3960",
X"87386280",
X"2e81e538",
X"83e0a408",
X"83e0a00c",
X"8bdf0b83",
X"e0a80c83",
X"e3c40851",
X"ffbf9a3f",
X"fae73f81",
X"c7396056",
X"80762599",
X"388af80b",
X"83e0a80c",
X"83e3a415",
X"70085255",
X"ffbefa3f",
X"74085291",
X"39758025",
X"913883e3",
X"a4150851",
X"cdd53f80",
X"52fd1951",
X"b8396280",
X"2e818d38",
X"83e3a415",
X"700883e3",
X"b008720c",
X"83e3b00c",
X"fd1a7053",
X"51558be9",
X"3f83e080",
X"08568051",
X"8bdf3f83",
X"e0800852",
X"745187fd",
X"3f755280",
X"5187f63f",
X"80d63960",
X"55807525",
X"b83883e0",
X"ac0883e0",
X"a00c8bdf",
X"0b83e0a8",
X"0c83e3c0",
X"0851ffbe",
X"843f83e3",
X"c00851ff",
X"bb9e3f83",
X"e0800881",
X"ff067052",
X"55f4f63f",
X"74802e9c",
X"388155a0",
X"39748025",
X"933883e3",
X"c00851cc",
X"c63f8051",
X"f4db3f84",
X"39628738",
X"7a802efa",
X"8a388055",
X"7483e080",
X"0c943d0d",
X"04fe3d0d",
X"f5873f83",
X"e0800880",
X"2e863880",
X"51818b39",
X"f58c3f83",
X"e0800880",
X"ff38f5ac",
X"3f83e080",
X"08802eb9",
X"388151f2",
X"bb3f8051",
X"f4c23fef",
X"af3f800b",
X"83e3ac0c",
X"f9b43f83",
X"e0800853",
X"ff0b83e3",
X"ac0cf19b",
X"3f7280cc",
X"3883e3a8",
X"3351f49c",
X"3f7251f2",
X"8b3f80c1",
X"39f4d43f",
X"83e08008",
X"802eb638",
X"8151f1f8",
X"3f8051f3",
X"ff3feeec",
X"3f8af80b",
X"83e0a80c",
X"83e3b008",
X"51ffbcb5",
X"3fff0b83",
X"e3ac0cf0",
X"d63f83e3",
X"b0085280",
X"5185f23f",
X"8151f5b0",
X"3f843d0d",
X"04fb3d0d",
X"800b83e3",
X"a8349080",
X"80528684",
X"808051cf",
X"813f83e0",
X"80088193",
X"3889b73f",
X"80f19851",
X"d3c23f83",
X"e0800855",
X"9c800a54",
X"80c08053",
X"80ede852",
X"83e08008",
X"51f7853f",
X"83e3c408",
X"5380edf8",
X"527451ce",
X"8b3f83e0",
X"80088438",
X"f7933f83",
X"e3c80853",
X"80ee8452",
X"7451cdf4",
X"3f83e080",
X"08b53887",
X"3dfc0554",
X"84808053",
X"86a88080",
X"5283e3c8",
X"0851cc80",
X"3f83e080",
X"08933875",
X"8480802e",
X"09810689",
X"38810b83",
X"e3a83487",
X"39800b83",
X"e3a83483",
X"e3a83351",
X"f2aa3f81",
X"51f4813f",
X"92f33f81",
X"51f3f93f",
X"fda73ffc",
X"3983e08c",
X"080283e0",
X"8c0cfb3d",
X"0d0280ee",
X"900b83e0",
X"a40c80ee",
X"940b83e0",
X"9c0c80ee",
X"980b83e0",
X"ac0c83e0",
X"8c08fc05",
X"0c800b83",
X"e3b00b83",
X"e08c08f8",
X"050c83e0",
X"8c08f405",
X"0ccc933f",
X"83e08008",
X"8605fc06",
X"83e08c08",
X"f0050c02",
X"83e08c08",
X"f0050831",
X"0d833d70",
X"83e08c08",
X"f8050870",
X"840583e0",
X"8c08f805",
X"0c0c51c8",
X"da3f83e0",
X"8c08f405",
X"08810583",
X"e08c08f4",
X"050c83e0",
X"8c08f405",
X"08872e09",
X"8106ffad",
X"38869480",
X"8051ebad",
X"3fff0b83",
X"e3ac0c80",
X"0b83e3d0",
X"0c84d8c0",
X"0b83e3cc",
X"0c8151ee",
X"d73f8151",
X"eefc3f80",
X"51eef73f",
X"8151ef9d",
X"3f8151ef",
X"f23f8251",
X"efc03f80",
X"51f0963f",
X"8051f0c0",
X"3f80c6c3",
X"528051c6",
X"943ffce5",
X"3f83e08c",
X"08fc0508",
X"0d800b83",
X"e0800c87",
X"3d0d83e0",
X"8c0c0480",
X"3d0d81ff",
X"51800b83",
X"e3dc1234",
X"ff115170",
X"f438823d",
X"0d04ff3d",
X"0d737033",
X"53518111",
X"33713471",
X"81123483",
X"3d0d04fb",
X"3d0d7779",
X"56568070",
X"71555552",
X"717525ac",
X"38721670",
X"33701470",
X"81ff0655",
X"51515171",
X"74278938",
X"81127081",
X"ff065351",
X"71811470",
X"83ffff06",
X"55525474",
X"7324d638",
X"7183e080",
X"0c873d0d",
X"04fc3d0d",
X"7655ffbf",
X"c03f83e0",
X"8008802e",
X"f53883e5",
X"f8088605",
X"7081ff06",
X"5253ffbd",
X"c13f8439",
X"fa933fff",
X"bf9f3f83",
X"e0800881",
X"2ef23880",
X"54731553",
X"ffbe863f",
X"83e08008",
X"73348114",
X"5473852e",
X"098106e9",
X"388439f9",
X"e83fffbe",
X"f43f83e0",
X"8008802e",
X"f2387433",
X"83e3dc34",
X"81153383",
X"e3dd3482",
X"153383e3",
X"de348315",
X"3383e3df",
X"34845283",
X"e3dc51fe",
X"ba3f83e0",
X"800881ff",
X"06841633",
X"56537275",
X"2e098106",
X"8d38ffbd",
X"e93f83e0",
X"8008802e",
X"9a3883e5",
X"f808a82e",
X"09810689",
X"38860b83",
X"e5f80c87",
X"39a80b83",
X"e5f80c80",
X"e451eed9",
X"3f863d0d",
X"04f43d0d",
X"7e605955",
X"805d8075",
X"822b7183",
X"e5fc120c",
X"83e69017",
X"5b5b5776",
X"79347777",
X"2e83b238",
X"76527751",
X"c7a23f8e",
X"3dfc0554",
X"905383e5",
X"e4527751",
X"c6de3f7c",
X"5675902e",
X"09810683",
X"903883e5",
X"e451fd96",
X"3f83e5e6",
X"51fd8f3f",
X"83e5e851",
X"fd883f76",
X"83e5f40c",
X"7751c4a9",
X"3f80eca4",
X"5283e080",
X"0851ffb3",
X"e53f83e0",
X"8008812e",
X"09810680",
X"d3387683",
X"e68c0c82",
X"0b83e5e4",
X"34ff960b",
X"83e5e534",
X"7751c6f1",
X"3f83e080",
X"085583e0",
X"80087725",
X"883883e0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83e5e634",
X"7483e5e7",
X"347683e5",
X"e834ff80",
X"0b83e5e9",
X"34818f39",
X"83e5e433",
X"83e5e533",
X"71882b07",
X"565b7483",
X"ffff2e09",
X"810680e7",
X"38fe800b",
X"83e68c0c",
X"810b83e5",
X"f40cff0b",
X"83e5e434",
X"ff0b83e5",
X"e5347751",
X"c5ff3f83",
X"e0800883",
X"e6940c83",
X"e0800855",
X"83e08008",
X"80258838",
X"83e08008",
X"8f055574",
X"842c7083",
X"ffff0670",
X"882a5851",
X"557583e5",
X"e6347483",
X"e5e73476",
X"83e5e834",
X"ff800b83",
X"e5e93481",
X"0b83e5f3",
X"34a43974",
X"85962e09",
X"810680fd",
X"387583e6",
X"8c0c7751",
X"c5b43f83",
X"e5f33383",
X"e0800807",
X"557483e5",
X"f33483e5",
X"f3338106",
X"5574802e",
X"83388457",
X"83e5e833",
X"83e5e933",
X"71882b07",
X"565c7481",
X"802e0981",
X"06a13883",
X"e5e63383",
X"e5e73371",
X"882b0756",
X"5bad8075",
X"27873876",
X"8207579c",
X"39768107",
X"57963974",
X"82802e09",
X"81068738",
X"76830757",
X"87397481",
X"ff268a38",
X"7783e5fc",
X"1b0c7679",
X"348e3d0d",
X"04803d0d",
X"72842983",
X"e5fc0570",
X"0883e080",
X"0c51823d",
X"0d04fe3d",
X"0d800b83",
X"e5e00c80",
X"0b83e5dc",
X"0cff0b83",
X"e3d80ca8",
X"0b83e5f8",
X"0cae51ff",
X"b8903f80",
X"0b83e5fc",
X"54528073",
X"70840555",
X"0c811252",
X"71842e09",
X"8106ef38",
X"843d0d04",
X"fe3d0d74",
X"02840596",
X"05225353",
X"71802e97",
X"38727081",
X"05543351",
X"ffb89a3f",
X"ff127083",
X"ffff0651",
X"52e63984",
X"3d0d04fe",
X"3d0d0292",
X"05225382",
X"ac51e9f1",
X"3f80c351",
X"ffb7f63f",
X"819651e9",
X"e43f7252",
X"83e3dc51",
X"ffb23f72",
X"5283e3dc",
X"51f8f43f",
X"83e08008",
X"81ff0651",
X"ffb7d23f",
X"843d0d04",
X"ffb13d0d",
X"80d13df8",
X"0551f99d",
X"3f83e5e0",
X"08810583",
X"e5e00c80",
X"cf3d33cf",
X"117081ff",
X"06515656",
X"74832688",
X"ed38758f",
X"06ff0556",
X"7583e3d8",
X"082e9b38",
X"75832696",
X"387583e3",
X"d80c7584",
X"2983e5fc",
X"05700853",
X"557551fa",
X"9c3f8076",
X"2488c938",
X"75842983",
X"e5fc0555",
X"7408802e",
X"88ba3883",
X"e3d80884",
X"2983e5fc",
X"05700802",
X"880582b9",
X"0533525b",
X"557480d2",
X"2e84b138",
X"7480d224",
X"903874bf",
X"2e9c3874",
X"80d02e81",
X"d73887f8",
X"397480d3",
X"2e80d238",
X"7480d72e",
X"81c63887",
X"e7390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290556",
X"56ffb6cd",
X"3f80c151",
X"ffb6863f",
X"f6ed3f86",
X"0b83e3dc",
X"34815283",
X"e3dc51ff",
X"b7a83f81",
X"51fde43f",
X"74893886",
X"0b83e5f8",
X"0c8739a8",
X"0b83e5f8",
X"0cffb699",
X"3f80c151",
X"ffb5d23f",
X"f6b93f90",
X"0b83e5f3",
X"33810656",
X"5674802e",
X"83389856",
X"83e5e833",
X"83e5e933",
X"71882b07",
X"56597481",
X"802e0981",
X"069c3883",
X"e5e63383",
X"e5e73371",
X"882b0756",
X"57ad8075",
X"278c3875",
X"81800756",
X"853975a0",
X"07567583",
X"e3dc34ff",
X"0b83e3dd",
X"34e00b83",
X"e3de3480",
X"0b83e3df",
X"34845283",
X"e3dc51ff",
X"b69c3f84",
X"51869e39",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"055659ff",
X"b58b3f79",
X"51ffbffa",
X"3f83e080",
X"08802e8b",
X"3880ce51",
X"ffb4b63f",
X"85f23980",
X"c151ffb4",
X"ac3fffb5",
X"a03fffb3",
X"d43f83e6",
X"8c085883",
X"75259b38",
X"83e5e833",
X"83e5e933",
X"71882b07",
X"fc177129",
X"7a058380",
X"055a5157",
X"8d397481",
X"802918ff",
X"80055881",
X"80578056",
X"76762e93",
X"38ffb485",
X"3f83e080",
X"0883e3dc",
X"17348116",
X"56ea39ff",
X"b3f33f83",
X"e0800881",
X"ff067753",
X"83e3dc52",
X"56f4dc3f",
X"83e08008",
X"81ff0655",
X"75752e09",
X"8106818a",
X"38ffb3f1",
X"3f80c151",
X"ffb3aa3f",
X"ffb49e3f",
X"77527951",
X"ffbe893f",
X"805e80d1",
X"3dfdf405",
X"54765383",
X"e3dc5279",
X"51ffbc95",
X"3f0282b9",
X"05335581",
X"587480d7",
X"2e098106",
X"bd3880d1",
X"3dfdf005",
X"5476538f",
X"3d70537a",
X"5259ffbd",
X"9b3f8056",
X"76762ea2",
X"38751983",
X"e3dc1733",
X"71337072",
X"32703070",
X"80257030",
X"7e06811d",
X"5d5e5151",
X"51525b55",
X"db3982ac",
X"51e4aa3f",
X"77802e86",
X"3880c351",
X"843980ce",
X"51ffb2a5",
X"3fffb399",
X"3fffb1cd",
X"3f83dd39",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"05595580",
X"705d59ff",
X"b2bf3f80",
X"c151ffb1",
X"f83f83e5",
X"f408792e",
X"82de3883",
X"e6940880",
X"fc055580",
X"fd527451",
X"86d73f83",
X"e080085b",
X"778224b2",
X"38ff1870",
X"872b83ff",
X"ff800680",
X"efe40583",
X"e3dc5957",
X"55818055",
X"75708105",
X"57337770",
X"81055934",
X"ff157081",
X"ff065155",
X"74ea3882",
X"8d397782",
X"e82e81ab",
X"387782e9",
X"2e098106",
X"81b23880",
X"ee9c51ff",
X"b7fa3f78",
X"58778732",
X"70307072",
X"0780257a",
X"8a327030",
X"70720780",
X"25730753",
X"545a5157",
X"5575802e",
X"97387878",
X"269238a0",
X"0b83e3dc",
X"1a348119",
X"7081ff06",
X"5a55eb39",
X"81187081",
X"ff065955",
X"8a7827ff",
X"bc388f58",
X"83e3d718",
X"3383e3dc",
X"1934ff18",
X"7081ff06",
X"59557784",
X"26ea3890",
X"58800b83",
X"e3dc1934",
X"81187081",
X"ff067098",
X"2b525955",
X"748025e9",
X"3880c655",
X"7a858f24",
X"843880c2",
X"557483e3",
X"dc3480f1",
X"0b83e3df",
X"34810b83",
X"e3e0347a",
X"83e3dd34",
X"7a882c55",
X"7483e3de",
X"3480cb39",
X"82f07825",
X"80c43877",
X"80fd29fd",
X"97d30552",
X"7951ffba",
X"b73f80d1",
X"3dfdec05",
X"5480fd53",
X"83e3dc52",
X"7951ffb9",
X"ef3f7b81",
X"19595675",
X"80fc2483",
X"38785877",
X"882c5574",
X"83e4d934",
X"7783e4da",
X"347583e4",
X"db348180",
X"5980cc39",
X"83e68c08",
X"57837825",
X"9b3883e5",
X"e83383e5",
X"e9337188",
X"2b07fc1a",
X"71297905",
X"83800559",
X"51598d39",
X"77818029",
X"17ff8005",
X"57818059",
X"76527951",
X"ffb9c53f",
X"80d13dfd",
X"ec055478",
X"5383e3dc",
X"527951ff",
X"b8fe3f78",
X"51f6b83f",
X"ffafb63f",
X"ffadea3f",
X"8b3983e5",
X"dc088105",
X"83e5dc0c",
X"80d13d0d",
X"04f6d93f",
X"eab73ff9",
X"39fc3d0d",
X"76787184",
X"2983e5fc",
X"05700851",
X"53535370",
X"9e3880ce",
X"723480cf",
X"0b811334",
X"80ce0b82",
X"133480c5",
X"0b831334",
X"70841334",
X"80e73983",
X"e6901333",
X"5480d272",
X"3473822a",
X"70810651",
X"5180cf53",
X"70843880",
X"d7537281",
X"1334a00b",
X"82133473",
X"83065170",
X"812e9e38",
X"70812488",
X"3870802e",
X"8f389f39",
X"70822e92",
X"3870832e",
X"92389339",
X"80d8558e",
X"3980d355",
X"893980cd",
X"55843980",
X"c4557483",
X"133480c4",
X"0b841334",
X"800b8513",
X"34863d0d",
X"04fd3d0d",
X"75538073",
X"0c800b84",
X"140c800b",
X"88140c87",
X"a6803370",
X"81ff0670",
X"812a8132",
X"71813271",
X"81067181",
X"06318418",
X"0c555670",
X"832a8132",
X"71822a81",
X"32718106",
X"71810631",
X"770c5254",
X"515187a0",
X"90337009",
X"81068815",
X"0c51853d",
X"0d04fe3d",
X"0d747654",
X"527151ff",
X"a03f7281",
X"2ea23881",
X"73268d38",
X"72822eab",
X"3872832e",
X"9f38e639",
X"7108e238",
X"841208dd",
X"38881208",
X"d838a039",
X"88120881",
X"2e098106",
X"cc389439",
X"88120881",
X"2e8d3871",
X"08893884",
X"1208802e",
X"ffb73884",
X"3d0d04fc",
X"3d0d7678",
X"53548153",
X"80558739",
X"71107310",
X"54527372",
X"26517280",
X"2ea73870",
X"802e8638",
X"718025e8",
X"3872802e",
X"98387174",
X"26893873",
X"72317574",
X"07565472",
X"812a7281",
X"2a5353e5",
X"39735178",
X"83387451",
X"7083e080",
X"0c863d0d",
X"04fe3d0d",
X"80537552",
X"7451ffa3",
X"3f843d0d",
X"04fe3d0d",
X"81537552",
X"7451ff93",
X"3f843d0d",
X"04fb3d0d",
X"77795555",
X"80567476",
X"25863874",
X"30558156",
X"73802588",
X"38733076",
X"81325754",
X"80537352",
X"7451fee7",
X"3f83e080",
X"08547580",
X"2e873883",
X"e0800830",
X"547383e0",
X"800c873d",
X"0d04fa3d",
X"0d787a57",
X"55805774",
X"77258638",
X"74305581",
X"57759f2c",
X"54815375",
X"74327431",
X"527451fe",
X"aa3f83e0",
X"80085476",
X"802e8738",
X"83e08008",
X"30547383",
X"e0800c88",
X"3d0d04ff",
X"3d0d7352",
X"7183e69c",
X"082ea638",
X"71a00a07",
X"90809c0c",
X"90808c08",
X"5170802e",
X"f738800b",
X"90809c0c",
X"90808c08",
X"5170f938",
X"7183e69c",
X"0c833d0d",
X"04ff0b83",
X"e69c0c81",
X"80800b83",
X"e6980c80",
X"0b83e080",
X"0c04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"9e3f7280",
X"2ea33883",
X"e6980814",
X"52713375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552da",
X"39800b83",
X"e0800c86",
X"3d0d04f7",
X"3d0d7b7d",
X"7f115855",
X"59805573",
X"762eb138",
X"83e69808",
X"8b3d5957",
X"74197033",
X"75fc0619",
X"70085d76",
X"83067b07",
X"53545451",
X"72713479",
X"720c8114",
X"81165654",
X"73762e09",
X"8106d938",
X"800b83e0",
X"800c8b3d",
X"0d04803d",
X"0d83e69c",
X"08900a07",
X"90809c0c",
X"90808c08",
X"5170802e",
X"f738800b",
X"90809c0c",
X"90808c08",
X"5170f938",
X"823d0d04",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"000025f4",
X"00002635",
X"00002657",
X"0000267e",
X"0000267e",
X"0000267e",
X"0000267e",
X"000026ef",
X"00002741",
X"25732025",
X"73000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"66726565",
X"7a65722e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"6e616d65",
X"20000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00003650",
X"00003654",
X"0000365c",
X"00003668",
X"00003674",
X"00003680",
X"0000368c",
X"00003690",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
