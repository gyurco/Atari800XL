
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f5",
X"b4738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80f9",
X"c80c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f2",
X"e22d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580f2a1",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80dcb004",
X"fd3d0d75",
X"705254ae",
X"ab3f83e0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83e0",
X"8008732e",
X"a13883e0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183e0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83e2c008",
X"248a38b4",
X"fc3fff0b",
X"83e2c00c",
X"800b83e0",
X"800c04ff",
X"3d0d7352",
X"83e09c08",
X"722e8d38",
X"d93f7151",
X"96a03f71",
X"83e09c0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"55805681",
X"54bc1508",
X"762e0981",
X"06819138",
X"7451c83f",
X"7958757a",
X"2580f738",
X"83e2f008",
X"70892a57",
X"83ff0678",
X"84807231",
X"56565773",
X"78258338",
X"73557583",
X"e2c0082e",
X"8438ff82",
X"3f83e2c0",
X"088025a6",
X"3875892b",
X"5198dc3f",
X"83e2f008",
X"8f3dfc11",
X"555c5481",
X"52f81b51",
X"96c63f76",
X"1483e2f0",
X"0c7583e2",
X"c00c7453",
X"76527851",
X"b3a63f83",
X"e0800883",
X"e2f00816",
X"83e2f00c",
X"78763176",
X"1b5b5956",
X"778024ff",
X"8b38617a",
X"710c5475",
X"5475802e",
X"83388154",
X"7383e080",
X"0c8e3d0d",
X"04fc3d0d",
X"fe943f76",
X"51fea83f",
X"863dfc05",
X"53785277",
X"5195e93f",
X"7975710c",
X"5483e080",
X"085483e0",
X"8008802e",
X"83388154",
X"7383e080",
X"0c863d0d",
X"04fe3d0d",
X"7583e2c0",
X"08535380",
X"72248938",
X"71732e84",
X"38fdcf3f",
X"7451fde3",
X"3f725197",
X"ae3f83e0",
X"80085283",
X"e0800880",
X"2e833881",
X"527183e0",
X"800c843d",
X"0d04803d",
X"0d7280c0",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d72bc",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"c40b83e0",
X"800c04fd",
X"3d0d7577",
X"71547053",
X"5553a9fc",
X"3f82c813",
X"08bc150c",
X"82c01308",
X"80c0150c",
X"fce43f73",
X"5193ab3f",
X"7383e09c",
X"0c83e080",
X"085383e0",
X"8008802e",
X"83388153",
X"7283e080",
X"0c853d0d",
X"04fd3d0d",
X"75775553",
X"fcb83f72",
X"802ea538",
X"bc130852",
X"7351a986",
X"3f83e080",
X"088f3877",
X"527251ff",
X"9a3f83e0",
X"8008538a",
X"3982cc13",
X"0853d839",
X"81537283",
X"e0800c85",
X"3d0d04fe",
X"3d0dff0b",
X"83e2c00c",
X"7483e0a0",
X"0c7583e2",
X"bc0cafda",
X"3f83e080",
X"0881ff06",
X"52815371",
X"993883e2",
X"d8518e94",
X"3f83e080",
X"085283e0",
X"8008802e",
X"83387252",
X"71537283",
X"e0800c84",
X"3d0d04fa",
X"3d0d787a",
X"82c41208",
X"82c41208",
X"70722459",
X"56565757",
X"73732e09",
X"81069138",
X"80c01652",
X"80c01751",
X"a6f73f83",
X"e0800855",
X"7483e080",
X"0c883d0d",
X"04f63d0d",
X"7c5b807b",
X"715c5457",
X"7a772e8c",
X"38811a82",
X"cc140854",
X"5a72f638",
X"805980d9",
X"397a5481",
X"5780707b",
X"7b315a57",
X"55ff1853",
X"74732580",
X"c13882cc",
X"14085273",
X"51ff8c3f",
X"800b83e0",
X"800825a1",
X"3882cc14",
X"0882cc11",
X"0882cc16",
X"0c7482cc",
X"120c5375",
X"802e8638",
X"7282cc17",
X"0c725480",
X"577382cc",
X"15088117",
X"575556ff",
X"b8398119",
X"59800bff",
X"1b545478",
X"73258338",
X"81547681",
X"32707506",
X"515372ff",
X"90388c3d",
X"0d04f73d",
X"0d7b7d5a",
X"5a82d052",
X"83e2bc08",
X"5180e19d",
X"3f83e080",
X"0857f9da",
X"3f795283",
X"e2c45195",
X"b73f83e0",
X"80085480",
X"5383e080",
X"08732e09",
X"81068283",
X"3883e0a0",
X"080b0b80",
X"f6ec5370",
X"5256a6b4",
X"3f0b0b80",
X"f6ec5280",
X"c01651a6",
X"a73f75bc",
X"170c7382",
X"c0170c81",
X"0b82c417",
X"0c810b82",
X"c8170c73",
X"82cc170c",
X"ff1782d0",
X"17555781",
X"913983e0",
X"ac337082",
X"2a708106",
X"51545572",
X"81803874",
X"812a8106",
X"587780f6",
X"3874842a",
X"810682c4",
X"150c83e0",
X"ac338106",
X"82c8150c",
X"79527351",
X"a5ce3f73",
X"51a5e53f",
X"83e08008",
X"1453af73",
X"70810555",
X"3472bc15",
X"0c83e0ad",
X"527251a5",
X"af3f83e0",
X"a40882c0",
X"150c83e0",
X"ba5280c0",
X"1451a59c",
X"3f78802e",
X"8d387351",
X"782d83e0",
X"8008802e",
X"99387782",
X"cc150c75",
X"802e8638",
X"7382cc17",
X"0c7382d0",
X"15ff1959",
X"55567680",
X"2e9b3883",
X"e0a45283",
X"e2c45194",
X"ad3f83e0",
X"80088a38",
X"83e0ad33",
X"5372fed2",
X"3878802e",
X"893883e0",
X"a00851fc",
X"b83f83e0",
X"a0085372",
X"83e0800c",
X"8b3d0d04",
X"ff3d0d80",
X"527351fd",
X"b53f833d",
X"0d04f03d",
X"0d627052",
X"54f6893f",
X"83e08008",
X"7453873d",
X"70535555",
X"f6a93ff7",
X"893f7351",
X"d33f6353",
X"745283e0",
X"800851fa",
X"b83f923d",
X"0d047183",
X"e0800c04",
X"80c01283",
X"e0800c04",
X"803d0d72",
X"82c01108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"7282cc11",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282c4",
X"110883e0",
X"800c5182",
X"3d0d04f9",
X"3d0d7983",
X"e0900857",
X"57817727",
X"81963876",
X"88170827",
X"818e3875",
X"33557482",
X"2e893874",
X"832eb338",
X"80fe3974",
X"54761083",
X"fe065376",
X"882a8c17",
X"08055289",
X"3dfc0551",
X"aa883f83",
X"e0800880",
X"df38029d",
X"0533893d",
X"3371882b",
X"07565680",
X"d1398454",
X"76822b83",
X"fc065376",
X"872a8c17",
X"08055289",
X"3dfc0551",
X"a9d83f83",
X"e08008b0",
X"38029f05",
X"33028405",
X"9e053371",
X"982b7190",
X"2b07028c",
X"059d0533",
X"70882b72",
X"078d3d33",
X"7180ffff",
X"fe800607",
X"51525357",
X"58568339",
X"81557483",
X"e0800c89",
X"3d0d04fb",
X"3d0d83e0",
X"9008fe19",
X"881208fe",
X"05555654",
X"80567473",
X"278d3882",
X"14337571",
X"29941608",
X"05575375",
X"83e0800c",
X"873d0d04",
X"fc3d0d76",
X"52800b83",
X"e0900870",
X"33515253",
X"70832e09",
X"81069138",
X"95123394",
X"13337198",
X"2b71902b",
X"07555551",
X"9b12339a",
X"13337188",
X"2b077407",
X"83e0800c",
X"55863d0d",
X"04fc3d0d",
X"7683e090",
X"08555580",
X"75238815",
X"08537281",
X"2e883888",
X"14087326",
X"85388152",
X"b2397290",
X"38733352",
X"71832e09",
X"81068538",
X"90140853",
X"728c160c",
X"72802e8d",
X"387251fe",
X"d63f83e0",
X"80085285",
X"39901408",
X"52719016",
X"0c805271",
X"83e0800c",
X"863d0d04",
X"fa3d0d78",
X"83e09008",
X"71228105",
X"7083ffff",
X"06575457",
X"5573802e",
X"88389015",
X"08537286",
X"38835280",
X"e739738f",
X"06527180",
X"da388113",
X"90160c8c",
X"15085372",
X"9038830b",
X"84172257",
X"52737627",
X"80c638bf",
X"39821633",
X"ff057484",
X"2a065271",
X"b2387251",
X"fcb13f81",
X"527183e0",
X"800827a8",
X"38835283",
X"e0800888",
X"1708279c",
X"3883e080",
X"088c160c",
X"83e08008",
X"51fdbc3f",
X"83e08008",
X"90160c73",
X"75238052",
X"7183e080",
X"0c883d0d",
X"04f23d0d",
X"60626458",
X"5e5b7533",
X"5574a02e",
X"09810688",
X"38811670",
X"4456ef39",
X"62703356",
X"5674af2e",
X"09810684",
X"38811643",
X"800b881c",
X"0c627033",
X"5155749f",
X"2691387a",
X"51fdd23f",
X"83e08008",
X"56807d34",
X"83813993",
X"3d841c08",
X"7058595f",
X"8a55a076",
X"70810558",
X"34ff1555",
X"74ff2e09",
X"8106ef38",
X"80705a5c",
X"887f085f",
X"5a7b811d",
X"7081ff06",
X"60137033",
X"70af3270",
X"30a07327",
X"71802507",
X"5151525b",
X"535e5755",
X"7480e738",
X"76ae2e09",
X"81068338",
X"8155787a",
X"27750755",
X"74802e9f",
X"38798832",
X"703078ae",
X"32703070",
X"73079f2a",
X"53515751",
X"5675bb38",
X"88598b5a",
X"ffab3976",
X"982b5574",
X"80258738",
X"80f4c417",
X"3357ff9f",
X"17557499",
X"268938e0",
X"177081ff",
X"06585578",
X"811a7081",
X"ff06721b",
X"535b5755",
X"767534fe",
X"f8397b1e",
X"7f0c8055",
X"76a02683",
X"38815574",
X"8b19347a",
X"51fc823f",
X"83e08008",
X"80f538a0",
X"547a2270",
X"852b83e0",
X"06545590",
X"1b08527c",
X"51a4933f",
X"83e08008",
X"5783e080",
X"08818138",
X"7c335574",
X"802e80f4",
X"388b1d33",
X"70832a70",
X"81065156",
X"5674b438",
X"8b7d841d",
X"0883e080",
X"08595b5b",
X"58ff1858",
X"77ff2e9a",
X"38797081",
X"055b3379",
X"7081055b",
X"33717131",
X"52565675",
X"802ee238",
X"86397580",
X"2e96387a",
X"51fbe53f",
X"ff863983",
X"e0800856",
X"83e08008",
X"b6388339",
X"7656841b",
X"088b1133",
X"515574a7",
X"388b1d33",
X"70842a70",
X"81065156",
X"56748938",
X"83569439",
X"81569039",
X"7c51fa94",
X"3f83e080",
X"08881c0c",
X"fd813975",
X"83e0800c",
X"903d0d04",
X"f83d0d7a",
X"7c595782",
X"5483fe53",
X"77527651",
X"a2d83f83",
X"5683e080",
X"0880ec38",
X"81173377",
X"3371882b",
X"07565682",
X"567482d4",
X"d52e0981",
X"0680d438",
X"7554b653",
X"77527651",
X"a2ac3f83",
X"e0800898",
X"38811733",
X"77337188",
X"2b0783e0",
X"80085256",
X"56748182",
X"c62eac38",
X"825480d2",
X"53775276",
X"51a2833f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62e83",
X"38815675",
X"83e0800c",
X"8a3d0d04",
X"eb3d0d67",
X"5a800b83",
X"e0900ca1",
X"a53f83e0",
X"80088106",
X"55825674",
X"83ef3874",
X"75538f3d",
X"70535759",
X"feca3f83",
X"e0800881",
X"ff065776",
X"812e0981",
X"0680d438",
X"905483be",
X"53745275",
X"51a1973f",
X"83e08008",
X"80c9388f",
X"3d335574",
X"802e80c9",
X"3802bf05",
X"33028405",
X"be053371",
X"982b7190",
X"2b07028c",
X"05bd0533",
X"70882b72",
X"07953d33",
X"71077058",
X"7b575e52",
X"5e575957",
X"fdee3f83",
X"e0800881",
X"ff065776",
X"832e0981",
X"06863881",
X"5682f239",
X"76802e86",
X"38865682",
X"e839a454",
X"8d537852",
X"7551a0ae",
X"3f815683",
X"e0800882",
X"d43802be",
X"05330284",
X"05bd0533",
X"71882b07",
X"595d77ab",
X"380280ce",
X"05330284",
X"0580cd05",
X"3371982b",
X"71902b07",
X"973d3370",
X"882b7207",
X"02940580",
X"cb053371",
X"0754525e",
X"57595602",
X"b7053378",
X"71290288",
X"05b60533",
X"028c05b5",
X"05337188",
X"2b07701d",
X"707f8c05",
X"0c5f5957",
X"595d8e3d",
X"33821b34",
X"02b90533",
X"903d3371",
X"882b075a",
X"5c78841b",
X"2302bb05",
X"33028405",
X"ba053371",
X"882b0756",
X"5c74ab38",
X"0280ca05",
X"33028405",
X"80c90533",
X"71982b71",
X"902b0796",
X"3d337088",
X"2b720702",
X"940580c7",
X"05337107",
X"51525357",
X"5e5c7476",
X"31783179",
X"842a903d",
X"33547171",
X"31535656",
X"80d2823f",
X"83e08008",
X"82057088",
X"1c0c83e0",
X"8008e08a",
X"05565674",
X"83dffe26",
X"83388257",
X"83fff676",
X"27853883",
X"57893986",
X"5676802e",
X"80db3876",
X"7a347683",
X"2e098106",
X"b0380280",
X"d6053302",
X"840580d5",
X"05337198",
X"2b71902b",
X"07993d33",
X"70882b72",
X"07029405",
X"80d30533",
X"71077f90",
X"050c525e",
X"57585686",
X"39771b90",
X"1b0c841a",
X"228c1b08",
X"1971842a",
X"05941c0c",
X"5d800b81",
X"1b347983",
X"e0900c80",
X"567583e0",
X"800c973d",
X"0d04e93d",
X"0d83e090",
X"08568554",
X"75802e81",
X"8238800b",
X"81173499",
X"3de01146",
X"6a548a3d",
X"705458ec",
X"0551f6e5",
X"3f83e080",
X"085483e0",
X"800880df",
X"38893d33",
X"5473802e",
X"913802ab",
X"05337084",
X"2a810651",
X"5574802e",
X"86388354",
X"80c13976",
X"51f4893f",
X"83e08008",
X"a0170c02",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"9c1c0c52",
X"78981b0c",
X"53565957",
X"810b8117",
X"34745473",
X"83e0800c",
X"993d0d04",
X"f53d0d7d",
X"7f617283",
X"e090085a",
X"5d5d595c",
X"807b0c85",
X"5775802e",
X"81e03881",
X"16338106",
X"55845774",
X"802e81d2",
X"38913974",
X"81173486",
X"39800b81",
X"17348157",
X"81c0399c",
X"16089817",
X"08315574",
X"78278338",
X"74587780",
X"2e81a938",
X"98160870",
X"83ff0656",
X"577480cf",
X"38821633",
X"ff057789",
X"2a067081",
X"ff065a55",
X"78a03876",
X"8738a016",
X"08558d39",
X"a4160851",
X"f0e93f83",
X"e0800855",
X"817527ff",
X"a83874a4",
X"170ca416",
X"0851f283",
X"3f83e080",
X"085583e0",
X"8008802e",
X"ff893883",
X"e0800819",
X"a8170c98",
X"160883ff",
X"06848071",
X"31515577",
X"75278338",
X"77557483",
X"ffff0654",
X"98160883",
X"ff0653a8",
X"16085279",
X"577b8338",
X"7b577651",
X"9ad43f83",
X"e08008fe",
X"d0389816",
X"08159817",
X"0c741a78",
X"76317c08",
X"177d0c59",
X"5afed339",
X"80577683",
X"e0800c8d",
X"3d0d04fa",
X"3d0d7883",
X"e0900855",
X"56855573",
X"802e81e3",
X"38811433",
X"81065384",
X"5572802e",
X"81d5389c",
X"14085372",
X"76278338",
X"72569814",
X"0857800b",
X"98150c75",
X"802e81b9",
X"38821433",
X"70892b56",
X"5376802e",
X"b7387452",
X"ff165180",
X"cd833f83",
X"e08008ff",
X"18765470",
X"53585380",
X"ccf33f83",
X"e0800873",
X"26963874",
X"30707806",
X"7098170c",
X"777131a4",
X"17085258",
X"51538939",
X"a0140870",
X"a4160c53",
X"747627b9",
X"387251ee",
X"d63f83e0",
X"80085381",
X"0b83e080",
X"08278b38",
X"88140883",
X"e0800826",
X"8838800b",
X"811534b0",
X"3983e080",
X"08a4150c",
X"98140815",
X"98150c75",
X"753156c4",
X"39981408",
X"16709816",
X"0c735256",
X"efc53f83",
X"e080088c",
X"3883e080",
X"08811534",
X"81559439",
X"821433ff",
X"0576892a",
X"0683e080",
X"0805a815",
X"0c805574",
X"83e0800c",
X"883d0d04",
X"ef3d0d63",
X"56855583",
X"e0900880",
X"2e80d238",
X"933df405",
X"84170c64",
X"53883d70",
X"53765257",
X"f1cf3f83",
X"e0800855",
X"83e08008",
X"b438883d",
X"33547380",
X"2ea13802",
X"a7053370",
X"842a7081",
X"06515555",
X"83557380",
X"2e973876",
X"51eef53f",
X"83e08008",
X"88170c75",
X"51efa63f",
X"83e08008",
X"557483e0",
X"800c933d",
X"0d04e43d",
X"0d6ea13d",
X"08405e85",
X"5683e090",
X"08802e84",
X"85389e3d",
X"f405841f",
X"0c7e9838",
X"7d51eef5",
X"3f83e080",
X"085683ee",
X"39814181",
X"f6398341",
X"81f13993",
X"3d7f9605",
X"4159807f",
X"8295055e",
X"56756081",
X"ff053483",
X"41901e08",
X"762e81d3",
X"38a0547d",
X"2270852b",
X"83e00654",
X"58901e08",
X"52785196",
X"dd3f83e0",
X"80084183",
X"e08008ff",
X"b8387833",
X"5c7b802e",
X"ffb4388b",
X"193370bf",
X"06718106",
X"52435574",
X"802e80de",
X"387b81bf",
X"0655748f",
X"2480d338",
X"9a193355",
X"7480cb38",
X"f31d7058",
X"5d815675",
X"8b2e0981",
X"0685388e",
X"568b3975",
X"9a2e0981",
X"0683389c",
X"56751970",
X"70810552",
X"33713381",
X"1a821a5f",
X"5b525b55",
X"74863879",
X"77348539",
X"80df7734",
X"777b5757",
X"7aa02e09",
X"8106c038",
X"81567b81",
X"e5327030",
X"709f2a51",
X"51557bae",
X"2e933874",
X"802e8e38",
X"61832a70",
X"81065155",
X"74802e97",
X"387d51ed",
X"df3f83e0",
X"80084183",
X"e0800887",
X"38901e08",
X"feaf3880",
X"60347580",
X"2e88387c",
X"527f518e",
X"833f6080",
X"2e863880",
X"0b901f0c",
X"60566083",
X"2e853860",
X"81d03889",
X"1f57901e",
X"08802e81",
X"a8388056",
X"75197033",
X"515574a0",
X"2ea03874",
X"852e0981",
X"06843881",
X"e5557477",
X"70810559",
X"34811670",
X"81ff0657",
X"55877627",
X"d7388819",
X"335574a0",
X"2ea938ae",
X"77708105",
X"59348856",
X"75197033",
X"515574a0",
X"2e953874",
X"77708105",
X"59348116",
X"7081ff06",
X"57558a76",
X"27e2388b",
X"19337f88",
X"05349f19",
X"339e1a33",
X"71982b71",
X"902b079d",
X"1c337088",
X"2b72079c",
X"1e337107",
X"640c5299",
X"1d33981e",
X"3371882b",
X"07535153",
X"57595674",
X"7f840523",
X"97193396",
X"1a337188",
X"2b075656",
X"747f8605",
X"23807734",
X"7d51ebf0",
X"3f83e080",
X"08833270",
X"30707207",
X"9f2c83e0",
X"80080652",
X"5656961f",
X"3355748a",
X"38891f52",
X"961f518c",
X"8f3f7583",
X"e0800c9e",
X"3d0d04f4",
X"3d0d7e8f",
X"3dec1156",
X"56589053",
X"f0155277",
X"51e0d23f",
X"83e08008",
X"80d73878",
X"902e0981",
X"0680ce38",
X"02ab0533",
X"80f9d00b",
X"80f9d033",
X"5758568c",
X"3974762e",
X"8a388417",
X"70335657",
X"74f33876",
X"33705755",
X"74802ead",
X"38821722",
X"708a2b90",
X"3dec0556",
X"70555656",
X"84888080",
X"527751e0",
X"803f83e0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583e0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"558b953f",
X"83e08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"8114518a",
X"ad3f83e0",
X"80083070",
X"83e08008",
X"07802583",
X"e0800c53",
X"863d0d04",
X"fc3d0d76",
X"705255e6",
X"ed3f83e0",
X"80085481",
X"5383e080",
X"0880c138",
X"7451e6b0",
X"3f83e080",
X"0880f6fc",
X"5383e080",
X"085253ff",
X"913f83e0",
X"8008a138",
X"80f78052",
X"7251ff82",
X"3f83e080",
X"08923880",
X"f7845272",
X"51fef33f",
X"83e08008",
X"802e8338",
X"81547353",
X"7283e080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"e68c3f81",
X"5383e080",
X"08983873",
X"51e5d53f",
X"83e38808",
X"5283e080",
X"0851feba",
X"3f83e080",
X"08537283",
X"e0800c85",
X"3d0d04df",
X"3d0da43d",
X"0870525e",
X"dbf33f83",
X"e0800833",
X"953d5654",
X"73963880",
X"fd8c5274",
X"51898d3f",
X"9a397d52",
X"7851defb",
X"3f84d039",
X"7d51dbd9",
X"3f83e080",
X"08527451",
X"db893f80",
X"43804280",
X"41804083",
X"e3900852",
X"943d7052",
X"5de1e33f",
X"83e08008",
X"59800b83",
X"e0800855",
X"5b83e080",
X"087b2e94",
X"38811b74",
X"525be4e5",
X"3f83e080",
X"085483e0",
X"8008ee38",
X"805aff5f",
X"7909709f",
X"2c7b065b",
X"547a7a24",
X"8438ff1b",
X"5af61a70",
X"09709f2c",
X"72067bff",
X"125a5a52",
X"55558075",
X"25953876",
X"51e4aa3f",
X"83e08008",
X"76ff1858",
X"55577380",
X"24ed3874",
X"7f2e8638",
X"a1b53f74",
X"5f78ff1b",
X"70585d58",
X"807a2595",
X"387751e4",
X"803f83e0",
X"800876ff",
X"18585558",
X"738024ed",
X"38800b83",
X"e7c00c80",
X"0b83e7e8",
X"0c80f788",
X"518d8c3f",
X"81800b83",
X"e7e80c80",
X"f790518c",
X"fe3fa80b",
X"83e7c00c",
X"76802e80",
X"e43883e7",
X"c0087779",
X"32703070",
X"72078025",
X"70872b83",
X"e7e80c51",
X"56785356",
X"56e3b73f",
X"83e08008",
X"802e8838",
X"80f79851",
X"8cc53f76",
X"51e2f93f",
X"83e08008",
X"5280f8b8",
X"518cb43f",
X"7651e381",
X"3f83e080",
X"0883e7c0",
X"08555775",
X"74258638",
X"a81656f7",
X"397583e7",
X"c00c86f0",
X"7624ff98",
X"3887980b",
X"83e7c00c",
X"77802eb1",
X"387751e2",
X"b73f83e0",
X"80087852",
X"55e2d73f",
X"80f7a054",
X"83e08008",
X"8d388739",
X"80763481",
X"d03980f7",
X"9c547453",
X"735280f6",
X"f0518bd3",
X"3f805480",
X"f6f8518b",
X"ca3f8114",
X"5473a82e",
X"098106ef",
X"38868da0",
X"519da83f",
X"8052903d",
X"70525780",
X"c2e73f83",
X"52765180",
X"c2df3f62",
X"818f3861",
X"802e80fb",
X"387b5473",
X"ff2e9638",
X"78802e81",
X"8a387851",
X"e1db3f83",
X"e08008ff",
X"155559e7",
X"3978802e",
X"80f53878",
X"51e1d73f",
X"83e08008",
X"802efc8e",
X"387851e1",
X"9f3f83e0",
X"80085280",
X"f6ec5183",
X"e03f83e0",
X"8008a338",
X"7c518598",
X"3f83e080",
X"085574ff",
X"16565480",
X"7425ae38",
X"741d7033",
X"555673af",
X"2efecd38",
X"e9397851",
X"e0e03f83",
X"e0800852",
X"7c5184d0",
X"3f8f397f",
X"88296010",
X"057a0561",
X"055afc90",
X"3962802e",
X"fbd13880",
X"52765180",
X"c1bf3fa3",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067084",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d38a8",
X"0b9088b8",
X"34b80b90",
X"88b83470",
X"83e0800c",
X"823d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"852a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"980b9088",
X"b834b80b",
X"9088b834",
X"7083e080",
X"0c823d0d",
X"04930b90",
X"88bc34ff",
X"0b9088a8",
X"3404ff3d",
X"0d028f05",
X"3352800b",
X"9088bc34",
X"8a519aef",
X"3fdf3f80",
X"f80b9088",
X"a034800b",
X"90888834",
X"fa125271",
X"90888034",
X"800b9088",
X"98347190",
X"88903490",
X"88b85280",
X"7234b872",
X"34833d0d",
X"04803d0d",
X"028b0533",
X"51709088",
X"b434febf",
X"3f83e080",
X"08802ef6",
X"38823d0d",
X"04803d0d",
X"8439a5a4",
X"3ffed93f",
X"83e08008",
X"802ef338",
X"9088b433",
X"7081ff06",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"a30b9088",
X"bc34ff0b",
X"9088a834",
X"9088b851",
X"a87134b8",
X"7134823d",
X"0d04803d",
X"0d9088bc",
X"3370982b",
X"70802583",
X"e0800c51",
X"51823d0d",
X"04803d0d",
X"9088b833",
X"7081ff06",
X"70832a81",
X"32708106",
X"51515151",
X"70802ee8",
X"38b00b90",
X"88b834b8",
X"0b9088b8",
X"34823d0d",
X"04803d0d",
X"9080ac08",
X"810683e0",
X"800c823d",
X"0d04fd3d",
X"0d757754",
X"54807325",
X"94387370",
X"81055533",
X"5280f7a4",
X"5187843f",
X"ff1353e9",
X"39853d0d",
X"04fd3d0d",
X"75775354",
X"73335170",
X"89387133",
X"5170802e",
X"a1387333",
X"72335253",
X"72712785",
X"38ff5194",
X"39707327",
X"85388151",
X"8b398114",
X"81135354",
X"d3398051",
X"7083e080",
X"0c853d0d",
X"04fd3d0d",
X"75775454",
X"72337081",
X"ff065252",
X"70802ea3",
X"387181ff",
X"068114ff",
X"bf125354",
X"52709926",
X"8938a012",
X"7081ff06",
X"53517174",
X"70810556",
X"34d23980",
X"7434853d",
X"0d04ffbd",
X"3d0d80c6",
X"3d0852a5",
X"3d705254",
X"ffb33f80",
X"c73d0852",
X"853d7052",
X"53ffa63f",
X"72527351",
X"fedf3f80",
X"c53d0d04",
X"fe3d0d74",
X"76535371",
X"70810553",
X"33517073",
X"70810555",
X"3470f038",
X"843d0d04",
X"fe3d0d74",
X"52807233",
X"52537073",
X"2e8d3881",
X"12811471",
X"33535452",
X"70f53872",
X"83e0800c",
X"843d0d04",
X"f63d0d7c",
X"7e60625a",
X"5d5b5680",
X"59815585",
X"39747a29",
X"55745275",
X"51b9da3f",
X"83e08008",
X"7a27ee38",
X"74802e80",
X"dd387452",
X"7551b9c5",
X"3f83e080",
X"08755376",
X"5254b9c9",
X"3f83e080",
X"087a5375",
X"5256b9ad",
X"3f83e080",
X"08793070",
X"7b079f2a",
X"70778024",
X"07515154",
X"55728738",
X"83e08008",
X"c5387681",
X"18b01655",
X"58588974",
X"258b38b7",
X"14537a85",
X"3880d714",
X"53727834",
X"811959ff",
X"9f398077",
X"348c3d0d",
X"04f73d0d",
X"7b7d7f62",
X"029005bb",
X"05335759",
X"565a5ab0",
X"58728338",
X"a0587570",
X"70810552",
X"33715954",
X"55903980",
X"74258e38",
X"ff147770",
X"81055933",
X"545472ef",
X"3873ff15",
X"55538073",
X"25893877",
X"52795178",
X"2def3975",
X"33755753",
X"72802e90",
X"38725279",
X"51782d75",
X"70810557",
X"3353ed39",
X"8b3d0d04",
X"ee3d0d64",
X"66696970",
X"70810552",
X"335b4a5c",
X"5e5e7680",
X"2e82f938",
X"76a52e09",
X"810682e0",
X"38807041",
X"67707081",
X"05523371",
X"4a59575f",
X"76b02e09",
X"81068c38",
X"75708105",
X"57337648",
X"57815fd0",
X"17567589",
X"2680da38",
X"76675c59",
X"805c9339",
X"778a2480",
X"c3387b8a",
X"29187b70",
X"81055d33",
X"5a5cd019",
X"7081ff06",
X"58588977",
X"27a438ff",
X"9f197081",
X"ff06ffa9",
X"1b5a5156",
X"85762792",
X"38ffbf19",
X"7081ff06",
X"51567585",
X"268a38c9",
X"19587780",
X"25ffb938",
X"7a477b40",
X"7881ff06",
X"577680e4",
X"2e80e538",
X"7680e424",
X"a7387680",
X"d82e8186",
X"387680d8",
X"24903876",
X"802e81cc",
X"3876a52e",
X"81b63881",
X"b9397680",
X"e32e818c",
X"3881af39",
X"7680f52e",
X"9b387680",
X"f5248b38",
X"7680f32e",
X"81813881",
X"99397680",
X"f82e80ca",
X"38818f39",
X"913d7055",
X"5780538a",
X"5279841b",
X"7108535b",
X"56fc813f",
X"7655ab39",
X"79841b71",
X"08943d70",
X"5b5b525b",
X"56758025",
X"8c387530",
X"56ad7834",
X"0280c105",
X"57765480",
X"538a5275",
X"51fbd53f",
X"77557e54",
X"b839913d",
X"70557780",
X"d8327030",
X"70802556",
X"51585690",
X"5279841b",
X"7108535b",
X"57fbb13f",
X"7555db39",
X"79841b83",
X"1233545b",
X"56983979",
X"841b7108",
X"575b5680",
X"547f537c",
X"527d51fc",
X"9c3f8739",
X"76527d51",
X"7c2d6670",
X"33588105",
X"47fd8339",
X"943d0d04",
X"7283e094",
X"0c7183e0",
X"980c04fb",
X"3d0d883d",
X"70708405",
X"52085754",
X"755383e0",
X"94085283",
X"e0980851",
X"fcc63f87",
X"3d0d04ff",
X"3d0d7370",
X"08535102",
X"93053372",
X"34700881",
X"05710c83",
X"3d0d04fc",
X"3d0d873d",
X"88115578",
X"54bdbf53",
X"51fc993f",
X"8052873d",
X"51d13f86",
X"3d0d04fc",
X"3d0d7655",
X"7483e39c",
X"082eaf38",
X"80537451",
X"87c13f83",
X"e0800881",
X"ff06ff14",
X"7081ff06",
X"7230709f",
X"2a515255",
X"53547280",
X"2e843871",
X"dd3873fe",
X"387483e3",
X"9c0c863d",
X"0d04ff3d",
X"0dff0b83",
X"e39c0c84",
X"a53f8151",
X"87853f83",
X"e0800881",
X"ff065271",
X"ee3881d3",
X"3f7183e0",
X"800c833d",
X"0d04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"823f7280",
X"2ea03883",
X"e3b01433",
X"75708105",
X"57348114",
X"7083ffff",
X"06ff1570",
X"83ffff06",
X"56525552",
X"dd39800b",
X"83e0800c",
X"863d0d04",
X"fc3d0d76",
X"787a1156",
X"53558053",
X"71742e93",
X"38721551",
X"703383e3",
X"b0133481",
X"12811454",
X"52ea3980",
X"0b83e080",
X"0c863d0d",
X"04fd3d0d",
X"905483e3",
X"9c085186",
X"f43f83e0",
X"800881ff",
X"06ff1571",
X"30713070",
X"73079f2a",
X"729f2a06",
X"52555255",
X"5372db38",
X"853d0d04",
X"803d0d83",
X"e3a80810",
X"83e3a008",
X"079080a8",
X"0c823d0d",
X"04800b83",
X"e3a80ce4",
X"3f04810b",
X"83e3a80c",
X"db3f04ed",
X"3f047183",
X"e3a40c04",
X"803d0d80",
X"51f43f81",
X"0b83e3a8",
X"0c810b83",
X"e3a00cff",
X"bb3f823d",
X"0d04803d",
X"0d723070",
X"74078025",
X"83e3a00c",
X"51ffa53f",
X"823d0d04",
X"803d0d02",
X"8b053390",
X"80a40c90",
X"80a80870",
X"81065151",
X"70f53890",
X"80a40870",
X"81ff0683",
X"e0800c51",
X"823d0d04",
X"803d0d81",
X"ff51d13f",
X"83e08008",
X"81ff0683",
X"e0800c82",
X"3d0d0480",
X"3d0d7390",
X"2b730790",
X"80b40c82",
X"3d0d0404",
X"fb3d0d78",
X"0284059f",
X"05337098",
X"2b555755",
X"7280259b",
X"387580ff",
X"06568052",
X"80f751e0",
X"3f83e080",
X"0881ff06",
X"54738126",
X"80ff3880",
X"51fee73f",
X"ffa23f81",
X"51fedf3f",
X"ff9a3f75",
X"51feed3f",
X"74982a51",
X"fee63f74",
X"902a7081",
X"ff065253",
X"feda3f74",
X"882a7081",
X"ff065253",
X"fece3f74",
X"81ff0651",
X"fec63f81",
X"557580c0",
X"2e098106",
X"86388195",
X"558d3975",
X"80c82e09",
X"81068438",
X"81875574",
X"51fea53f",
X"8a55fec8",
X"3f83e080",
X"0881ff06",
X"70982b54",
X"54728025",
X"8c38ff15",
X"7081ff06",
X"565374e2",
X"387383e0",
X"800c873d",
X"0d04fa3d",
X"0dfdc53f",
X"8051fdda",
X"3f8a54fe",
X"933fff14",
X"7081ff06",
X"555373f3",
X"38737453",
X"5580c051",
X"fea63f83",
X"e0800881",
X"ff065473",
X"812e0981",
X"06829f38",
X"83aa5280",
X"c851fe8c",
X"3f83e080",
X"0881ff06",
X"5372812e",
X"09810681",
X"a8387454",
X"873d7411",
X"5456fdc8",
X"3f83e080",
X"08733481",
X"147081ff",
X"06555383",
X"7427e538",
X"029a0533",
X"5372812e",
X"09810681",
X"d938029b",
X"05335380",
X"ce905472",
X"81aa2e8d",
X"3881c739",
X"80e4518b",
X"9a3fff14",
X"5473802e",
X"81b83882",
X"0a5281e9",
X"51fda53f",
X"83e08008",
X"81ff0653",
X"72de3872",
X"5280fa51",
X"fd923f83",
X"e0800881",
X"ff065372",
X"81903872",
X"54731653",
X"fcd63f83",
X"e0800873",
X"34811470",
X"81ff0655",
X"53837427",
X"e838873d",
X"3370862a",
X"70810651",
X"54548c55",
X"7280e338",
X"845580de",
X"39745281",
X"e951fccc",
X"3f83e080",
X"0881ff06",
X"53825581",
X"e9568173",
X"27863873",
X"5580c156",
X"80ce9054",
X"8a3980e4",
X"518a8c3f",
X"ff145473",
X"802ea938",
X"80527551",
X"fc9a3f83",
X"e0800881",
X"ff065372",
X"e1388480",
X"5280d051",
X"fc863f83",
X"e0800881",
X"ff065372",
X"802e8338",
X"80557483",
X"e3ac3480",
X"51fb873f",
X"fbc23f88",
X"3d0d04fb",
X"3d0d7754",
X"800b83e3",
X"ac337083",
X"2a708106",
X"51555755",
X"72752e09",
X"81068538",
X"73892b54",
X"735280d1",
X"51fbbd3f",
X"83e08008",
X"81ff0653",
X"72bd3882",
X"b8c054fb",
X"833f83e0",
X"800881ff",
X"06537281",
X"ff2e0981",
X"068938ff",
X"145473e7",
X"389f3972",
X"81fe2e09",
X"81069638",
X"83e7b052",
X"83e3b051",
X"faed3ffa",
X"d33ffad0",
X"3f833981",
X"558051fa",
X"893ffac4",
X"3f7481ff",
X"0683e080",
X"0c873d0d",
X"04fb3d0d",
X"7783e3b0",
X"56548151",
X"f9ec3f83",
X"e3ac3370",
X"832a7081",
X"06515456",
X"72853873",
X"892b5473",
X"5280d851",
X"fab63f83",
X"e0800881",
X"ff065372",
X"80e43881",
X"ff51f9d4",
X"3f81fe51",
X"f9ce3f84",
X"80537470",
X"81055633",
X"51f9c13f",
X"ff137083",
X"ffff0651",
X"5372eb38",
X"7251f9b0",
X"3f7251f9",
X"ab3ff9d0",
X"3f83e080",
X"089f0653",
X"a7885472",
X"852e8c38",
X"993980e4",
X"5187c43f",
X"ff1454f9",
X"b33f83e0",
X"800881ff",
X"2e843873",
X"e9388051",
X"f8e43ff9",
X"9f3f800b",
X"83e0800c",
X"873d0d04",
X"7183e7b4",
X"0c888080",
X"0b83e7b0",
X"0c848080",
X"0b83e7b8",
X"0c04fd3d",
X"0d777017",
X"557705ff",
X"1a535371",
X"ff2e9438",
X"73708105",
X"55335170",
X"73708105",
X"5534ff12",
X"52e93985",
X"3d0d04fb",
X"3d0d87a6",
X"810b83e7",
X"b4085656",
X"753383a6",
X"801634a0",
X"5483a080",
X"5383e7b4",
X"085283e7",
X"b00851ff",
X"b13fa054",
X"83a48053",
X"83e7b408",
X"5283e7b0",
X"0851ff9e",
X"3f905483",
X"a8805383",
X"e7b40852",
X"83e7b008",
X"51ff8b3f",
X"a0538052",
X"83e7b808",
X"83a08005",
X"5186953f",
X"a0538052",
X"83e7b808",
X"83a48005",
X"5186853f",
X"90538052",
X"83e7b808",
X"83a88005",
X"5185f53f",
X"ff763483",
X"a0805480",
X"5383e7b4",
X"085283e7",
X"b80851fe",
X"c53f80d0",
X"805483b0",
X"805383e7",
X"b4085283",
X"e7b80851",
X"feb03f87",
X"ba3fa254",
X"805383e7",
X"b8088c80",
X"055280fa",
X"c451fe9a",
X"3f860b87",
X"a8833480",
X"0b87a882",
X"34800b87",
X"a09a34af",
X"0b87a096",
X"34bf0b87",
X"a0973480",
X"0b87a098",
X"349f0b87",
X"a0993480",
X"0b87a09b",
X"34e00b87",
X"a88934a2",
X"0b87a880",
X"34830b87",
X"a48f3482",
X"0b87a881",
X"34873d0d",
X"04fc3d0d",
X"83a08054",
X"805383e7",
X"b8085283",
X"e7b40851",
X"fdb83f80",
X"d0805483",
X"b0805383",
X"e7b80852",
X"83e7b408",
X"51fda33f",
X"a05483a0",
X"805383e7",
X"b8085283",
X"e7b40851",
X"fd903fa0",
X"5483a480",
X"5383e7b8",
X"085283e7",
X"b40851fc",
X"fd3f9054",
X"83a88053",
X"83e7b808",
X"5283e7b4",
X"0851fcea",
X"3f83e7b4",
X"085583a6",
X"80153387",
X"a6813486",
X"3d0d04fa",
X"3d0d7870",
X"5255c1e2",
X"3f83ffff",
X"0b83e080",
X"0825a938",
X"7451c1e3",
X"3f83e080",
X"089e3883",
X"e0800857",
X"883dfc05",
X"54848080",
X"5383e7b4",
X"08527451",
X"ffbf953f",
X"ffbedb3f",
X"883d0d04",
X"fa3d0d78",
X"705255c1",
X"a13f83ff",
X"ff0b83e0",
X"80082596",
X"38805788",
X"3dfc0554",
X"84808053",
X"83e7b408",
X"527451c0",
X"943f883d",
X"0d04803d",
X"0d908090",
X"08810683",
X"e0800c82",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe067607",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"812c8106",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fd06",
X"76100772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087082",
X"2cbf0683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fe8306",
X"76822b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"882c8706",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f1ff",
X"0676882b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70912cbf",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870fc",
X"87ffff06",
X"76912b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"992c8106",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870ffbf",
X"0a067699",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908080",
X"0870882c",
X"810683e0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"80087089",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8a2c8106",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708b2c81",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708c2c",
X"bf0683e0",
X"800c5182",
X"3d0d04fe",
X"3d0d7481",
X"e629872a",
X"9080a00c",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d848080",
X"53805288",
X"800a51ff",
X"b33f8180",
X"80538052",
X"82800a51",
X"c63f843d",
X"0d04803d",
X"0d8151fc",
X"aa3f7280",
X"2e903880",
X"51fdfe3f",
X"cd3f83e7",
X"bc3351fd",
X"f43f8151",
X"fcbb3f80",
X"51fcb63f",
X"8051fc87",
X"3f823d0d",
X"04fd3d0d",
X"75528054",
X"80ff7225",
X"8838810b",
X"ff801353",
X"54ffbf12",
X"51709926",
X"8638e012",
X"52b039ff",
X"9f125199",
X"7127a738",
X"d012e013",
X"54517089",
X"26853872",
X"52983972",
X"8f268538",
X"72528f39",
X"71ba2e09",
X"81068538",
X"9a528339",
X"80527380",
X"2e853881",
X"80125271",
X"81ff0683",
X"e0800c85",
X"3d0d0480",
X"3d0d84d8",
X"c0518071",
X"70810553",
X"347084e0",
X"c02e0981",
X"06f03882",
X"3d0d04fe",
X"3d0d0297",
X"053351fe",
X"f43f83e0",
X"800881ff",
X"0683e7c0",
X"08545280",
X"73249b38",
X"83e7e408",
X"137283e7",
X"e8080753",
X"53717334",
X"83e7c008",
X"810583e7",
X"c00c843d",
X"0d04fa3d",
X"0d82800a",
X"1b558057",
X"883dfc05",
X"54795374",
X"527851ff",
X"baab3f88",
X"3d0d04fe",
X"3d0d83e7",
X"d8085274",
X"51c18f3f",
X"83e08008",
X"8c387653",
X"755283e7",
X"d80851c6",
X"3f843d0d",
X"04fe3d0d",
X"83e7d808",
X"53755274",
X"51ffbbcd",
X"3f83e080",
X"088d3877",
X"53765283",
X"e7d80851",
X"ffa03f84",
X"3d0d04fe",
X"3d0d83e7",
X"d80851ff",
X"bac03f83",
X"e0800881",
X"80802e09",
X"81068738",
X"8f808053",
X"9b3983e7",
X"d80851ff",
X"baa43f83",
X"e0800880",
X"d0802e09",
X"81069238",
X"8fb08053",
X"83e08008",
X"5283e7d8",
X"0851fed6",
X"3f843d0d",
X"04803d0d",
X"f9fe3f83",
X"e0800884",
X"2980fae8",
X"05700883",
X"e0800c51",
X"823d0d04",
X"ed3d0d80",
X"44804380",
X"42804180",
X"705a5bfd",
X"ce3f800b",
X"83e7c00c",
X"800b83e7",
X"e80c80f7",
X"f051e9c7",
X"3f81800b",
X"83e7e80c",
X"80f7f451",
X"e9b93f80",
X"d00b83e7",
X"c00c7830",
X"707a0780",
X"2570872b",
X"83e7e80c",
X"5155f8ef",
X"3f83e080",
X"085280f7",
X"fc51e993",
X"3f80f80b",
X"83e7c00c",
X"78813270",
X"30707207",
X"80257087",
X"2b83e7e8",
X"0c515656",
X"9ced3f83",
X"e0800852",
X"80f88c51",
X"e8e93f81",
X"a00b83e7",
X"c00c7882",
X"32703070",
X"72078025",
X"70872b83",
X"e7e80c51",
X"5656fec5",
X"3f83e080",
X"085280f8",
X"9c51e8bf",
X"3f81c80b",
X"83e7c00c",
X"78833270",
X"30707207",
X"80257087",
X"2b83e7e8",
X"0c515683",
X"e7d80852",
X"56ffb599",
X"3f83e080",
X"085280f8",
X"a451e88f",
X"3f82980b",
X"83e7c00c",
X"810b83e7",
X"c45b5883",
X"e7c00883",
X"197a3270",
X"30707207",
X"80257087",
X"2b83e7e8",
X"0c51578e",
X"3d7055ff",
X"1b545757",
X"579aaf3f",
X"79708405",
X"5b0851ff",
X"b4cf3f74",
X"5483e080",
X"08537752",
X"80f8ac51",
X"e7c13fa8",
X"1783e7c0",
X"0c811858",
X"77852e09",
X"8106ffaf",
X"3883b80b",
X"83e7c00c",
X"78883270",
X"30707207",
X"80257087",
X"2b83e7e8",
X"0c515656",
X"f7bb3f80",
X"f8bc5583",
X"e0800880",
X"2e8f3883",
X"e7d40851",
X"ffb3fa3f",
X"83e08008",
X"55745280",
X"f8c451e6",
X"ee3f8488",
X"0b83e7c0",
X"0c788932",
X"70307072",
X"07802570",
X"872b83e7",
X"e80c5157",
X"80f8d052",
X"55e6cc3f",
X"868da051",
X"f8b53f80",
X"52913d70",
X"52559df5",
X"3f835274",
X"519dee3f",
X"63557483",
X"9c386119",
X"59788025",
X"85387459",
X"90398979",
X"25853889",
X"59873978",
X"892682fb",
X"3878822b",
X"5580f6c4",
X"150804f5",
X"d63f83e0",
X"80086157",
X"5575812e",
X"09810689",
X"3883e080",
X"08105590",
X"3975ff2e",
X"09810688",
X"3883e080",
X"08812c55",
X"90752585",
X"38905588",
X"39748024",
X"83388155",
X"7451f5b0",
X"3f82b039",
X"99b43f83",
X"e0800861",
X"05557480",
X"25853880",
X"55883987",
X"75258338",
X"87557451",
X"8d973f82",
X"8e39f5a0",
X"3f83e080",
X"08610555",
X"74802585",
X"38805588",
X"39837525",
X"83388355",
X"7451f599",
X"3f81ec39",
X"60873862",
X"802e81e3",
X"3883e38c",
X"0883e388",
X"0caded0b",
X"83e3900c",
X"83e7d808",
X"51d5e43f",
X"fa913f81",
X"c6396056",
X"80762598",
X"38ad8c0b",
X"83e3900c",
X"83e7b415",
X"70085255",
X"d5c53f74",
X"08529239",
X"75802592",
X"3883e7b4",
X"150851ff",
X"b1c13f80",
X"52fc1951",
X"b8396280",
X"2e818c38",
X"83e7b415",
X"700883e7",
X"c408720c",
X"83e7c40c",
X"fc1a7053",
X"51558be4",
X"3f83e080",
X"08568051",
X"8bda3f83",
X"e0800852",
X"745187f3",
X"3f755280",
X"5187ec3f",
X"80d53960",
X"55807525",
X"b63883e3",
X"980883e3",
X"880caded",
X"0b83e390",
X"0c83e7d4",
X"0851d4cf",
X"3f83e7d4",
X"0851d1ef",
X"3f83e080",
X"0881ff06",
X"705255f3",
X"f93f7480",
X"2e9d3881",
X"55a13974",
X"80259438",
X"83e7d408",
X"51ffb0b3",
X"3f8051f3",
X"dd3f8439",
X"6287387a",
X"802ef9b7",
X"38805574",
X"83e0800c",
X"953d0d04",
X"fe3d0df4",
X"893f83e0",
X"8008802e",
X"86388051",
X"818a39f4",
X"8e3f83e0",
X"800880fe",
X"38f4ae3f",
X"83e08008",
X"802eb938",
X"8151f1eb",
X"3f8051f3",
X"c43fede3",
X"3f800b83",
X"e7c00cf8",
X"df3f83e0",
X"800853ff",
X"0b83e7c0",
X"0cefd63f",
X"7280cb38",
X"83e7bc33",
X"51f39e3f",
X"7251f1bb",
X"3f80c039",
X"f3d63f83",
X"e0800880",
X"2eb53881",
X"51f1a83f",
X"8051f381",
X"3feda03f",
X"ad8c0b83",
X"e3900c83",
X"e7c40851",
X"d3813fff",
X"0b83e7c0",
X"0cef923f",
X"83e7c408",
X"52805185",
X"ea3f8151",
X"f4c83f84",
X"3d0d04fc",
X"3d0d800b",
X"83e7bc34",
X"84808052",
X"848a8080",
X"51ffb2f3",
X"3f83e080",
X"0880cd38",
X"89cf3f80",
X"fcfc51ff",
X"b7b23f83",
X"e0800855",
X"8e808054",
X"80c08053",
X"80f8d852",
X"83e08008",
X"51f6ae3f",
X"83e7d808",
X"5380f8e8",
X"527451ff",
X"b1fb3f83",
X"e0800884",
X"38f6bc3f",
X"83e7bc33",
X"51f1f23f",
X"8151f3de",
X"3f93ca3f",
X"8151f3d6",
X"3f8151fd",
X"eb3ffa39",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"0280f8f4",
X"0b83e38c",
X"0c80f8f8",
X"0b83e384",
X"0c80f8fc",
X"0b83e398",
X"0c80f980",
X"0b83e394",
X"0c83e08c",
X"08fc050c",
X"800b83e7",
X"c40b83e0",
X"8c08f805",
X"0c83e08c",
X"08f4050c",
X"ffb0c03f",
X"83e08008",
X"8605fc06",
X"83e08c08",
X"f0050c02",
X"83e08c08",
X"f0050831",
X"0d833d70",
X"83e08c08",
X"f8050870",
X"840583e0",
X"8c08f805",
X"0c0c51ff",
X"ad813f83",
X"e08c08f4",
X"05088105",
X"83e08c08",
X"f4050c83",
X"e08c08f4",
X"0508882e",
X"098106ff",
X"ab388484",
X"808051ea",
X"9b3fff0b",
X"83e7c00c",
X"800b83e7",
X"e80c84d8",
X"c00b83e7",
X"e40c8151",
X"eec13f81",
X"51eee63f",
X"8051eee1",
X"3f8151ef",
X"873f8251",
X"efaf3f80",
X"51efd73f",
X"8051f081",
X"3f80d1af",
X"528051de",
X"ff3ffda3",
X"3f83e08c",
X"08fc0508",
X"0d800b83",
X"e0800c87",
X"3d0d83e0",
X"8c0c0480",
X"3d0d81ff",
X"51800b83",
X"e7f81234",
X"ff115170",
X"f438823d",
X"0d04ff3d",
X"0d737033",
X"53518111",
X"33713471",
X"81123483",
X"3d0d04ff",
X"3d0d83ea",
X"9408a82e",
X"0981068b",
X"3883eaac",
X"0883ea94",
X"0c8739a8",
X"0b83ea94",
X"0c83ea94",
X"08860570",
X"81ff0652",
X"52d5873f",
X"833d0d04",
X"fb3d0d77",
X"79565680",
X"70715555",
X"52717525",
X"ac387216",
X"70337014",
X"7081ff06",
X"55515151",
X"71742789",
X"38811270",
X"81ff0653",
X"51718114",
X"7083ffff",
X"06555254",
X"747324d6",
X"387183e0",
X"800c873d",
X"0d04fb3d",
X"0d775689",
X"39fabd3f",
X"8351efaf",
X"3fd68e3f",
X"83e08008",
X"802eee38",
X"83ea9408",
X"86057081",
X"ff065253",
X"d4943f81",
X"0b9088d4",
X"34fa953f",
X"8351ef87",
X"3f9088d4",
X"337081ff",
X"06555373",
X"802eea38",
X"73862a70",
X"81065153",
X"72ffbe38",
X"73982b53",
X"80732480",
X"de38d4fe",
X"3f83e080",
X"085583e0",
X"800880cf",
X"38741675",
X"822b5454",
X"9088c013",
X"33743481",
X"15557485",
X"2e098106",
X"e8387533",
X"83e7f834",
X"81163383",
X"e7f93482",
X"163383e7",
X"fa348316",
X"3383e7fb",
X"34845283",
X"e7f851fe",
X"933f83e0",
X"800881ff",
X"06841733",
X"55537274",
X"2e8738fd",
X"ce3ffed1",
X"3980e451",
X"edf93f87",
X"3d0d04f4",
X"3d0d7e60",
X"5955805d",
X"8075822b",
X"7183ea98",
X"120c83ea",
X"b0175b5b",
X"57767934",
X"77772e83",
X"b7387652",
X"7751ffab",
X"9c3f8e3d",
X"fc055490",
X"5383ea80",
X"527751ff",
X"aad73f7c",
X"5675902e",
X"09810683",
X"933883ea",
X"8051fcde",
X"3f83ea82",
X"51fcd73f",
X"83ea8451",
X"fcd03f76",
X"83ea900c",
X"7751ffa8",
X"9c3f80f7",
X"805283e0",
X"800851ca",
X"bd3f83e0",
X"8008812e",
X"09810680",
X"d4387683",
X"eaa80c82",
X"0b83ea80",
X"34ff960b",
X"83ea8134",
X"7751ffaa",
X"e93f83e0",
X"80085583",
X"e0800877",
X"25883883",
X"e080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583ea82",
X"347483ea",
X"83347683",
X"ea8434ff",
X"800b83ea",
X"85348190",
X"3983ea80",
X"3383ea81",
X"3371882b",
X"07565b74",
X"83ffff2e",
X"09810680",
X"e838fe80",
X"0b83eaa8",
X"0c810b83",
X"ea900cff",
X"0b83ea80",
X"34ff0b83",
X"ea813477",
X"51ffa9f6",
X"3f83e080",
X"0883eab4",
X"0c83e080",
X"085583e0",
X"80088025",
X"883883e0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83ea8234",
X"7483ea83",
X"347683ea",
X"8434ff80",
X"0b83ea85",
X"34810b83",
X"ea8f34a5",
X"39748596",
X"2e098106",
X"80fe3875",
X"83eaa80c",
X"7751ffa9",
X"aa3f83ea",
X"8f3383e0",
X"80080755",
X"7483ea8f",
X"3483ea8f",
X"33810655",
X"74802e83",
X"38845783",
X"ea843383",
X"ea853371",
X"882b0756",
X"5c748180",
X"2e098106",
X"a13883ea",
X"823383ea",
X"83337188",
X"2b07565b",
X"ad807527",
X"87387682",
X"07579c39",
X"76810757",
X"96397482",
X"802e0981",
X"06873876",
X"83075787",
X"397481ff",
X"268a3877",
X"83ea981b",
X"0c767934",
X"8e3d0d04",
X"803d0d72",
X"842983ea",
X"98057008",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"727083e7",
X"f00c7084",
X"2980fcbc",
X"05700883",
X"eaac0c51",
X"51823d0d",
X"04fe3d0d",
X"8151de3f",
X"800b83e9",
X"fc0c800b",
X"83e9f80c",
X"ff0b83e7",
X"f40ca80b",
X"83ea940c",
X"ae51cec2",
X"3f800b83",
X"ea985452",
X"80737084",
X"05550c81",
X"12527184",
X"2e098106",
X"ef38843d",
X"0d04fe3d",
X"0d740284",
X"05960522",
X"53537180",
X"2e963872",
X"70810554",
X"3351cecd",
X"3fff1270",
X"83ffff06",
X"5152e739",
X"843d0d04",
X"fe3d0d02",
X"92052253",
X"82ac51e8",
X"ee3f80c3",
X"51ceaa3f",
X"819651e8",
X"e23f7252",
X"83e7f851",
X"ffb43f72",
X"5283e7f8",
X"51f8cd3f",
X"83e08008",
X"81ff0651",
X"ce873f84",
X"3d0d04ff",
X"b13d0d80",
X"d13df805",
X"51f8f73f",
X"83e9fc08",
X"810583e9",
X"fc0c80cf",
X"3d33cf11",
X"7081ff06",
X"51565674",
X"832688e6",
X"38758f06",
X"ff055675",
X"83e7f408",
X"2e9b3875",
X"83269638",
X"7583e7f4",
X"0c758429",
X"83ea9805",
X"70085355",
X"7551f9fb",
X"3f807624",
X"88c23875",
X"842983ea",
X"98055574",
X"08802e88",
X"b33883e7",
X"f4088429",
X"83ea9805",
X"70080288",
X"0582b905",
X"33525b55",
X"7480d22e",
X"84b03874",
X"80d22490",
X"3874bf2e",
X"9c387480",
X"d02e81d5",
X"3887f239",
X"7480d32e",
X"80d33874",
X"80d72e81",
X"c43887e1",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055656",
X"cd833f80",
X"c151ccbd",
X"3ff6983f",
X"83eaaf33",
X"83e7f834",
X"815283e7",
X"f851cdda",
X"3f8151fd",
X"e73f748b",
X"3883eaac",
X"0883ea94",
X"0c8739a8",
X"0b83ea94",
X"0cccce3f",
X"80c151cc",
X"883ff5e3",
X"3f900b83",
X"ea8f3381",
X"06565674",
X"802e8338",
X"985683ea",
X"843383ea",
X"85337188",
X"2b075659",
X"7481802e",
X"0981069c",
X"3883ea82",
X"3383ea83",
X"3371882b",
X"075657ad",
X"8075278c",
X"38758180",
X"07568539",
X"75a00756",
X"7583e7f8",
X"34ff0b83",
X"e7f934e0",
X"0b83e7fa",
X"34800b83",
X"e7fb3484",
X"5283e7f8",
X"51cccf3f",
X"8451869b",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055659",
X"cbc33f79",
X"51ffa3d7",
X"3f83e080",
X"08802e8a",
X"3880ce51",
X"caef3f85",
X"f13980c1",
X"51cae63f",
X"cbd73fca",
X"903f83ea",
X"a8085883",
X"75259b38",
X"83ea8433",
X"83ea8533",
X"71882b07",
X"fc177129",
X"7a058380",
X"055a5157",
X"8d397481",
X"802918ff",
X"80055881",
X"80578056",
X"76762e92",
X"38cac23f",
X"83e08008",
X"83e7f817",
X"34811656",
X"eb39cab1",
X"3f83e080",
X"0881ff06",
X"775383e7",
X"f85256f4",
X"bf3f83e0",
X"800881ff",
X"06557575",
X"2e098106",
X"81953894",
X"51e4ac3f",
X"caab3f80",
X"c151c9e5",
X"3fcad63f",
X"77527951",
X"ffa1ea3f",
X"805e80d1",
X"3dfdf405",
X"54765383",
X"e7f85279",
X"51ff9ff0",
X"3f0282b9",
X"05335581",
X"597480d7",
X"2e098106",
X"80c53877",
X"527951ff",
X"a1bb3f80",
X"d13dfdf0",
X"05547653",
X"8f3d7053",
X"7a5258ff",
X"a0f33f80",
X"5676762e",
X"a2387518",
X"83e7f817",
X"33713370",
X"72327030",
X"70802570",
X"307f0681",
X"1d5d5f51",
X"5151525b",
X"55db3982",
X"ac51e3a7",
X"3f78802e",
X"863880c3",
X"51843980",
X"ce51c8d9",
X"3fc9ca3f",
X"c8833f83",
X"d8390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290559",
X"5580705d",
X"5980e451",
X"e2f13fc8",
X"f03f80c1",
X"51c8aa3f",
X"83ea9008",
X"792e82d6",
X"3883eab4",
X"0880fc05",
X"5580fd52",
X"745185c1",
X"3f83e080",
X"085b7782",
X"24b238ff",
X"1870872b",
X"83ffff80",
X"0680fb88",
X"0583e7f8",
X"59575581",
X"80557570",
X"81055733",
X"77708105",
X"5934ff15",
X"7081ff06",
X"515574ea",
X"38828539",
X"7782e82e",
X"81a33877",
X"82e92e09",
X"810681aa",
X"38785877",
X"87327030",
X"70720780",
X"257a8a32",
X"70307072",
X"07802573",
X"0753545a",
X"51575575",
X"802e9738",
X"78782692",
X"38a00b83",
X"e7f81a34",
X"81197081",
X"ff065a55",
X"eb398118",
X"7081ff06",
X"59558a78",
X"27ffbc38",
X"8f5883e7",
X"f3183383",
X"e7f81934",
X"ff187081",
X"ff065955",
X"778426ea",
X"38905880",
X"0b83e7f8",
X"19348118",
X"7081ff06",
X"70982b52",
X"59557480",
X"25e93880",
X"c6557a85",
X"8f248438",
X"80c25574",
X"83e7f834",
X"80f10b83",
X"e7fb3481",
X"0b83e7fc",
X"347a83e7",
X"f9347a88",
X"2c557483",
X"e7fa3480",
X"cb3982f0",
X"782580c4",
X"387780fd",
X"29fd97d3",
X"05527951",
X"ff9e963f",
X"80d13dfd",
X"ec055480",
X"fd5383e7",
X"f8527951",
X"ff9dce3f",
X"7b811959",
X"567580fc",
X"24833878",
X"5877882c",
X"557483e8",
X"f5347783",
X"e8f63475",
X"83e8f734",
X"81805980",
X"cc3983ea",
X"a8085783",
X"78259b38",
X"83ea8433",
X"83ea8533",
X"71882b07",
X"fc1a7129",
X"79058380",
X"05595159",
X"8d397781",
X"802917ff",
X"80055781",
X"80597652",
X"7951ff9d",
X"a43f80d1",
X"3dfdec05",
X"54785383",
X"e7f85279",
X"51ff9cdd",
X"3f7851f6",
X"bf3fc5ed",
X"3fc4a63f",
X"8b3983e9",
X"f8088105",
X"83e9f80c",
X"80d13d0d",
X"04f6e03f",
X"fc39fc3d",
X"0d767871",
X"842983ea",
X"98057008",
X"51535353",
X"709e3880",
X"ce723480",
X"cf0b8113",
X"3480ce0b",
X"82133480",
X"c50b8313",
X"34708413",
X"3480e739",
X"83eab013",
X"335480d2",
X"72347382",
X"2a708106",
X"515180cf",
X"53708438",
X"80d75372",
X"811334a0",
X"0b821334",
X"73830651",
X"70812e9e",
X"38708124",
X"88387080",
X"2e8f389f",
X"3970822e",
X"92387083",
X"2e923893",
X"3980d855",
X"8e3980d3",
X"55893980",
X"cd558439",
X"80c45574",
X"83133480",
X"c40b8413",
X"34800b85",
X"1334863d",
X"0d0483e7",
X"f00883e0",
X"800c0480",
X"3d0d83e7",
X"f0088429",
X"80fcdc05",
X"700883e0",
X"800c5182",
X"3d0d04fc",
X"3d0d7678",
X"53548153",
X"80558739",
X"71107310",
X"54527372",
X"26517280",
X"2ea73870",
X"802e8638",
X"718025e8",
X"3872802e",
X"98387174",
X"26893873",
X"72317574",
X"07565472",
X"812a7281",
X"2a5353e5",
X"39735178",
X"83387451",
X"7083e080",
X"0c863d0d",
X"04fe3d0d",
X"80537552",
X"7451ffa3",
X"3f843d0d",
X"04fe3d0d",
X"81537552",
X"7451ff93",
X"3f843d0d",
X"04fb3d0d",
X"77795555",
X"80567476",
X"25863874",
X"30558156",
X"73802588",
X"38733076",
X"81325754",
X"80537352",
X"7451fee7",
X"3f83e080",
X"08547580",
X"2e873883",
X"e0800830",
X"547383e0",
X"800c873d",
X"0d04fa3d",
X"0d787a57",
X"55805774",
X"77258638",
X"74305581",
X"57759f2c",
X"54815375",
X"74327431",
X"527451fe",
X"aa3f83e0",
X"80085476",
X"802e8738",
X"83e08008",
X"30547383",
X"e0800c88",
X"3d0d04fd",
X"3d0d7554",
X"80740c80",
X"0b84150c",
X"800b8815",
X"0c800b8c",
X"150c87a6",
X"80337081",
X"ff067071",
X"842a0651",
X"5151dbb2",
X"3f70812a",
X"81327181",
X"32718106",
X"71810631",
X"84170c53",
X"5370832a",
X"81327182",
X"2a813270",
X"81067271",
X"31770c51",
X"525287a0",
X"903387a0",
X"91337081",
X"ff067073",
X"06813281",
X"0688180c",
X"51525283",
X"e0800880",
X"2e80c238",
X"83e08008",
X"812a7081",
X"0683e080",
X"08810631",
X"84160c51",
X"83e08008",
X"832a83e0",
X"8008822a",
X"71810671",
X"81063176",
X"0c525283",
X"e0800884",
X"2a810688",
X"150c83e0",
X"8008852a",
X"81068c15",
X"0c853d0d",
X"04fe3d0d",
X"74765452",
X"7151febb",
X"3f72812e",
X"a2388173",
X"268d3872",
X"822ea838",
X"72832e9c",
X"38e63971",
X"08e23884",
X"1208dd38",
X"881208d8",
X"38a53988",
X"1208812e",
X"9e389139",
X"88120881",
X"2e953871",
X"08913884",
X"12088c38",
X"8c120881",
X"2e098106",
X"ffb23884",
X"3d0d0400",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002b97",
X"00002bd8",
X"00002bfa",
X"00002c1c",
X"00002c42",
X"00002c42",
X"00002c42",
X"00002c42",
X"00002cb3",
X"00002d04",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"43505520",
X"54757262",
X"6f3a2564",
X"78000000",
X"44726976",
X"65205475",
X"72626f3a",
X"25730000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"4d454d00",
X"5374616e",
X"64617264",
X"00000000",
X"46617374",
X"28362900",
X"46617374",
X"28352900",
X"46617374",
X"28342900",
X"46617374",
X"28332900",
X"46617374",
X"28322900",
X"46617374",
X"28312900",
X"46617374",
X"28302900",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00003bac",
X"00003bb0",
X"00003bb8",
X"00003bc4",
X"00003bd0",
X"00003bdc",
X"00003be8",
X"00003bec",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00000028",
X"00000006",
X"00000005",
X"00000004",
X"00000003",
X"00000002",
X"00000001",
X"00000000",
X"00003c84",
X"00003c90",
X"00003c98",
X"00003ca0",
X"00003ca8",
X"00003cb0",
X"00003cb8",
X"00003cc0",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
