
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81d6",
X"a4738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81de",
X"c80c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757580f4",
X"8f2d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7580f3ce",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80de9204",
X"fd3d0d75",
X"705254ae",
X"a73f83c0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"c0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83c0",
X"8008732e",
X"a13883c0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183c0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83c2d008",
X"248a38b4",
X"f83fff0b",
X"83c2d00c",
X"800b83c0",
X"800c04ff",
X"3d0d7352",
X"83c0ac08",
X"722e8d38",
X"d93f7151",
X"96993f71",
X"83c0ac0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"558154bc",
X"15088191",
X"387451cf",
X"3f795880",
X"7a2580f7",
X"3883c380",
X"0870892a",
X"5783ff06",
X"78848072",
X"31565657",
X"73782583",
X"38735575",
X"83c2d008",
X"2e8438ff",
X"893f83c2",
X"d0088025",
X"a6387589",
X"2b5198dc",
X"3f83c380",
X"088f3dfc",
X"11555c54",
X"8152f81b",
X"5196c63f",
X"761483c3",
X"800c7583",
X"c2d00c74",
X"53765278",
X"51b3a93f",
X"83c08008",
X"83c38008",
X"1683c380",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8b3861",
X"7a710c54",
X"75547580",
X"2e833881",
X"547383c0",
X"800c8e3d",
X"0d04fc3d",
X"0dfe9b3f",
X"7651feaf",
X"3f863dfc",
X"05537852",
X"775195e9",
X"3f797571",
X"0c5483c0",
X"80085483",
X"c0800880",
X"2e833881",
X"547383c0",
X"800c863d",
X"0d04fe3d",
X"0d7583c2",
X"d0085353",
X"80722489",
X"3871732e",
X"8438fdd6",
X"3f7451fd",
X"ea3f7251",
X"97ae3f83",
X"c0800852",
X"83c08008",
X"802e8338",
X"81527183",
X"c0800c84",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"c0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"c0800c51",
X"823d0d04",
X"80c40b83",
X"c0800c04",
X"fd3d0d75",
X"77715470",
X"535553a9",
X"ff3f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfceb3f",
X"735193ab",
X"3f7383c0",
X"ac0c83c0",
X"80085383",
X"c0800880",
X"2e833881",
X"537283c0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcbf3f",
X"72802ea5",
X"38bc1308",
X"527351a9",
X"893f83c0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"c0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83c0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83c2d0",
X"0c7483c0",
X"b00c7583",
X"c2cc0caf",
X"dd3f83c0",
X"800881ff",
X"06528153",
X"71993883",
X"c2e8518e",
X"943f83c0",
X"80085283",
X"c0800880",
X"2e833872",
X"52715372",
X"83c0800c",
X"843d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"51a6fa3f",
X"83c08008",
X"557483c0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"c0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283c2cc",
X"085180e2",
X"d13f83c0",
X"800857f9",
X"e13f7952",
X"83c2d451",
X"95b73f83",
X"c0800854",
X"805383c0",
X"8008732e",
X"09810682",
X"833883c0",
X"b0080b0b",
X"81dbb853",
X"705256a6",
X"b73f0b0b",
X"81dbb852",
X"80c01651",
X"a6aa3f75",
X"bc170c73",
X"82c0170c",
X"810b82c4",
X"170c810b",
X"82c8170c",
X"7382cc17",
X"0cff1782",
X"d0175557",
X"81913983",
X"c0bc3370",
X"822a7081",
X"06515455",
X"72818038",
X"74812a81",
X"06587780",
X"f6387484",
X"2a810682",
X"c4150c83",
X"c0bc3381",
X"0682c815",
X"0c795273",
X"51a5d13f",
X"7351a5e8",
X"3f83c080",
X"081453af",
X"73708105",
X"553472bc",
X"150c83c0",
X"bd527251",
X"a5b23f83",
X"c0b40882",
X"c0150c83",
X"c0ca5280",
X"c01451a5",
X"9f3f7880",
X"2e8d3873",
X"51782d83",
X"c0800880",
X"2e993877",
X"82cc150c",
X"75802e86",
X"387382cc",
X"170c7382",
X"d015ff19",
X"59555676",
X"802e9b38",
X"83c0b452",
X"83c2d451",
X"94ad3f83",
X"c080088a",
X"3883c0bd",
X"335372fe",
X"d2387880",
X"2e893883",
X"c0b00851",
X"fcb83f83",
X"c0b00853",
X"7283c080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb53f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f690",
X"3f83c080",
X"08745387",
X"3d705355",
X"55f6b03f",
X"f7903f73",
X"51d33f63",
X"53745283",
X"c0800851",
X"fab83f92",
X"3d0d0471",
X"83c0800c",
X"0480c012",
X"83c0800c",
X"04803d0d",
X"7282c011",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"c0800c51",
X"823d0d04",
X"f93d0d79",
X"83c09008",
X"57578177",
X"27819638",
X"76881708",
X"27818e38",
X"75335574",
X"822e8938",
X"74832eb3",
X"3880fe39",
X"74547610",
X"83fe0653",
X"76882a8c",
X"17080552",
X"893dfc05",
X"51aa8b3f",
X"83c08008",
X"80df3802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d13984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"51a9db3f",
X"83c08008",
X"b038029f",
X"05330284",
X"059e0533",
X"71982b71",
X"902b0702",
X"8c059d05",
X"3370882b",
X"72078d3d",
X"337180ff",
X"fffe8006",
X"07515253",
X"57585683",
X"39815574",
X"83c0800c",
X"893d0d04",
X"fb3d0d83",
X"c09008fe",
X"19881208",
X"fe055556",
X"54805674",
X"73278d38",
X"82143375",
X"71299416",
X"08055753",
X"7583c080",
X"0c873d0d",
X"04fc3d0d",
X"7652800b",
X"83c09008",
X"70335152",
X"5370832e",
X"09810691",
X"38951233",
X"94133371",
X"982b7190",
X"2b075555",
X"519b1233",
X"9a133371",
X"882b0774",
X"0783c080",
X"0c55863d",
X"0d04fc3d",
X"0d7683c0",
X"90085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"fed63f83",
X"c0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183c080",
X"0c863d0d",
X"04fa3d0d",
X"7883c090",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fcb13f",
X"81527183",
X"c0800827",
X"a8388352",
X"83c08008",
X"88170827",
X"9c3883c0",
X"80088c16",
X"0c83c080",
X"0851fdbc",
X"3f83c080",
X"0890160c",
X"73752380",
X"527183c0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585e5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"9f269138",
X"7a51fdd2",
X"3f83c080",
X"0856807d",
X"34838139",
X"933d841c",
X"08705859",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"3880705a",
X"5c887f08",
X"5f5a7b81",
X"1d7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535e57",
X"557480e7",
X"3876ae2e",
X"09810683",
X"38815578",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675bb",
X"3888598b",
X"5affab39",
X"76982b55",
X"74802587",
X"3881d5b4",
X"173357ff",
X"9f175574",
X"99268938",
X"e0177081",
X"ff065855",
X"78811a70",
X"81ff0672",
X"1b535b57",
X"55767534",
X"fef8397b",
X"1e7f0c80",
X"5576a026",
X"83388155",
X"748b1934",
X"7a51fc82",
X"3f83c080",
X"0880f538",
X"a0547a22",
X"70852b83",
X"e0065455",
X"901b0852",
X"7c51a496",
X"3f83c080",
X"085783c0",
X"80088181",
X"387c3355",
X"74802e80",
X"f4388b1d",
X"3370832a",
X"70810651",
X"565674b4",
X"388b7d84",
X"1d0883c0",
X"8008595b",
X"5b58ff18",
X"5877ff2e",
X"9a387970",
X"81055b33",
X"79708105",
X"5b337171",
X"31525656",
X"75802ee2",
X"38863975",
X"802e9638",
X"7a51fbe5",
X"3fff8639",
X"83c08008",
X"5683c080",
X"08b63883",
X"39765684",
X"1b088b11",
X"33515574",
X"a7388b1d",
X"3370842a",
X"70810651",
X"56567489",
X"38835694",
X"39815690",
X"397c51fa",
X"943f83c0",
X"8008881c",
X"0cfd8139",
X"7583c080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"51a2db3f",
X"835683c0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"51a2af3f",
X"83c08008",
X"98388117",
X"33773371",
X"882b0783",
X"c0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"7651a286",
X"3f83c080",
X"08983881",
X"17337733",
X"71882b07",
X"83c08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583c080",
X"0c8a3d0d",
X"04eb3d0d",
X"675a800b",
X"83c0900c",
X"a1a83f83",
X"c0800881",
X"06558256",
X"7483ef38",
X"7475538f",
X"3d705357",
X"59feca3f",
X"83c08008",
X"81ff0657",
X"76812e09",
X"810680d4",
X"38905483",
X"be537452",
X"7551a19a",
X"3f83c080",
X"0880c938",
X"8f3d3355",
X"74802e80",
X"c93802bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"33710770",
X"587b575e",
X"525e5759",
X"57fdee3f",
X"83c08008",
X"81ff0657",
X"76832e09",
X"81068638",
X"815682f2",
X"3976802e",
X"86388656",
X"82e839a4",
X"548d5378",
X"527551a0",
X"b13f8156",
X"83c08008",
X"82d43802",
X"be053302",
X"8405bd05",
X"3371882b",
X"07595d77",
X"ab380280",
X"ce053302",
X"840580cd",
X"05337198",
X"2b71902b",
X"07973d33",
X"70882b72",
X"07029405",
X"80cb0533",
X"71075452",
X"5e575956",
X"02b70533",
X"78712902",
X"8805b605",
X"33028c05",
X"b5053371",
X"882b0770",
X"1d707f8c",
X"050c5f59",
X"57595d8e",
X"3d33821b",
X"3402b905",
X"33903d33",
X"71882b07",
X"5a5c7884",
X"1b2302bb",
X"05330284",
X"05ba0533",
X"71882b07",
X"565c74ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"07515253",
X"575e5c74",
X"76317831",
X"79842a90",
X"3d335471",
X"71315356",
X"5680d3b6",
X"3f83c080",
X"08820570",
X"881c0c83",
X"c08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83c0900c",
X"80567583",
X"c0800c97",
X"3d0d04e9",
X"3d0d83c0",
X"90085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e53f83c0",
X"80085483",
X"c0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f489",
X"3f83c080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383c080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83c09008",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0e93f",
X"83c08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"833f83c0",
X"80085583",
X"c0800880",
X"2eff8938",
X"83c08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"519ad73f",
X"83c08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83c0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83c09008",
X"55568555",
X"73802e81",
X"e3388114",
X"33810653",
X"84557280",
X"2e81d538",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b9388214",
X"3370892b",
X"56537680",
X"2eb73874",
X"52ff1651",
X"80ceb73f",
X"83c08008",
X"ff187654",
X"70535853",
X"80cea73f",
X"83c08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed63f83",
X"c0800853",
X"810b83c0",
X"8008278b",
X"38881408",
X"83c08008",
X"26883880",
X"0b811534",
X"b03983c0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc53f",
X"83c08008",
X"8c3883c0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683c0",
X"800805a8",
X"150c8055",
X"7483c080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83c09008",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1cf3f",
X"83c08008",
X"5583c080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef5",
X"3f83c080",
X"0888170c",
X"7551efa6",
X"3f83c080",
X"08557483",
X"c0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683c0",
X"9008802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f53f83c0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"96e03f83",
X"c0800841",
X"83c08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"eddf3f83",
X"c0800841",
X"83c08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"8e863f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f03f83c0",
X"80088332",
X"70307072",
X"079f2c83",
X"c0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"8c923f75",
X"83c0800c",
X"9e3d0d04",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"7751e0d2",
X"3f83c080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3381ded0",
X"0b81ded0",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"527751e0",
X"813f83c0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583c0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"558b993f",
X"83c08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"8114518a",
X"b13f83c0",
X"80083070",
X"83c08008",
X"07802583",
X"c0800c53",
X"863d0d04",
X"fc3d0d76",
X"705255e6",
X"ee3f83c0",
X"80085481",
X"5383c080",
X"0880c138",
X"7451e6b1",
X"3f83c080",
X"0881dbc8",
X"5383c080",
X"085253ff",
X"913f83c0",
X"8008a138",
X"81dbcc52",
X"7251ff82",
X"3f83c080",
X"08923881",
X"dbd05272",
X"51fef33f",
X"83c08008",
X"802e8338",
X"81547353",
X"7283c080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"e68d3f81",
X"5383c080",
X"08983873",
X"51e5d63f",
X"83c39808",
X"5283c080",
X"0851feba",
X"3f83c080",
X"08537283",
X"c0800c85",
X"3d0d04df",
X"3d0da43d",
X"0870525e",
X"dbfb3f83",
X"c0800833",
X"953d5654",
X"73963881",
X"e2a05274",
X"5189913f",
X"9a397d52",
X"7851defc",
X"3f84d039",
X"7d51dbe1",
X"3f83c080",
X"08527451",
X"db913f80",
X"43804280",
X"41804083",
X"c3a00852",
X"943d7052",
X"5de1e43f",
X"83c08008",
X"59800b83",
X"c0800855",
X"5b83c080",
X"087b2e94",
X"38811b74",
X"525be4e6",
X"3f83c080",
X"085483c0",
X"8008ee38",
X"805aff5f",
X"7909709f",
X"2c7b065b",
X"547a7a24",
X"8438ff1b",
X"5af61a70",
X"09709f2c",
X"72067bff",
X"125a5a52",
X"55558075",
X"25953876",
X"51e4ab3f",
X"83c08008",
X"76ff1858",
X"55577380",
X"24ed3874",
X"7f2e8638",
X"a1b93f74",
X"5f78ff1b",
X"70585d58",
X"807a2595",
X"387751e4",
X"813f83c0",
X"800876ff",
X"18585558",
X"738024ed",
X"38800b83",
X"c7d00c80",
X"0b83c884",
X"0c81dbd4",
X"518d903f",
X"81800b83",
X"c8840c81",
X"dbdc518d",
X"823fa80b",
X"83c7d00c",
X"76802e80",
X"e43883c7",
X"d0087779",
X"32703070",
X"72078025",
X"70872b83",
X"c8840c51",
X"56785356",
X"56e3b83f",
X"83c08008",
X"802e8838",
X"81dbe451",
X"8cc93f76",
X"51e2fa3f",
X"83c08008",
X"5281dd84",
X"518cb83f",
X"7651e382",
X"3f83c080",
X"0883c7d0",
X"08555775",
X"74258638",
X"a81656f7",
X"397583c7",
X"d00c86f0",
X"7624ff98",
X"3887980b",
X"83c7d00c",
X"77802eb1",
X"387751e2",
X"b83f83c0",
X"80087852",
X"55e2d83f",
X"81dbec54",
X"83c08008",
X"8d388739",
X"80763481",
X"d03981db",
X"e8547453",
X"735281db",
X"bc518bd7",
X"3f805481",
X"dbc4518b",
X"ce3f8114",
X"5473a82e",
X"098106ef",
X"38868da0",
X"519dac3f",
X"8052903d",
X"70525780",
X"c4913f83",
X"52765180",
X"c4893f62",
X"818f3861",
X"802e80fb",
X"387b5473",
X"ff2e9638",
X"78802e81",
X"8a387851",
X"e1dc3f83",
X"c08008ff",
X"155559e7",
X"3978802e",
X"80f53878",
X"51e1d83f",
X"83c08008",
X"802efc8e",
X"387851e1",
X"a03f83c0",
X"80085281",
X"dbb85183",
X"e43f83c0",
X"8008a338",
X"7c51859c",
X"3f83c080",
X"085574ff",
X"16565480",
X"7425ae38",
X"741d7033",
X"555673af",
X"2efecd38",
X"e9397851",
X"e0e13f83",
X"c0800852",
X"7c5184d4",
X"3f8f397f",
X"88296010",
X"057a0561",
X"055afc90",
X"3962802e",
X"fbd13880",
X"52765180",
X"c2e93fa3",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067084",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d38a8",
X"0b9088b8",
X"34b80b90",
X"88b83470",
X"83c0800c",
X"823d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"852a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"980b9088",
X"b834b80b",
X"9088b834",
X"7083c080",
X"0c823d0d",
X"04930b90",
X"88bc34ff",
X"0b9088a8",
X"3404ff3d",
X"0d028f05",
X"3352800b",
X"9088bc34",
X"8a519af3",
X"3fdf3f80",
X"f80b9088",
X"a034800b",
X"90888834",
X"fa125271",
X"90888034",
X"800b9088",
X"98347190",
X"88903490",
X"88b85280",
X"7234b872",
X"34833d0d",
X"04803d0d",
X"028b0533",
X"51709088",
X"b434febf",
X"3f83c080",
X"08802ef6",
X"38823d0d",
X"04803d0d",
X"8439a6b2",
X"3ffed93f",
X"83c08008",
X"802ef338",
X"9088b433",
X"7081ff06",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"a30b9088",
X"bc34ff0b",
X"9088a834",
X"9088b851",
X"a87134b8",
X"7134823d",
X"0d04803d",
X"0d9088bc",
X"337081c0",
X"06703070",
X"802583c0",
X"800c5151",
X"51823d0d",
X"04803d0d",
X"9088b833",
X"7081ff06",
X"70832a81",
X"32708106",
X"51515151",
X"70802ee8",
X"38b00b90",
X"88b834b8",
X"0b9088b8",
X"34823d0d",
X"04803d0d",
X"9080ac08",
X"810683c0",
X"800c823d",
X"0d04fd3d",
X"0d757754",
X"54807325",
X"94387370",
X"81055533",
X"5281dbf0",
X"5187843f",
X"ff1353e9",
X"39853d0d",
X"04fd3d0d",
X"75775354",
X"73335170",
X"89387133",
X"5170802e",
X"a1387333",
X"72335253",
X"72712785",
X"38ff5194",
X"39707327",
X"85388151",
X"8b398114",
X"81135354",
X"d3398051",
X"7083c080",
X"0c853d0d",
X"04fd3d0d",
X"75775454",
X"72337081",
X"ff065252",
X"70802ea3",
X"387181ff",
X"068114ff",
X"bf125354",
X"52709926",
X"8938a012",
X"7081ff06",
X"53517174",
X"70810556",
X"34d23980",
X"7434853d",
X"0d04ffbd",
X"3d0d80c6",
X"3d0852a5",
X"3d705254",
X"ffb33f80",
X"c73d0852",
X"853d7052",
X"53ffa63f",
X"72527351",
X"fedf3f80",
X"c53d0d04",
X"fe3d0d74",
X"76535371",
X"70810553",
X"33517073",
X"70810555",
X"3470f038",
X"843d0d04",
X"fe3d0d74",
X"52807233",
X"52537073",
X"2e8d3881",
X"12811471",
X"33535452",
X"70f53872",
X"83c0800c",
X"843d0d04",
X"f63d0d7c",
X"7e60625a",
X"5d5b5680",
X"59815585",
X"39747a29",
X"55745275",
X"51bb8b3f",
X"83c08008",
X"7a27ee38",
X"74802e80",
X"dd387452",
X"7551baf6",
X"3f83c080",
X"08755376",
X"5254bafa",
X"3f83c080",
X"087a5375",
X"5256bade",
X"3f83c080",
X"08793070",
X"7b079f2a",
X"70778024",
X"07515154",
X"55728738",
X"83c08008",
X"c5387681",
X"18b01655",
X"58588974",
X"258b38b7",
X"14537a85",
X"3880d714",
X"53727834",
X"811959ff",
X"9f398077",
X"348c3d0d",
X"04f73d0d",
X"7b7d7f62",
X"029005bb",
X"05335759",
X"565a5ab0",
X"58728338",
X"a0587570",
X"70810552",
X"33715954",
X"55903980",
X"74258e38",
X"ff147770",
X"81055933",
X"545472ef",
X"3873ff15",
X"55538073",
X"25893877",
X"52795178",
X"2def3975",
X"33755753",
X"72802e90",
X"38725279",
X"51782d75",
X"70810557",
X"3353ed39",
X"8b3d0d04",
X"ee3d0d64",
X"66696970",
X"70810552",
X"335b4a5c",
X"5e5e7680",
X"2e82f938",
X"76a52e09",
X"810682e0",
X"38807041",
X"67707081",
X"05523371",
X"4a59575f",
X"76b02e09",
X"81068c38",
X"75708105",
X"57337648",
X"57815fd0",
X"17567589",
X"2680da38",
X"76675c59",
X"805c9339",
X"778a2480",
X"c3387b8a",
X"29187b70",
X"81055d33",
X"5a5cd019",
X"7081ff06",
X"58588977",
X"27a438ff",
X"9f197081",
X"ff06ffa9",
X"1b5a5156",
X"85762792",
X"38ffbf19",
X"7081ff06",
X"51567585",
X"268a38c9",
X"19587780",
X"25ffb938",
X"7a477b40",
X"7881ff06",
X"577680e4",
X"2e80e538",
X"7680e424",
X"a7387680",
X"d82e8186",
X"387680d8",
X"24903876",
X"802e81cc",
X"3876a52e",
X"81b63881",
X"b9397680",
X"e32e818c",
X"3881af39",
X"7680f52e",
X"9b387680",
X"f5248b38",
X"7680f32e",
X"81813881",
X"99397680",
X"f82e80ca",
X"38818f39",
X"913d7055",
X"5780538a",
X"5279841b",
X"7108535b",
X"56fc813f",
X"7655ab39",
X"79841b71",
X"08943d70",
X"5b5b525b",
X"56758025",
X"8c387530",
X"56ad7834",
X"0280c105",
X"57765480",
X"538a5275",
X"51fbd53f",
X"77557e54",
X"b839913d",
X"70557780",
X"d8327030",
X"70802556",
X"51585690",
X"5279841b",
X"7108535b",
X"57fbb13f",
X"7555db39",
X"79841b83",
X"1233545b",
X"56983979",
X"841b7108",
X"575b5680",
X"547f537c",
X"527d51fc",
X"9c3f8739",
X"76527d51",
X"7c2d6670",
X"33588105",
X"47fd8339",
X"943d0d04",
X"7283c094",
X"0c7183c0",
X"980c04fb",
X"3d0d883d",
X"70708405",
X"52085754",
X"755383c0",
X"94085283",
X"c0980851",
X"fcc63f87",
X"3d0d04ff",
X"3d0d7370",
X"08535102",
X"93053372",
X"34700881",
X"05710c83",
X"3d0d04fc",
X"3d0d873d",
X"88115578",
X"54bdbb53",
X"51fc993f",
X"8052873d",
X"51d13f86",
X"3d0d04fc",
X"3d0d7655",
X"7483c3ac",
X"082eaf38",
X"80537451",
X"87c13f83",
X"c0800881",
X"ff06ff14",
X"7081ff06",
X"7230709f",
X"2a515255",
X"53547280",
X"2e843871",
X"dd3873fe",
X"387483c3",
X"ac0c863d",
X"0d04ff3d",
X"0dff0b83",
X"c3ac0c84",
X"a53f8151",
X"87853f83",
X"c0800881",
X"ff065271",
X"ee3881d3",
X"3f7183c0",
X"800c833d",
X"0d04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"823f7280",
X"2ea03883",
X"c3c01433",
X"75708105",
X"57348114",
X"7083ffff",
X"06ff1570",
X"83ffff06",
X"56525552",
X"dd39800b",
X"83c0800c",
X"863d0d04",
X"fc3d0d76",
X"787a1156",
X"53558053",
X"71742e93",
X"38721551",
X"703383c3",
X"c0133481",
X"12811454",
X"52ea3980",
X"0b83c080",
X"0c863d0d",
X"04fd3d0d",
X"905483c3",
X"ac085186",
X"f43f83c0",
X"800881ff",
X"06ff1571",
X"30713070",
X"73079f2a",
X"729f2a06",
X"52555255",
X"5372db38",
X"853d0d04",
X"803d0d83",
X"c3b80810",
X"83c3b008",
X"079080a8",
X"0c823d0d",
X"04800b83",
X"c3b80ce4",
X"3f04810b",
X"83c3b80c",
X"db3f04ed",
X"3f047183",
X"c3b40c04",
X"803d0d80",
X"51f43f81",
X"0b83c3b8",
X"0c810b83",
X"c3b00cff",
X"bb3f823d",
X"0d04803d",
X"0d723070",
X"74078025",
X"83c3b00c",
X"51ffa53f",
X"823d0d04",
X"803d0d02",
X"8b053390",
X"80a40c90",
X"80a80870",
X"81065151",
X"70f53890",
X"80a40870",
X"81ff0683",
X"c0800c51",
X"823d0d04",
X"803d0d81",
X"ff51d13f",
X"83c08008",
X"81ff0683",
X"c0800c82",
X"3d0d0480",
X"3d0d7390",
X"2b730790",
X"80b40c82",
X"3d0d0404",
X"fb3d0d78",
X"0284059f",
X"05337098",
X"2b555755",
X"7280259b",
X"387580ff",
X"06568052",
X"80f751e0",
X"3f83c080",
X"0881ff06",
X"54738126",
X"80ff3880",
X"51fee73f",
X"ffa23f81",
X"51fedf3f",
X"ff9a3f75",
X"51feed3f",
X"74982a51",
X"fee63f74",
X"902a7081",
X"ff065253",
X"feda3f74",
X"882a7081",
X"ff065253",
X"fece3f74",
X"81ff0651",
X"fec63f81",
X"557580c0",
X"2e098106",
X"86388195",
X"558d3975",
X"80c82e09",
X"81068438",
X"81875574",
X"51fea53f",
X"8a55fec8",
X"3f83c080",
X"0881ff06",
X"70982b54",
X"54728025",
X"8c38ff15",
X"7081ff06",
X"565374e2",
X"387383c0",
X"800c873d",
X"0d04fa3d",
X"0dfdc53f",
X"8051fdda",
X"3f8a54fe",
X"933fff14",
X"7081ff06",
X"555373f3",
X"38737453",
X"5580c051",
X"fea63f83",
X"c0800881",
X"ff065473",
X"812e0981",
X"06829f38",
X"83aa5280",
X"c851fe8c",
X"3f83c080",
X"0881ff06",
X"5372812e",
X"09810681",
X"a8387454",
X"873d7411",
X"5456fdc8",
X"3f83c080",
X"08733481",
X"147081ff",
X"06555383",
X"7427e538",
X"029a0533",
X"5372812e",
X"09810681",
X"d938029b",
X"05335380",
X"ce905472",
X"81aa2e8d",
X"3881c739",
X"80e4518b",
X"9a3fff14",
X"5473802e",
X"81b83882",
X"0a5281e9",
X"51fda53f",
X"83c08008",
X"81ff0653",
X"72de3872",
X"5280fa51",
X"fd923f83",
X"c0800881",
X"ff065372",
X"81903872",
X"54731653",
X"fcd63f83",
X"c0800873",
X"34811470",
X"81ff0655",
X"53837427",
X"e838873d",
X"3370862a",
X"70810651",
X"54548c55",
X"7280e338",
X"845580de",
X"39745281",
X"e951fccc",
X"3f83c080",
X"0881ff06",
X"53825581",
X"e9568173",
X"27863873",
X"5580c156",
X"80ce9054",
X"8a3980e4",
X"518a8c3f",
X"ff145473",
X"802ea938",
X"80527551",
X"fc9a3f83",
X"c0800881",
X"ff065372",
X"e1388480",
X"5280d051",
X"fc863f83",
X"c0800881",
X"ff065372",
X"802e8338",
X"80557483",
X"c3bc3480",
X"51fb873f",
X"fbc23f88",
X"3d0d04fb",
X"3d0d7754",
X"800b83c3",
X"bc337083",
X"2a708106",
X"51555755",
X"72752e09",
X"81068538",
X"73892b54",
X"735280d1",
X"51fbbd3f",
X"83c08008",
X"81ff0653",
X"72bd3882",
X"b8c054fb",
X"833f83c0",
X"800881ff",
X"06537281",
X"ff2e0981",
X"068938ff",
X"145473e7",
X"389f3972",
X"81fe2e09",
X"81069638",
X"83c7c052",
X"83c3c051",
X"faed3ffa",
X"d33ffad0",
X"3f833981",
X"558051fa",
X"893ffac4",
X"3f7481ff",
X"0683c080",
X"0c873d0d",
X"04fb3d0d",
X"7783c3c0",
X"56548151",
X"f9ec3f83",
X"c3bc3370",
X"832a7081",
X"06515456",
X"72853873",
X"892b5473",
X"5280d851",
X"fab63f83",
X"c0800881",
X"ff065372",
X"80e43881",
X"ff51f9d4",
X"3f81fe51",
X"f9ce3f84",
X"80537470",
X"81055633",
X"51f9c13f",
X"ff137083",
X"ffff0651",
X"5372eb38",
X"7251f9b0",
X"3f7251f9",
X"ab3ff9d0",
X"3f83c080",
X"089f0653",
X"a7885472",
X"852e8c38",
X"993980e4",
X"5187c43f",
X"ff1454f9",
X"b33f83c0",
X"800881ff",
X"2e843873",
X"e9388051",
X"f8e43ff9",
X"9f3f800b",
X"83c0800c",
X"873d0d04",
X"7183c7c4",
X"0c888080",
X"0b83c7c0",
X"0c848080",
X"0b83c7c8",
X"0c04fd3d",
X"0d777017",
X"557705ff",
X"1a535371",
X"ff2e9438",
X"73708105",
X"55335170",
X"73708105",
X"5534ff12",
X"52e93985",
X"3d0d04fb",
X"3d0d87a6",
X"810b83c7",
X"c4085656",
X"753383a6",
X"801634a0",
X"5483a080",
X"5383c7c4",
X"085283c7",
X"c00851ff",
X"b13fa054",
X"83a48053",
X"83c7c408",
X"5283c7c0",
X"0851ff9e",
X"3f905483",
X"a8805383",
X"c7c40852",
X"83c7c008",
X"51ff8b3f",
X"a0538052",
X"83c7c808",
X"83a08005",
X"5186953f",
X"a0538052",
X"83c7c808",
X"83a48005",
X"5186853f",
X"90538052",
X"83c7c808",
X"83a88005",
X"5185f53f",
X"ff763483",
X"a0805480",
X"5383c7c4",
X"085283c7",
X"c80851fe",
X"c53f80d0",
X"805483b0",
X"805383c7",
X"c4085283",
X"c7c80851",
X"feb03f87",
X"ba3fa254",
X"805383c7",
X"c8088c80",
X"055281df",
X"c451fe9a",
X"3f860b87",
X"a8833480",
X"0b87a882",
X"34800b87",
X"a09a34af",
X"0b87a096",
X"34bf0b87",
X"a0973480",
X"0b87a098",
X"349f0b87",
X"a0993480",
X"0b87a09b",
X"34e00b87",
X"a88934a2",
X"0b87a880",
X"34830b87",
X"a48f3482",
X"0b87a881",
X"34873d0d",
X"04fc3d0d",
X"83a08054",
X"805383c7",
X"c8085283",
X"c7c40851",
X"fdb83f80",
X"d0805483",
X"b0805383",
X"c7c80852",
X"83c7c408",
X"51fda33f",
X"a05483a0",
X"805383c7",
X"c8085283",
X"c7c40851",
X"fd903fa0",
X"5483a480",
X"5383c7c8",
X"085283c7",
X"c40851fc",
X"fd3f9054",
X"83a88053",
X"83c7c808",
X"5283c7c4",
X"0851fcea",
X"3f83c7c4",
X"085583a6",
X"80153387",
X"a6813486",
X"3d0d04fa",
X"3d0d7870",
X"5255c1df",
X"3f83ffff",
X"0b83c080",
X"0825a938",
X"7451c1e0",
X"3f83c080",
X"089e3883",
X"c0800857",
X"883dfc05",
X"54848080",
X"5383c7c4",
X"08527451",
X"ffbf993f",
X"ffbedf3f",
X"883d0d04",
X"fa3d0d78",
X"705255c1",
X"9e3f83ff",
X"ff0b83c0",
X"80082596",
X"38805788",
X"3dfc0554",
X"84808053",
X"83c7c408",
X"527451c0",
X"913f883d",
X"0d04803d",
X"0d908090",
X"08810683",
X"c0800c82",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe067607",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"812c8106",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fd06",
X"76100772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087082",
X"2cbf0683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fe8306",
X"76822b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"882c8706",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f1ff",
X"0676882b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70912cbf",
X"0683c080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870fc",
X"87ffff06",
X"76912b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"992c8106",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870ffbf",
X"0a067699",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908080",
X"0870882c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"80087089",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8a2c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708b2c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708c2c",
X"bf0683c0",
X"800c5182",
X"3d0d04fe",
X"3d0d7481",
X"e629872a",
X"9080a00c",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d848080",
X"53805288",
X"800a51ff",
X"b33f8180",
X"80538052",
X"82800a51",
X"c63f843d",
X"0d04803d",
X"0d8151fc",
X"aa3f7280",
X"2e903880",
X"51fdfe3f",
X"cd3f83c7",
X"cc3351fd",
X"f43f8151",
X"fcbb3f80",
X"51fcb63f",
X"8051fc87",
X"3f823d0d",
X"04fd3d0d",
X"75528054",
X"80ff7225",
X"8838810b",
X"ff801353",
X"54ffbf12",
X"51709926",
X"8638e012",
X"52b039ff",
X"9f125199",
X"7127a738",
X"d012e013",
X"54517089",
X"26853872",
X"52983972",
X"8f268538",
X"72528f39",
X"71ba2e09",
X"81068538",
X"9a528339",
X"80527380",
X"2e853881",
X"80125271",
X"81ff0683",
X"c0800c85",
X"3d0d0480",
X"3d0d84d8",
X"c0518071",
X"70810553",
X"347084e0",
X"c02e0981",
X"06f03882",
X"3d0d04fe",
X"3d0d0297",
X"053351fe",
X"f43f83c0",
X"800881ff",
X"0683c7d0",
X"08545280",
X"73249b38",
X"83c88008",
X"137283c8",
X"84080753",
X"53717334",
X"83c7d008",
X"810583c7",
X"d00c843d",
X"0d04fa3d",
X"0d82800a",
X"1b558057",
X"883dfc05",
X"54795374",
X"527851ff",
X"baa83f88",
X"3d0d04fe",
X"3d0d83c7",
X"e8085274",
X"51c18c3f",
X"83c08008",
X"8c387653",
X"755283c7",
X"e80851c6",
X"3f843d0d",
X"04fe3d0d",
X"83c7e808",
X"53755274",
X"51ffbbca",
X"3f83c080",
X"088d3877",
X"53765283",
X"c7e80851",
X"ffa03f84",
X"3d0d04fe",
X"3d0d83c7",
X"e80851ff",
X"babd3f83",
X"c0800881",
X"80802e09",
X"81068838",
X"83c18080",
X"539c3983",
X"c7e80851",
X"ffbaa03f",
X"83c08008",
X"80d0802e",
X"09810693",
X"3883c1b0",
X"805383c0",
X"80085283",
X"c7e80851",
X"fed43f84",
X"3d0d0480",
X"3d0df9fc",
X"3f83c080",
X"08842981",
X"dfe80570",
X"0883c080",
X"0c51823d",
X"0d04ed3d",
X"0d804480",
X"43804280",
X"4180705a",
X"5bfdcc3f",
X"800b83c7",
X"d00c800b",
X"83c8840c",
X"81dcbc51",
X"e9c53f81",
X"800b83c8",
X"840c81dc",
X"c051e9b7",
X"3f80d00b",
X"83c7d00c",
X"7830707a",
X"07802570",
X"872b83c8",
X"840c5155",
X"f8ed3f83",
X"c0800852",
X"81dcc851",
X"e9913f80",
X"f80b83c7",
X"d00c7881",
X"32703070",
X"72078025",
X"70872b83",
X"c8840c51",
X"56569e9c",
X"3f83c080",
X"085281dc",
X"d851e8e7",
X"3f81a00b",
X"83c7d00c",
X"78823270",
X"30707207",
X"80257087",
X"2b83c884",
X"0c515656",
X"fec53f83",
X"c0800852",
X"81dce851",
X"e8bd3f81",
X"c80b83c7",
X"d00c7883",
X"32703070",
X"72078025",
X"70872b83",
X"c8840c51",
X"5683c7e8",
X"085256ff",
X"b59b3f83",
X"c0800852",
X"81dcf051",
X"e88d3f82",
X"980b83c7",
X"d00c810b",
X"83c7d45b",
X"5883c7d0",
X"0883197a",
X"32703070",
X"72078025",
X"70872b83",
X"c8840c51",
X"578e3d70",
X"55ff1b54",
X"5757579b",
X"de3f7970",
X"84055b08",
X"51ffb4d1",
X"3f745483",
X"c0800853",
X"775281dc",
X"f851e7bf",
X"3fa81783",
X"c7d00c81",
X"18587785",
X"2e098106",
X"ffaf3883",
X"b80b83c7",
X"d00c7888",
X"32703070",
X"72078025",
X"70872b83",
X"c8840c51",
X"5656f7b9",
X"3f81dd88",
X"5583c080",
X"08802e8f",
X"3883c7e4",
X"0851ffb3",
X"fc3f83c0",
X"80085574",
X"5281dd90",
X"51e6ec3f",
X"84880b83",
X"c7d00c78",
X"89327030",
X"70720780",
X"2570872b",
X"83c8840c",
X"515681dd",
X"9c5256e6",
X"ca3f84b0",
X"0b83c7d0",
X"0c788a32",
X"70307072",
X"07802570",
X"872b83c8",
X"840c5156",
X"81dda852",
X"56e6a83f",
X"85800b83",
X"c7d00c78",
X"8b327030",
X"70720780",
X"2570872b",
X"83c8840c",
X"515681dd",
X"c45256e6",
X"863f868d",
X"a051f7ef",
X"3f805291",
X"3d705255",
X"9ed53f83",
X"5274519e",
X"ce3f6355",
X"7483e038",
X"61195978",
X"80258538",
X"74599039",
X"8b792585",
X"388b5987",
X"39788b26",
X"83bf3878",
X"822b5581",
X"d7b41508",
X"04f5903f",
X"83c08008",
X"61575575",
X"812e0981",
X"06893883",
X"c0800810",
X"55903975",
X"ff2e0981",
X"06883883",
X"c0800881",
X"2c559075",
X"25853890",
X"55883974",
X"80248338",
X"81557451",
X"f4ea3f82",
X"f4399a9f",
X"3f83c080",
X"08610555",
X"74802585",
X"38805588",
X"39877525",
X"83388755",
X"74518e82",
X"3f82d239",
X"f4da3f83",
X"c0800861",
X"05557480",
X"25853880",
X"55883986",
X"75258338",
X"86557451",
X"f4d33f82",
X"b0396087",
X"3862802e",
X"82a73883",
X"c39c0883",
X"c3980cad",
X"e50b83c3",
X"a00c83c7",
X"e80851d5",
X"9a3ff9cb",
X"3f828a39",
X"60568076",
X"259838ad",
X"840b83c3",
X"a00c83c7",
X"c4157008",
X"5255d4fb",
X"3f740852",
X"92397580",
X"25923883",
X"c7c41508",
X"51ffb0ff",
X"3f8052fc",
X"1951b839",
X"62802e81",
X"d03883c7",
X"c4157008",
X"83c7d408",
X"720c83c7",
X"d40cfc1a",
X"70535155",
X"8ccf3f83",
X"c0800856",
X"80518cc5",
X"3f83c080",
X"08527451",
X"88de3f75",
X"52805188",
X"d73f8199",
X"39605580",
X"7525b838",
X"83c3a808",
X"83c3980c",
X"ade50b83",
X"c3a00c83",
X"c7e40851",
X"d4853f83",
X"c7e40851",
X"d1a63f83",
X"c0800881",
X"ff067052",
X"55f3b33f",
X"74802e80",
X"e0388155",
X"80e33974",
X"802580d5",
X"3883c7e4",
X"0851ffaf",
X"ee3f8051",
X"f3943f80",
X"c4396280",
X"2ebf3883",
X"c3a40883",
X"c3980cad",
X"e50b83c3",
X"a00c83c7",
X"ec0851d3",
X"b23f7889",
X"2e098106",
X"8b3883c7",
X"ec0851f0",
X"f73f9639",
X"788a2e09",
X"81068e38",
X"83c7ec08",
X"51f0a43f",
X"84396287",
X"387a802e",
X"f8af3880",
X"557483c0",
X"800c953d",
X"0d04fe3d",
X"0d83c7f0",
X"5180f48e",
X"3ff2f73f",
X"83c08008",
X"802e8638",
X"8051818a",
X"39f2fc3f",
X"83c08008",
X"80fe38f3",
X"9c3f83c0",
X"8008802e",
X"b9388151",
X"f0d93f80",
X"51f2b23f",
X"ecd13f80",
X"0b83c7d0",
X"0cf7cf3f",
X"83c08008",
X"53ff0b83",
X"c7d00cee",
X"c43f7280",
X"cb3883c7",
X"cc3351f2",
X"8c3f7251",
X"f0a93f80",
X"c039f2c4",
X"3f83c080",
X"08802eb5",
X"388151f0",
X"963f8051",
X"f1ef3fec",
X"8e3fad84",
X"0b83c3a0",
X"0c83c7d4",
X"0851d1eb",
X"3fff0b83",
X"c7d00cee",
X"803f83c7",
X"d4085280",
X"5186893f",
X"8151f3b6",
X"3f843d0d",
X"04fb3d0d",
X"805283c7",
X"f05180e3",
X"9d3f800b",
X"83c7cc34",
X"90808052",
X"86848080",
X"51ffb1d4",
X"3f83c080",
X"08819738",
X"89e43f81",
X"e28851ff",
X"b6933f83",
X"c0800855",
X"9c800a54",
X"80c08053",
X"81ddcc52",
X"83c08008",
X"51f5923f",
X"83c7e808",
X"5381dddc",
X"527451ff",
X"b0dc3f83",
X"c0800884",
X"38f5a03f",
X"83c7ec08",
X"5381dde8",
X"527451ff",
X"b0c43f83",
X"c08008b6",
X"38873dfc",
X"05548480",
X"805386a8",
X"80805283",
X"c7ec0851",
X"ffaecf3f",
X"83c08008",
X"93387584",
X"80802e09",
X"81068938",
X"810b83c7",
X"cc348739",
X"800b83c7",
X"cc3483c7",
X"cc3351f0",
X"8c3f8151",
X"f1f83f93",
X"953f8151",
X"f1f03f81",
X"51fd8f3f",
X"fa3983c0",
X"8c080283",
X"c08c0cfb",
X"3d0d0281",
X"ddf40b83",
X"c39c0c81",
X"ddf80b83",
X"c3940c81",
X"ddfc0b83",
X"c3a80c81",
X"de800b83",
X"c3a40c83",
X"c08c08fc",
X"050c800b",
X"83c7d40b",
X"83c08c08",
X"f8050c83",
X"c08c08f4",
X"050cffae",
X"d73f83c0",
X"80088605",
X"fc0683c0",
X"8c08f005",
X"0c0283c0",
X"8c08f005",
X"08310d83",
X"3d7083c0",
X"8c08f805",
X"08708405",
X"83c08c08",
X"f8050c0c",
X"51ffab9f",
X"3f83c08c",
X"08f40508",
X"810583c0",
X"8c08f405",
X"0c83c08c",
X"08f40508",
X"872e0981",
X"06ffab38",
X"86948080",
X"51e8b53f",
X"ff0b83c7",
X"d00c800b",
X"83c8840c",
X"84d8c00b",
X"83c8800c",
X"8151ecdb",
X"3f8151ed",
X"803f8051",
X"ecfb3f81",
X"51eda13f",
X"8251edc9",
X"3f8051ed",
X"f13f8051",
X"ee9b3f80",
X"d1ab5280",
X"51dd993f",
X"fccf3f83",
X"c08c08fc",
X"05080d80",
X"0b83c080",
X"0c873d0d",
X"83c08c0c",
X"04803d0d",
X"81ff5180",
X"0b83c894",
X"1234ff11",
X"5170f438",
X"823d0d04",
X"ff3d0d73",
X"70335351",
X"81113371",
X"34718112",
X"34833d0d",
X"04fb3d0d",
X"77795656",
X"80707155",
X"55527175",
X"25ac3872",
X"16703370",
X"147081ff",
X"06555151",
X"51717427",
X"89388112",
X"7081ff06",
X"53517181",
X"147083ff",
X"ff065552",
X"54747324",
X"d6387183",
X"c0800c87",
X"3d0d04fb",
X"3d0d7756",
X"d4e33f83",
X"c0800880",
X"2ef63883",
X"cab00886",
X"057081ff",
X"065253d2",
X"e53f810b",
X"9088d434",
X"9088d433",
X"7081ff06",
X"5153728b",
X"38f9e73f",
X"8351edcf",
X"3fea3980",
X"55741675",
X"822b5454",
X"9088c013",
X"33743481",
X"15557485",
X"2e098106",
X"e838810b",
X"9088d434",
X"753383c8",
X"94348116",
X"3383c895",
X"34821633",
X"83c89634",
X"83163383",
X"c8973484",
X"5283c894",
X"51feba3f",
X"83c08008",
X"81ff0684",
X"17335753",
X"72762e09",
X"81068c38",
X"d38c3f83",
X"c0800880",
X"2e9c3883",
X"cab008a8",
X"2e098106",
X"8b3883ca",
X"c80883ca",
X"b00c8739",
X"a80b83ca",
X"b00c80e4",
X"51ecc83f",
X"873d0d04",
X"f43d0d7e",
X"60595580",
X"5d807582",
X"2b7183ca",
X"b4120c83",
X"cacc175b",
X"5b577679",
X"3477772e",
X"83b73876",
X"527751ff",
X"a9e83f8e",
X"3dfc0554",
X"905383ca",
X"9c527751",
X"ffa9a33f",
X"7c567590",
X"2e098106",
X"83933883",
X"ca9c51fd",
X"933f83ca",
X"9e51fd8c",
X"3f83caa0",
X"51fd853f",
X"7683caac",
X"0c7751ff",
X"a6ef3f81",
X"dbcc5283",
X"c0800851",
X"c9883f83",
X"c0800881",
X"2e098106",
X"80d43876",
X"83cac40c",
X"820b83ca",
X"9c34ff96",
X"0b83ca9d",
X"347751ff",
X"a9b53f83",
X"c0800855",
X"83c08008",
X"77258838",
X"83c08008",
X"8f055574",
X"842c7083",
X"ffff0670",
X"882a5851",
X"557583ca",
X"9e347483",
X"ca9f3476",
X"83caa034",
X"ff800b83",
X"caa13481",
X"903983ca",
X"9c3383ca",
X"9d337188",
X"2b07565b",
X"7483ffff",
X"2e098106",
X"80e838fe",
X"800b83ca",
X"c40c810b",
X"83caac0c",
X"ff0b83ca",
X"9c34ff0b",
X"83ca9d34",
X"7751ffa8",
X"c23f83c0",
X"800883ca",
X"d00c83c0",
X"80085583",
X"c0800880",
X"25883883",
X"c080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583ca9e",
X"347483ca",
X"9f347683",
X"caa034ff",
X"800b83ca",
X"a134810b",
X"83caab34",
X"a5397485",
X"962e0981",
X"0680fe38",
X"7583cac4",
X"0c7751ff",
X"a7f63f83",
X"caab3383",
X"c0800807",
X"557483ca",
X"ab3483ca",
X"ab338106",
X"5574802e",
X"83388457",
X"83caa033",
X"83caa133",
X"71882b07",
X"565c7481",
X"802e0981",
X"06a13883",
X"ca9e3383",
X"ca9f3371",
X"882b0756",
X"5bad8075",
X"27873876",
X"8207579c",
X"39768107",
X"57963974",
X"82802e09",
X"81068738",
X"76830757",
X"87397481",
X"ff268a38",
X"7783cab4",
X"1b0c7679",
X"348e3d0d",
X"04803d0d",
X"72842983",
X"cab40570",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d727083",
X"c88c0c70",
X"842981e1",
X"bc057008",
X"83cac80c",
X"5151823d",
X"0d04fe3d",
X"0d8151de",
X"3f800b83",
X"ca980c80",
X"0b83ca94",
X"0cff0b83",
X"c8900ca8",
X"0b83cab0",
X"0cae51cd",
X"8d3f800b",
X"83cab454",
X"52807370",
X"8405550c",
X"81125271",
X"842e0981",
X"06ef3884",
X"3d0d04fe",
X"3d0d7402",
X"84059605",
X"22535371",
X"802e9638",
X"72708105",
X"543351cd",
X"983fff12",
X"7083ffff",
X"065152e7",
X"39843d0d",
X"04fe3d0d",
X"02920522",
X"5382ac51",
X"e7bd3f80",
X"c351ccf5",
X"3f819651",
X"e7b13f72",
X"5283c894",
X"51ffb43f",
X"725283c8",
X"9451f8d1",
X"3f83c080",
X"0881ff06",
X"51ccd23f",
X"843d0d04",
X"ffb13d0d",
X"80d13df8",
X"0551f8fb",
X"3f83ca98",
X"08810583",
X"ca980c80",
X"cf3d33cf",
X"117081ff",
X"06515656",
X"74832688",
X"e638758f",
X"06ff0556",
X"7583c890",
X"082e9b38",
X"75832696",
X"387583c8",
X"900c7584",
X"2983cab4",
X"05700853",
X"557551f9",
X"fb3f8076",
X"2488c238",
X"75842983",
X"cab40555",
X"7408802e",
X"88b33883",
X"c8900884",
X"2983cab4",
X"05700802",
X"880582b9",
X"0533525b",
X"557480d2",
X"2e84b038",
X"7480d224",
X"903874bf",
X"2e9c3874",
X"80d02e81",
X"d53887f2",
X"397480d3",
X"2e80d338",
X"7480d72e",
X"81c43887",
X"e1390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290556",
X"56cbce3f",
X"80c151cb",
X"883ff6cd",
X"3f83cacb",
X"3383c894",
X"34815283",
X"c89451cc",
X"a93f8151",
X"fde73f74",
X"8b3883ca",
X"c80883ca",
X"b00c8739",
X"a80b83ca",
X"b00ccb99",
X"3f80c151",
X"cad33ff6",
X"983f900b",
X"83caab33",
X"81065656",
X"74802e83",
X"38985683",
X"caa03383",
X"caa13371",
X"882b0756",
X"59748180",
X"2e098106",
X"9c3883ca",
X"9e3383ca",
X"9f337188",
X"2b075657",
X"ad807527",
X"8c387581",
X"80075685",
X"3975a007",
X"567583c8",
X"9434ff0b",
X"83c89534",
X"e00b83c8",
X"9634800b",
X"83c89734",
X"845283c8",
X"9451cb9e",
X"3f845186",
X"9b390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290556",
X"59ca8e3f",
X"7951ffa2",
X"a33f83c0",
X"8008802e",
X"8a3880ce",
X"51c9ba3f",
X"85f13980",
X"c151c9b1",
X"3fcaa63f",
X"c8db3f83",
X"cac40858",
X"8375259b",
X"3883caa0",
X"3383caa1",
X"3371882b",
X"07fc1771",
X"297a0583",
X"80055a51",
X"578d3974",
X"81802918",
X"ff800558",
X"81805780",
X"5676762e",
X"9238c98d",
X"3f83c080",
X"0883c894",
X"17348116",
X"56eb39c8",
X"fc3f83c0",
X"800881ff",
X"06775383",
X"c8945256",
X"f4c33f83",
X"c0800881",
X"ff065575",
X"752e0981",
X"06819538",
X"9451e2fb",
X"3fc8f63f",
X"80c151c8",
X"b03fc9a5",
X"3f775279",
X"51ffa0b6",
X"3f805e80",
X"d13dfdf4",
X"05547653",
X"83c89452",
X"7951ff9e",
X"c33f0282",
X"b9053355",
X"81597480",
X"d72e0981",
X"0680c538",
X"77527951",
X"ffa0873f",
X"80d13dfd",
X"f0055476",
X"538f3d70",
X"537a5258",
X"ff9fbf3f",
X"80567676",
X"2ea23875",
X"1883c894",
X"17337133",
X"70723270",
X"30708025",
X"70307f06",
X"811d5d5f",
X"51515152",
X"5b55db39",
X"82ac51e1",
X"f63f7880",
X"2e863880",
X"c3518439",
X"80ce51c7",
X"a43fc899",
X"3fc6ce3f",
X"83d83902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"59558070",
X"5d5980e4",
X"51e1c03f",
X"c7bb3f80",
X"c151c6f5",
X"3f83caac",
X"08792e82",
X"d63883ca",
X"d00880fc",
X"055580fd",
X"52745185",
X"c13f83c0",
X"80085b77",
X"8224b238",
X"ff187087",
X"2b83ffff",
X"800681e0",
X"880583c8",
X"94595755",
X"81805575",
X"70810557",
X"33777081",
X"055934ff",
X"157081ff",
X"06515574",
X"ea388285",
X"397782e8",
X"2e81a338",
X"7782e92e",
X"09810681",
X"aa387858",
X"77873270",
X"30707207",
X"80257a8a",
X"32703070",
X"72078025",
X"73075354",
X"5a515755",
X"75802e97",
X"38787826",
X"9238a00b",
X"83c8941a",
X"34811970",
X"81ff065a",
X"55eb3981",
X"187081ff",
X"0659558a",
X"7827ffbc",
X"388f5883",
X"c88f1833",
X"83c89419",
X"34ff1870",
X"81ff0659",
X"55778426",
X"ea389058",
X"800b83c8",
X"94193481",
X"187081ff",
X"0670982b",
X"52595574",
X"8025e938",
X"80c6557a",
X"858f2484",
X"3880c255",
X"7483c894",
X"3480f10b",
X"83c89734",
X"810b83c8",
X"98347a83",
X"c895347a",
X"882c5574",
X"83c89634",
X"80cb3982",
X"f0782580",
X"c4387780",
X"fd29fd97",
X"d3055279",
X"51ff9ce2",
X"3f80d13d",
X"fdec0554",
X"80fd5383",
X"c8945279",
X"51ff9c9a",
X"3f7b8119",
X"59567580",
X"fc248338",
X"78587788",
X"2c557483",
X"c9913477",
X"83c99234",
X"7583c993",
X"34818059",
X"80cc3983",
X"cac40857",
X"8378259b",
X"3883caa0",
X"3383caa1",
X"3371882b",
X"07fc1a71",
X"29790583",
X"80055951",
X"598d3977",
X"81802917",
X"ff800557",
X"81805976",
X"527951ff",
X"9bf03f80",
X"d13dfdec",
X"05547853",
X"83c89452",
X"7951ff9b",
X"a93f7851",
X"f6bf3fc4",
X"bc3fc2f1",
X"3f8b3983",
X"ca940881",
X"0583ca94",
X"0c80d13d",
X"0d04f6e0",
X"3ffc39fc",
X"3d0d7678",
X"71842983",
X"cab40570",
X"08515353",
X"53709e38",
X"80ce7234",
X"80cf0b81",
X"133480ce",
X"0b821334",
X"80c50b83",
X"13347084",
X"133480e7",
X"3983cacc",
X"13335480",
X"d2723473",
X"822a7081",
X"06515180",
X"cf537084",
X"3880d753",
X"72811334",
X"a00b8213",
X"34738306",
X"5170812e",
X"9e387081",
X"24883870",
X"802e8f38",
X"9f397082",
X"2e923870",
X"832e9238",
X"933980d8",
X"558e3980",
X"d3558939",
X"80cd5584",
X"3980c455",
X"74831334",
X"80c40b84",
X"1334800b",
X"85133486",
X"3d0d0483",
X"c88c0883",
X"c0800c04",
X"803d0d83",
X"c88c0884",
X"2981e1dc",
X"05700883",
X"c0800c51",
X"823d0d04",
X"fc3d0d76",
X"78535481",
X"53805587",
X"39711073",
X"10545273",
X"72265172",
X"802ea738",
X"70802e86",
X"38718025",
X"e8387280",
X"2e983871",
X"74268938",
X"73723175",
X"74075654",
X"72812a72",
X"812a5353",
X"e5397351",
X"78833874",
X"517083c0",
X"800c863d",
X"0d04fe3d",
X"0d805375",
X"527451ff",
X"a33f843d",
X"0d04fe3d",
X"0d815375",
X"527451ff",
X"933f843d",
X"0d04fb3d",
X"0d777955",
X"55805674",
X"76258638",
X"74305581",
X"56738025",
X"88387330",
X"76813257",
X"54805373",
X"527451fe",
X"e73f83c0",
X"80085475",
X"802e8738",
X"83c08008",
X"30547383",
X"c0800c87",
X"3d0d04fa",
X"3d0d787a",
X"57558057",
X"74772586",
X"38743055",
X"8157759f",
X"2c548153",
X"75743274",
X"31527451",
X"feaa3f83",
X"c0800854",
X"76802e87",
X"3883c080",
X"08305473",
X"83c0800c",
X"883d0d04",
X"fc3d0d76",
X"5580750c",
X"800b8416",
X"0c800b88",
X"160c800b",
X"8c160c83",
X"c7f05180",
X"dacc3f87",
X"a6803370",
X"81ff0651",
X"52d9ff3f",
X"71812a81",
X"32728132",
X"71810671",
X"81063184",
X"180c5454",
X"71832a81",
X"3272822a",
X"81327181",
X"06718106",
X"31770c53",
X"5387a090",
X"33700981",
X"0688170c",
X"5283c080",
X"08802e80",
X"c23883c0",
X"8008812a",
X"70810683",
X"c0800881",
X"06318417",
X"0c5283c0",
X"8008832a",
X"83c08008",
X"822a7181",
X"06718106",
X"31770c53",
X"5383c080",
X"08842a81",
X"0688160c",
X"83c08008",
X"852a8106",
X"8c160c86",
X"3d0d04fe",
X"3d0d7476",
X"54527151",
X"fec63f72",
X"812ea238",
X"8173268d",
X"3872822e",
X"a8387283",
X"2e9c38e6",
X"397108e2",
X"38841208",
X"dd388812",
X"08d838a5",
X"39881208",
X"812e9e38",
X"91398812",
X"08812e95",
X"38710891",
X"38841208",
X"8c388c12",
X"08812e09",
X"8106ffb2",
X"38843d0d",
X"04fb3d0d",
X"78028405",
X"9f053355",
X"56800b81",
X"d9d05653",
X"81732b74",
X"06527180",
X"2e833881",
X"52747082",
X"05562270",
X"73902b07",
X"90809c0c",
X"51811353",
X"72882e09",
X"8106d938",
X"805383ca",
X"d8133351",
X"7081ff2e",
X"b2387010",
X"81d7f005",
X"70225551",
X"80731770",
X"33701081",
X"d7f00570",
X"22515151",
X"52527371",
X"2e913881",
X"12527186",
X"2e098106",
X"f1387390",
X"809c0c81",
X"13537286",
X"2e098106",
X"ffb83880",
X"53721670",
X"33515170",
X"81ff2e94",
X"38701081",
X"d7f00570",
X"22708480",
X"80079080",
X"9c0c5151",
X"81135372",
X"862e0981",
X"06d73880",
X"53721651",
X"703383ca",
X"d8143481",
X"13537286",
X"2e098106",
X"ec38873d",
X"0d0404ff",
X"3d0d7402",
X"84058f05",
X"33525270",
X"88387190",
X"80940c8e",
X"3970812e",
X"09810686",
X"38719080",
X"980c833d",
X"0d04fb3d",
X"0d029f05",
X"3379982b",
X"70982c7c",
X"982b7098",
X"2c83caf4",
X"15703370",
X"982b7098",
X"2c51585c",
X"5a515551",
X"54547073",
X"2e098106",
X"943883ca",
X"d4143370",
X"982b7098",
X"2c515256",
X"70722eb1",
X"38727534",
X"7183cad4",
X"153483ca",
X"d53383ca",
X"f5337198",
X"2b71902b",
X"0783cad4",
X"3370882b",
X"720783ca",
X"f4337107",
X"9080b80c",
X"52595354",
X"52873d0d",
X"04fe3d0d",
X"74811133",
X"71337188",
X"2b0783c0",
X"800c5351",
X"843d0d04",
X"83cae033",
X"83c0800c",
X"04f53d0d",
X"02bb0533",
X"028405bf",
X"05330288",
X"0580c305",
X"33028c05",
X"80c60522",
X"665c5a5e",
X"5c567a55",
X"7b548953",
X"a1527d51",
X"80d0c03f",
X"83c08008",
X"81ff0683",
X"c0800c8d",
X"3d0d0483",
X"c08c0802",
X"83c08c0c",
X"f53d0d83",
X"c08c0888",
X"050883c0",
X"8c088f05",
X"3383c08c",
X"08920522",
X"028c0573",
X"900583c0",
X"8c08e805",
X"0c83c08c",
X"08f8050c",
X"83c08c08",
X"f0050c83",
X"c08c08ec",
X"050c83c0",
X"8c08f405",
X"0c800b83",
X"c08c08f0",
X"050883c0",
X"8c08e005",
X"0c83c08c",
X"08fc050c",
X"83c08c08",
X"f0050889",
X"278a3889",
X"0b83c08c",
X"08e0050c",
X"83c08c08",
X"e0050886",
X"0587fffc",
X"0683c08c",
X"08e0050c",
X"0283c08c",
X"08e00508",
X"310d853d",
X"705583c0",
X"8c08ec05",
X"085483c0",
X"8c08f005",
X"085383c0",
X"8c08f405",
X"085283c0",
X"8c08e405",
X"0c80d9f2",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"e4050883",
X"c08c08ec",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"802e8c38",
X"83c08c08",
X"f805080d",
X"89c83983",
X"c08c08f0",
X"0508802e",
X"89a63883",
X"c08c08ec",
X"05088105",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e0050884",
X"2ea93884",
X"0b83c08c",
X"08e00508",
X"2588c738",
X"83c08c08",
X"e0050885",
X"2e859b38",
X"83c08c08",
X"e00508a1",
X"2e87ad38",
X"88ac3980",
X"0b83c08c",
X"08ec0508",
X"85053383",
X"c08c08e0",
X"050c83c0",
X"8c08fc05",
X"0c83c08c",
X"08e00508",
X"832e0981",
X"06888338",
X"83c08c08",
X"e8050881",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"812687e6",
X"38810b83",
X"c08c08e0",
X"050880d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"fc050c83",
X"c08c08ec",
X"05088205",
X"3383c08c",
X"08e00508",
X"87053483",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c80",
X"0b83c08c",
X"08e00508",
X"8b053483",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"f4050c80",
X"0b83c08c",
X"08e00508",
X"8c053483",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c80",
X"0b83c08c",
X"08e00508",
X"8d053483",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"f4050c80",
X"0b83c08c",
X"08e00508",
X"8e052383",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c80",
X"0b83c08c",
X"08e00508",
X"8a053483",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"05709405",
X"08fcffff",
X"06719405",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"ec050886",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"83c08c08",
X"e0050883",
X"c08c08fc",
X"05082e09",
X"8106b638",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"83c08c08",
X"fc050883",
X"c08c08e0",
X"05088b05",
X"3483c08c",
X"08ec0508",
X"87053383",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08812e8f",
X"3883c08c",
X"08e00508",
X"822eb738",
X"848c3983",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"f4050c82",
X"0b83c08c",
X"08e00508",
X"8a053483",
X"d93983c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c83c0",
X"8c08fc05",
X"0883c08c",
X"08e00508",
X"8a053483",
X"a13983c0",
X"8c08fc05",
X"08802e83",
X"953883c0",
X"8c08ec05",
X"08830533",
X"830683c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"832e0981",
X"0682f338",
X"83c08c08",
X"ec050882",
X"05337098",
X"2b83c08c",
X"08e0050c",
X"83c08c08",
X"e4050c83",
X"c08c08e0",
X"05088025",
X"82cc3883",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"f4050c83",
X"c08c08ec",
X"05088605",
X"3383c08c",
X"08e00508",
X"80d60534",
X"83c08c08",
X"e0050884",
X"0583c08c",
X"08ec0508",
X"8205338f",
X"0683c08c",
X"08e4050c",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050883c0",
X"8c08e005",
X"083483c0",
X"8c08ec05",
X"08840533",
X"83c08c08",
X"e0050881",
X"0534800b",
X"83c08c08",
X"e0050882",
X"053483c0",
X"8c08e005",
X"0808ff83",
X"ff068280",
X"0783c08c",
X"08e00508",
X"0c83c08c",
X"08e80508",
X"81053381",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e0050883",
X"c08c08e8",
X"05088105",
X"34818339",
X"83c08c08",
X"fc050880",
X"2e80f738",
X"83c08c08",
X"ec050886",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"a22e0981",
X"0680d738",
X"83c08c08",
X"ec050888",
X"053383c0",
X"8c08ec05",
X"08870533",
X"71828029",
X"0583c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c5283",
X"c08c08e4",
X"050c83c0",
X"8c08f405",
X"0c83c08c",
X"08e40508",
X"83c08c08",
X"e0050888",
X"052383c0",
X"8c08ec05",
X"083383c0",
X"8c08f005",
X"08713170",
X"83ffff06",
X"83c08c08",
X"f0050c83",
X"c08c08e0",
X"050c83c0",
X"8c08ec05",
X"080583c0",
X"8c08ec05",
X"0cf6d039",
X"83c08c08",
X"f805080d",
X"83c08c08",
X"f0050883",
X"c08c08e0",
X"050c83c0",
X"8c08f805",
X"080d83c0",
X"8c08e005",
X"0883c080",
X"0c8d3d0d",
X"83c08c0c",
X"0483c08c",
X"080283c0",
X"8c0ce63d",
X"0d83c08c",
X"08880508",
X"02840583",
X"c08c08e8",
X"050c83c0",
X"8c08d405",
X"0c800b83",
X"cafc3483",
X"c08c08d4",
X"05089005",
X"83c08c08",
X"c0050c80",
X"0b83c08c",
X"08c00508",
X"34800b83",
X"c08c08c0",
X"05088105",
X"34800b83",
X"c08c08c4",
X"050c83c0",
X"8c08c405",
X"0880d829",
X"83c08c08",
X"c0050805",
X"83c08c08",
X"ffb4050c",
X"800b83c0",
X"8c08ffb4",
X"050880d8",
X"050c83c0",
X"8c08ffb4",
X"05088405",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"c4050883",
X"c08c08ff",
X"b4050834",
X"880b83c0",
X"8c08ffb4",
X"05088105",
X"34800b83",
X"c08c08ff",
X"b4050882",
X"053483c0",
X"8c08ffb4",
X"050808ff",
X"a1ff06a0",
X"800783c0",
X"8c08ffb4",
X"05080c83",
X"c08c08c4",
X"05088105",
X"7081ff06",
X"83c08c08",
X"c4050c83",
X"c08c08ff",
X"b4050c81",
X"0b83c08c",
X"08c40508",
X"27fedb38",
X"83c08c08",
X"ec057054",
X"83c08c08",
X"c8050c92",
X"5283c08c",
X"08d40508",
X"5180cd99",
X"3f83c080",
X"0881ff06",
X"7083c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"088dea38",
X"83c08c08",
X"f40551f1",
X"8c3f83c0",
X"800883ff",
X"ff0683c0",
X"8c08f605",
X"5283c08c",
X"08e4050c",
X"f0f33f83",
X"c0800883",
X"ffff0683",
X"c08c08fd",
X"053383c0",
X"8c08ffb8",
X"050883c0",
X"8c08c405",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"c4050883",
X"c08c08ff",
X"bc050827",
X"80fe3883",
X"c08c08c8",
X"05085483",
X"c08c08c4",
X"05085389",
X"5283c08c",
X"08d40508",
X"5180cc9e",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"80f23883",
X"c08c08ee",
X"0551eff1",
X"3f83c080",
X"0883ffff",
X"065383c0",
X"8c08c405",
X"085283c0",
X"8c08d405",
X"0851f0b3",
X"3f83c08c",
X"08c40508",
X"81057081",
X"ff0683c0",
X"8c08c405",
X"0c83c08c",
X"08ffb405",
X"0cfef139",
X"83c08c08",
X"c0050881",
X"053383c0",
X"8c08ffb4",
X"050c81db",
X"0b83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffb405",
X"08802e8b",
X"e0389439",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"ffbc050c",
X"8bcb3983",
X"c08c08f1",
X"05335283",
X"c08c08d4",
X"05085180",
X"cb9c3f80",
X"0b83c08c",
X"08c00508",
X"81053383",
X"c08c08ff",
X"b4050c83",
X"c08c08c4",
X"050c83c0",
X"8c08c405",
X"0883c08c",
X"08ffb405",
X"082789e6",
X"3883c08c",
X"08c40508",
X"80d82970",
X"83c08c08",
X"c0050805",
X"70880570",
X"83053383",
X"c08c08cc",
X"050c83c0",
X"8c08c805",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08d8050c",
X"83c08c08",
X"cc050887",
X"a63883c0",
X"8c08c805",
X"08220284",
X"05718605",
X"87fffc06",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"dc050c83",
X"c08c08ff",
X"b8050c02",
X"83c08c08",
X"ffb40508",
X"310d893d",
X"705983c0",
X"8c08ffb8",
X"05085883",
X"c08c08ff",
X"bc050887",
X"05335783",
X"c08c08ff",
X"b4050ca2",
X"5583c08c",
X"08cc0508",
X"54865381",
X"815283c0",
X"8c08d405",
X"0851be93",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"d0050c83",
X"c08c08d0",
X"050881c1",
X"3883c08c",
X"08ffbc05",
X"08960553",
X"83c08c08",
X"ffb80508",
X"5283c08c",
X"08ffb405",
X"0851a1c6",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb40508",
X"802e8185",
X"3883c08c",
X"08ffbc05",
X"08940583",
X"c08c08ff",
X"bc050896",
X"05337086",
X"2a83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08cc050c",
X"83c08c08",
X"ffb40508",
X"832e0981",
X"0680c638",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"c8050882",
X"053483ca",
X"e0337081",
X"0583c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb405",
X"0883cae0",
X"3483c08c",
X"08ffb805",
X"0883c08c",
X"08cc0508",
X"3483c08c",
X"08dc0508",
X"0d83c08c",
X"08d00508",
X"81ff0683",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b80508fb",
X"ff3883c0",
X"8c08d805",
X"0883c08c",
X"08c00508",
X"05880570",
X"82053351",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb40508",
X"832e0981",
X"0680e338",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb40508",
X"81057081",
X"ff065183",
X"c08c08ff",
X"b4050c81",
X"0b83c08c",
X"08ffb405",
X"0827dd38",
X"800b83c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb4",
X"05088105",
X"7081ff06",
X"5183c08c",
X"08ffb405",
X"0c970b83",
X"c08c08ff",
X"b4050827",
X"dd3883c0",
X"8c08e405",
X"0880f932",
X"70307080",
X"25515183",
X"c08c08ff",
X"b4050c83",
X"c08c08e0",
X"0508912e",
X"09810680",
X"f93883c0",
X"8c08ffb4",
X"0508802e",
X"80ec3883",
X"c08c08c4",
X"050880e2",
X"38850b83",
X"c08c08c0",
X"0508a605",
X"34a00b83",
X"c08c08c0",
X"0508a705",
X"34850b83",
X"c08c08c0",
X"0508a805",
X"3480c00b",
X"83c08c08",
X"c00508a9",
X"0534860b",
X"83c08c08",
X"c00508aa",
X"0534900b",
X"83c08c08",
X"c00508ab",
X"0534860b",
X"83c08c08",
X"c00508ac",
X"0534a00b",
X"83c08c08",
X"c00508ad",
X"053483c0",
X"8c08e405",
X"0889d832",
X"70307080",
X"25515183",
X"c08c08ff",
X"b4050c83",
X"c08c08e0",
X"050883ed",
X"ec2e0981",
X"0680f638",
X"817083c0",
X"8c08ffb4",
X"05080683",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b4050880",
X"2e80ce38",
X"83c08c08",
X"c4050880",
X"c438840b",
X"83c08c08",
X"c00508aa",
X"053480c0",
X"0b83c08c",
X"08c00508",
X"ab053484",
X"0b83c08c",
X"08c00508",
X"ac053490",
X"0b83c08c",
X"08c00508",
X"ad053483",
X"c08c08ff",
X"b8050883",
X"c08c08c0",
X"05088c05",
X"3483c08c",
X"08e40508",
X"80f93270",
X"30708025",
X"515183c0",
X"8c08ffb4",
X"050c83c0",
X"8c08e005",
X"08862e09",
X"810680c3",
X"38817083",
X"c08c08ff",
X"b4050806",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb40508",
X"802e9c38",
X"83c08c08",
X"c4050893",
X"3883c08c",
X"08ffb805",
X"0883c08c",
X"08c00508",
X"8d053483",
X"c08c08c4",
X"050880d8",
X"2983c08c",
X"08c00508",
X"05708405",
X"70830533",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"c8050c83",
X"c08c08ff",
X"bc050c80",
X"58805783",
X"c08c08ff",
X"b4050856",
X"80558054",
X"8a53a152",
X"83c08c08",
X"d4050851",
X"b78d3f83",
X"c0800881",
X"ff067030",
X"709f2a51",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"a02e8c38",
X"83c08c08",
X"ffb40508",
X"f6c23883",
X"c08c08ff",
X"bc05088b",
X"053383c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb4",
X"0508802e",
X"b33883c0",
X"8c08c805",
X"08830533",
X"83c08c08",
X"ffb4050c",
X"80588057",
X"83c08c08",
X"ffb40508",
X"56805580",
X"548b53a1",
X"5283c08c",
X"08d40508",
X"51b6883f",
X"83c08c08",
X"c4050881",
X"057081ff",
X"0683c08c",
X"08c00508",
X"81053352",
X"83c08c08",
X"c4050c83",
X"c08c08ff",
X"b4050cf6",
X"8939800b",
X"83c08c08",
X"c4050c83",
X"c08c08c4",
X"050880d8",
X"2983c08c",
X"08d40508",
X"05709a05",
X"3383c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb405",
X"08822e09",
X"8106a938",
X"83cafc56",
X"81558054",
X"83c08c08",
X"ffb40508",
X"5383c08c",
X"08ffb805",
X"08970533",
X"5283c08c",
X"08d40508",
X"51e48a3f",
X"83c08c08",
X"c4050881",
X"057081ff",
X"0683c08c",
X"08c4050c",
X"83c08c08",
X"ffb4050c",
X"810b83c0",
X"8c08c405",
X"0827fefb",
X"38810b83",
X"c08c08c0",
X"05083480",
X"0b83c08c",
X"08ffbc05",
X"0c83c08c",
X"08e80508",
X"0d83c08c",
X"08ffbc05",
X"0883c080",
X"0c9c3d0d",
X"83c08c0c",
X"04f53d0d",
X"901e5780",
X"0b811833",
X"54597873",
X"27819d38",
X"7880d829",
X"178a1133",
X"54547283",
X"2e098106",
X"80f83894",
X"14335ba9",
X"8c3f83c0",
X"80085a80",
X"567581c4",
X"291a8711",
X"33545472",
X"802e80c0",
X"38730881",
X"d7e42e09",
X"8106b538",
X"80745955",
X"7480d829",
X"189a1133",
X"54547283",
X"2e098106",
X"9238a414",
X"70335454",
X"7a732787",
X"38ff1353",
X"72743481",
X"157081ff",
X"06565381",
X"7527d138",
X"81167081",
X"ff065753",
X"8f7627ff",
X"a43883ca",
X"e033ff05",
X"537283ca",
X"e0348119",
X"7081ff06",
X"8119335e",
X"5a537b79",
X"26fee538",
X"800b83c0",
X"800c8d3d",
X"0d0483c0",
X"8c080283",
X"c08c0ce6",
X"3d0d83c0",
X"8c088805",
X"08028405",
X"71900570",
X"337083c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08c805",
X"0c83c08c",
X"08dc050c",
X"83c08c08",
X"e0050c83",
X"c08c08ff",
X"a4050880",
X"2e94b538",
X"800b83c0",
X"8c08c805",
X"08810533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"d4050c83",
X"c08c08d4",
X"050883c0",
X"8c08ffa4",
X"05082593",
X"fd3883c0",
X"8c08d405",
X"0880d829",
X"83c08c08",
X"c8050805",
X"84057086",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"938938a6",
X"b23f83c0",
X"8c08ffb8",
X"050880d4",
X"050883c0",
X"80082692",
X"f2380283",
X"c08c08ff",
X"b8050881",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08d805",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08fc0523",
X"83c08c08",
X"ffa40508",
X"860583fc",
X"0683c08c",
X"08ffa405",
X"0c0283c0",
X"8c08ffa4",
X"0508310d",
X"853d7055",
X"83c08c08",
X"fc055483",
X"c08c08ff",
X"b8050853",
X"83c08c08",
X"e0050852",
X"83c08c08",
X"c0050cae",
X"8a3f83c0",
X"800881ff",
X"0683c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"0891bb38",
X"83c08c08",
X"ffb80508",
X"87053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e80d538",
X"83c08c08",
X"ffb80508",
X"86053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050882",
X"2e098106",
X"b33883c0",
X"8c08fc05",
X"2283c08c",
X"08ffa405",
X"0c870b83",
X"c08c08ff",
X"a4050827",
X"973883c0",
X"8c08c005",
X"08820552",
X"83c08c08",
X"c0050833",
X"51dba63f",
X"83c08c08",
X"ffb80508",
X"86053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050883",
X"2e098106",
X"90a43883",
X"c08c08ff",
X"b8050892",
X"05708205",
X"3383c08c",
X"08fc0522",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"c4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"a8050826",
X"8fe43880",
X"0b83c08c",
X"08e4050c",
X"800b83c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffb0",
X"05081083",
X"c08c0805",
X"f80583c0",
X"8c08ffb0",
X"05088429",
X"83c08c08",
X"ffb00508",
X"100583c0",
X"8c08c405",
X"08057084",
X"05703383",
X"c08c08c0",
X"05080570",
X"3383c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffb405",
X"0883c08c",
X"08ffbc05",
X"082383c0",
X"8c08ffa8",
X"05088105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08902e09",
X"8106be38",
X"83c08c08",
X"ffa80508",
X"3383c08c",
X"08c00508",
X"05810570",
X"33708280",
X"2983c08c",
X"08ffb405",
X"08055151",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffbc0508",
X"2383c08c",
X"08ffac05",
X"08860522",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa80508",
X"a23883c0",
X"8c08ffac",
X"05088805",
X"2283c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"0881ff2e",
X"80e53883",
X"c08c08ff",
X"bc050822",
X"7083c08c",
X"08ffa805",
X"08317082",
X"80297131",
X"83c08c08",
X"ffac0508",
X"88052270",
X"83c08c08",
X"ffa80508",
X"31707335",
X"5383c08c",
X"08ffa805",
X"0c83c08c",
X"08ffac05",
X"0c5183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffbc",
X"05082383",
X"c08c08ff",
X"b0050881",
X"057081ff",
X"0683c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa405",
X"0c810b83",
X"c08c08ff",
X"b0050827",
X"fce03883",
X"c08c08f8",
X"052283c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508bf26",
X"913883c0",
X"8c08e405",
X"08820783",
X"c08c08e4",
X"050c81c0",
X"0b83c08c",
X"08ffa405",
X"08279138",
X"83c08c08",
X"e4050881",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"fa052283",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a40508bf",
X"26913883",
X"c08c08e4",
X"05088807",
X"83c08c08",
X"e4050c81",
X"c00b83c0",
X"8c08ffa4",
X"05082791",
X"3883c08c",
X"08e40508",
X"840783c0",
X"8c08e405",
X"0c800b83",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"b0050810",
X"83c08c08",
X"c4050805",
X"70900570",
X"3383c08c",
X"08c00508",
X"05703372",
X"81053370",
X"72065153",
X"5183c08c",
X"08ffa805",
X"0c5183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"9b38900b",
X"83c08c08",
X"ffb00508",
X"2b83c08c",
X"08e40508",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"ffb00508",
X"81057081",
X"ff0683c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa4",
X"050c970b",
X"83c08c08",
X"ffb00508",
X"27fef438",
X"83c08c08",
X"ffb80508",
X"90053383",
X"c08c08e4",
X"050883c0",
X"8c08ffb4",
X"050c83c0",
X"8c08c405",
X"0c83c08c",
X"08ffb405",
X"0883c08c",
X"08ffb805",
X"088c0508",
X"2e83ff38",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffb80508",
X"8c050c83",
X"c08c08ff",
X"b8050889",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"83b93883",
X"c08c08e4",
X"0583c08c",
X"08ffb405",
X"088f0683",
X"c08c08e4",
X"050c83c0",
X"8c08cc05",
X"0c800b83",
X"c08c08f0",
X"050c800b",
X"83c08c08",
X"f4052380",
X"0b81d9e0",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffbc05",
X"082e82d3",
X"3883c08c",
X"08f00581",
X"d9e00b83",
X"c08c08ff",
X"ac050c83",
X"c08c08d0",
X"050c83c0",
X"8c08ffac",
X"05083383",
X"c08c08ff",
X"ac050881",
X"05338172",
X"2b81722b",
X"077083c0",
X"8c08ffb4",
X"05080652",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffa80508",
X"2e098106",
X"81be3883",
X"c08c08ff",
X"bc050885",
X"2680f638",
X"83c08c08",
X"ffac0508",
X"82053370",
X"81ff0683",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a4050880",
X"2e80ca38",
X"83c08c08",
X"ffbc0508",
X"83c08c08",
X"ffbc0508",
X"81057081",
X"ff0683c0",
X"8c08d005",
X"08730553",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb00508",
X"83c08c08",
X"ffa40508",
X"3483c08c",
X"08ffac05",
X"08830533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9d38",
X"810b83c0",
X"8c08ffa4",
X"05082b83",
X"c08c08cc",
X"05080807",
X"83c08c08",
X"cc05080c",
X"83c08c08",
X"ffac0508",
X"84057033",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa40508",
X"fdc83883",
X"c08c08f0",
X"05528051",
X"d0c33f83",
X"c08c08e4",
X"05085283",
X"c08c08c4",
X"050851d1",
X"fe3f83c0",
X"8c08fb05",
X"33708180",
X"0a29810a",
X"0570982c",
X"5583c08c",
X"08ffa405",
X"0c83c08c",
X"08f90533",
X"7081800a",
X"29810a05",
X"70982c55",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"c4050853",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa8050c",
X"d1d43f83",
X"c08c08ff",
X"b8050888",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"84e03883",
X"c08c08ff",
X"b8050890",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"05088126",
X"84c03880",
X"7081da94",
X"0b81da94",
X"0b810533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffb40508",
X"2e81ae38",
X"83c08c08",
X"ffac0508",
X"842983c0",
X"8c08ffa8",
X"05080570",
X"3383c08c",
X"08c00508",
X"05703372",
X"81053370",
X"72065153",
X"5183c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802eaa",
X"38810b83",
X"c08c08ff",
X"ac05082b",
X"83c08c08",
X"ffb40508",
X"077083ff",
X"ff0683c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffac",
X"05088105",
X"7081ff06",
X"81da9471",
X"84297105",
X"70810533",
X"515383c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508fed4",
X"3883c08c",
X"08ffb805",
X"088a0522",
X"83c08c08",
X"c0050c83",
X"c08c08ff",
X"b4050883",
X"c08c08c0",
X"05082e82",
X"ad38800b",
X"83c08c08",
X"e8050c80",
X"0b83c08c",
X"08ec0523",
X"807083c0",
X"8c08e805",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffb0050c",
X"81af3983",
X"c08c08ff",
X"b4050883",
X"c08c08ff",
X"ac05082c",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e80e7",
X"3883c08c",
X"08ffb005",
X"0883c08c",
X"08ffb005",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"bc050873",
X"0583c08c",
X"08ffb805",
X"08900533",
X"83c08c08",
X"ffac0508",
X"84290553",
X"5383c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa805",
X"0881da96",
X"053383c0",
X"8c08ffa4",
X"05083483",
X"c08c08ff",
X"ac050881",
X"057081ff",
X"0683c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa405",
X"0c8f0b83",
X"c08c08ff",
X"ac050827",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb00508",
X"85268c38",
X"83c08c08",
X"ffa40508",
X"fea93883",
X"c08c08e8",
X"05528051",
X"caf33f83",
X"c08c08ff",
X"b4050883",
X"c08c08ff",
X"b805088a",
X"052383c0",
X"8c08ffb8",
X"050880d2",
X"053383c0",
X"8c08ffb8",
X"050880d4",
X"05080583",
X"c08c08ff",
X"b8050880",
X"d4050c83",
X"c08c08d8",
X"05080d83",
X"c08c08d4",
X"05088180",
X"0a298180",
X"0a057098",
X"2c83c08c",
X"08c80508",
X"81053383",
X"c08c08ff",
X"a8050c51",
X"83c08c08",
X"d4050c83",
X"c08c08ff",
X"a8050883",
X"c08c08d4",
X"050824ec",
X"8538800b",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"dc05080d",
X"83c08c08",
X"ffa80508",
X"83c0800c",
X"9c3d0d83",
X"c08c0c04",
X"f33d0d02",
X"bf053302",
X"840580c3",
X"053383ca",
X"fc335a5b",
X"5979802e",
X"8d387878",
X"06577680",
X"2e8e3881",
X"89397878",
X"06577680",
X"2e80ff38",
X"83cafc33",
X"707a0758",
X"58798838",
X"78097079",
X"06515776",
X"83cafc34",
X"92973f83",
X"c080085e",
X"805c8f5d",
X"7d1c8711",
X"33585876",
X"802e80c1",
X"38770881",
X"d7e42e09",
X"8106b638",
X"805b815a",
X"7d1c701c",
X"9a113359",
X"59597682",
X"2e098106",
X"943883ca",
X"fc568155",
X"80547653",
X"97183352",
X"7851cbc5",
X"3fff1a80",
X"d81c5c5a",
X"798025d0",
X"38ff1d81",
X"c41d5d5d",
X"7c8025ff",
X"a7388f3d",
X"0d04e93d",
X"0d696c02",
X"880580ea",
X"05225c5a",
X"5b807071",
X"415e58ff",
X"78797a7b",
X"7c7d464c",
X"4a45405d",
X"4362993d",
X"34620284",
X"0580dd05",
X"34777922",
X"80ffff06",
X"54457279",
X"2379782e",
X"8887387a",
X"7081055c",
X"3370842a",
X"718c0670",
X"822a5a56",
X"568306ff",
X"1b7083ff",
X"ff065c54",
X"56805475",
X"742e9138",
X"7a708105",
X"5c33ff1b",
X"7083ffff",
X"065c5454",
X"8176279b",
X"387381ff",
X"067b7081",
X"055d3355",
X"74828029",
X"05ff1b70",
X"83ffff06",
X"5c545482",
X"7627aa38",
X"7383ffff",
X"067b7081",
X"055d3370",
X"902b7207",
X"7d708105",
X"5f337098",
X"2b7207fe",
X"1f7083ff",
X"ff064052",
X"52525254",
X"547e802e",
X"80c43876",
X"86f73874",
X"8a2e0981",
X"06943881",
X"1f7081ff",
X"06811e70",
X"81ff065f",
X"52405386",
X"dc39748c",
X"2e098106",
X"86d338ff",
X"1f7081ff",
X"06ff1e70",
X"81ff065f",
X"5240537b",
X"632586bd",
X"38ff4386",
X"b8397681",
X"2e83bb38",
X"76812489",
X"3876802e",
X"8d3886a5",
X"3976822e",
X"84a63886",
X"9c39f815",
X"53728426",
X"84953872",
X"842981da",
X"d4055372",
X"08046480",
X"2e80cd38",
X"78228380",
X"80065372",
X"8380802e",
X"098106bc",
X"38805675",
X"6427a438",
X"751e7083",
X"ffff0677",
X"101b9011",
X"72832a58",
X"51575153",
X"73753472",
X"87068171",
X"2b515372",
X"81163481",
X"167081ff",
X"06575397",
X"7627cc38",
X"7f840740",
X"800b993d",
X"43566116",
X"70337098",
X"2b70982c",
X"51515153",
X"80732480",
X"fb386073",
X"291e7083",
X"ffff067a",
X"22838080",
X"06525853",
X"72838080",
X"2e098106",
X"80de3860",
X"88327030",
X"70720780",
X"25639032",
X"70307072",
X"07802573",
X"07535458",
X"51555373",
X"802ebd38",
X"76870653",
X"72b63875",
X"84297610",
X"05791184",
X"1179832a",
X"57575153",
X"73753460",
X"81163465",
X"86142366",
X"88142375",
X"87387f81",
X"07408d39",
X"75812e09",
X"81068538",
X"7f820740",
X"81167081",
X"ff065753",
X"817627fe",
X"e5386361",
X"291e7083",
X"ffff065f",
X"53807046",
X"42ff0284",
X"0580dd05",
X"34ff0b99",
X"3d3483f5",
X"39811c70",
X"81ff065d",
X"53804273",
X"812e0981",
X"068e3877",
X"81800a29",
X"81800a05",
X"5880d339",
X"73802e89",
X"3873822e",
X"0981068d",
X"387c8180",
X"0a298180",
X"0a055da4",
X"39815f83",
X"b839ff1c",
X"7081ff06",
X"5d537b63",
X"258338ff",
X"437c802e",
X"92387c81",
X"800a2981",
X"ff0a055d",
X"7c982c5d",
X"83933977",
X"802e9238",
X"7781800a",
X"2981ff0a",
X"05587798",
X"2c5882fd",
X"39775383",
X"9e397489",
X"2680f438",
X"74842981",
X"dae80553",
X"72080473",
X"872e82e1",
X"3873852e",
X"82db3873",
X"882e82d5",
X"38738c2e",
X"82cf3873",
X"892e0981",
X"06863881",
X"4582c239",
X"73812e09",
X"810682b9",
X"38628025",
X"82b3387b",
X"982b7098",
X"2c514382",
X"a8397383",
X"ffff0646",
X"829f3973",
X"83ffff06",
X"47829639",
X"7381ff06",
X"41828e39",
X"73811a34",
X"82873973",
X"81ff0644",
X"81ff397e",
X"5382a039",
X"74812e81",
X"e3387481",
X"24893874",
X"802e8d38",
X"81e73974",
X"822e81d8",
X"3881de39",
X"74567b83",
X"38815674",
X"5373862e",
X"09810697",
X"38758106",
X"5372802e",
X"8e387822",
X"82ffff06",
X"fe808007",
X"53b6397b",
X"83388153",
X"73822e09",
X"81069738",
X"72810653",
X"72802e8e",
X"38782281",
X"ffff0681",
X"80800753",
X"93397b96",
X"38fc1453",
X"7281268e",
X"387822ff",
X"80800753",
X"72792380",
X"e5398055",
X"73812e09",
X"81068338",
X"73557753",
X"77802e89",
X"38748106",
X"537280ca",
X"3872d015",
X"54557281",
X"26833881",
X"5577802e",
X"b9387481",
X"06537280",
X"2eb03878",
X"22838080",
X"06537283",
X"80802e09",
X"81069f38",
X"73b02e09",
X"81068738",
X"61993d34",
X"913973b1",
X"2e098106",
X"89386102",
X"840580dd",
X"05346181",
X"05538c39",
X"61743181",
X"05538439",
X"61145372",
X"83ffff06",
X"4279f7fb",
X"387d832a",
X"5372821a",
X"34782283",
X"80800653",
X"72838080",
X"2e098106",
X"88388153",
X"7f872e83",
X"38805372",
X"83c0800c",
X"993d0d04",
X"fd3d0d75",
X"83113382",
X"12337198",
X"2b71902b",
X"07811433",
X"70882b72",
X"07753371",
X"0783c080",
X"0c525354",
X"56545285",
X"3d0d04f6",
X"3d0d02b7",
X"05330284",
X"05bb0533",
X"028805bf",
X"05335b5b",
X"5b805880",
X"5778882b",
X"7a075680",
X"557a5481",
X"53a3527c",
X"5192cc3f",
X"83c08008",
X"81ff0683",
X"c0800c8c",
X"3d0d04f6",
X"3d0d02b7",
X"05330284",
X"05bb0533",
X"028805bf",
X"05335b5b",
X"5b805880",
X"5778882b",
X"7a075680",
X"557a5483",
X"53a3527c",
X"5192903f",
X"83c08008",
X"81ff0683",
X"c0800c8c",
X"3d0d04f7",
X"3d0d02b3",
X"05330284",
X"05b60522",
X"605a5856",
X"80558054",
X"805381a3",
X"527b5191",
X"e23f83c0",
X"800881ff",
X"0683c080",
X"0c8b3d0d",
X"04ee3d0d",
X"6490115c",
X"5c807b34",
X"800b841c",
X"0c800b88",
X"1c34810b",
X"891c3488",
X"0b8a1c34",
X"800b8b1c",
X"34881b08",
X"c1068107",
X"881c0c8f",
X"3d70545d",
X"88527b51",
X"9beb3f83",
X"c0800881",
X"ff06705b",
X"597881a9",
X"38903d33",
X"5e81db5a",
X"7d892e09",
X"81068199",
X"387c5392",
X"527b519b",
X"c43f83c0",
X"800881ff",
X"06705b59",
X"78818238",
X"7c588857",
X"7856a955",
X"78548653",
X"81a0527b",
X"5190d03f",
X"83c08008",
X"81ff0670",
X"5b597880",
X"e03802ba",
X"05337b34",
X"7c547853",
X"7d527b51",
X"9bac3f83",
X"c0800881",
X"ff06705b",
X"597880c1",
X"3802bd05",
X"33527b51",
X"9bc43f83",
X"c0800881",
X"ff06705b",
X"5978aa38",
X"817b335a",
X"5a797926",
X"99388054",
X"79538852",
X"7b51fdbb",
X"3f811a70",
X"81ff067c",
X"33525b59",
X"e439810b",
X"881c3480",
X"5a7983c0",
X"800c943d",
X"0d04800b",
X"83c0800c",
X"04f93d0d",
X"79028405",
X"ab05338e",
X"3d705458",
X"5858ffbe",
X"b03f8a3d",
X"8a0551ff",
X"bea73f75",
X"51fc8d3f",
X"83c08008",
X"8486812e",
X"be3883c0",
X"80088486",
X"81269938",
X"83c08008",
X"8482802e",
X"80e63883",
X"c0800884",
X"82812e9f",
X"3881b439",
X"83c08008",
X"80c08283",
X"2e80f438",
X"83c08008",
X"80c08683",
X"2e80e838",
X"81993983",
X"c09c3355",
X"80567476",
X"2e098106",
X"818b3874",
X"54765391",
X"527751fb",
X"d63f7454",
X"76539052",
X"7751fbcb",
X"3f745476",
X"53845277",
X"51fbfc3f",
X"810b83c0",
X"9c3481b1",
X"5680de39",
X"80547653",
X"91527751",
X"fba93f80",
X"54765390",
X"527751fb",
X"9e3f800b",
X"83c09c34",
X"76528718",
X"33519796",
X"3fb53980",
X"54765394",
X"527751fb",
X"823f8054",
X"76539052",
X"7751faf7",
X"3f7551ff",
X"bcdb3f83",
X"c0800889",
X"2a810653",
X"76528718",
X"335190cd",
X"3f800b83",
X"c09c3480",
X"567583c0",
X"800c893d",
X"0d04f23d",
X"0d609011",
X"5a58800b",
X"881a3371",
X"59565674",
X"762e82a5",
X"3882ac3f",
X"84190883",
X"c0800826",
X"82953878",
X"335a810b",
X"8e3d2390",
X"3df81155",
X"f4055399",
X"18527751",
X"8ae53f83",
X"c0800881",
X"ff067057",
X"5574772e",
X"09810681",
X"d9388639",
X"745681d2",
X"39815682",
X"578e3d33",
X"77065574",
X"802ebb38",
X"800b8d3d",
X"34903df0",
X"05548453",
X"75527751",
X"facd3f83",
X"c0800881",
X"ff065574",
X"9d387b53",
X"75527751",
X"fce73f83",
X"c0800881",
X"ff065574",
X"81b12e81",
X"8b3874ff",
X"b3387610",
X"81fc0681",
X"177081ff",
X"06585657",
X"877627ff",
X"a8388156",
X"757a2680",
X"eb38800b",
X"8d3d348c",
X"3d705557",
X"84537552",
X"7751f9f7",
X"3f83c080",
X"0881ff06",
X"557480c1",
X"387651ff",
X"bad73f83",
X"c0800882",
X"87065574",
X"82812e09",
X"8106aa38",
X"02ae0533",
X"81075574",
X"028405ae",
X"05347b53",
X"75527751",
X"fbeb3f83",
X"c0800881",
X"ff065574",
X"81b12e90",
X"3874feb8",
X"38811670",
X"81ff0657",
X"55ff9139",
X"80567581",
X"ff065697",
X"3f83c080",
X"088fd005",
X"841a0c75",
X"577683c0",
X"800c903d",
X"0d040490",
X"80a00883",
X"c0800c04",
X"ff3d0d73",
X"87e82951",
X"ff8fa83f",
X"833d0d04",
X"0483cb80",
X"0b83c080",
X"0c04fd3d",
X"0d757754",
X"54800b83",
X"cae03472",
X"8a389090",
X"800b8415",
X"0c903972",
X"812e0981",
X"06883890",
X"98800b84",
X"150c8414",
X"0883caf8",
X"0c800b88",
X"150c800b",
X"8c150c83",
X"caf80853",
X"820b8780",
X"14348151",
X"ff9e3f83",
X"caf80853",
X"800b8814",
X"3483caf8",
X"0853810b",
X"87801434",
X"83caf808",
X"53800b8c",
X"143483ca",
X"f8085380",
X"0ba41434",
X"91743480",
X"0b83c0a0",
X"34800b83",
X"c0a43480",
X"0b83c0a8",
X"34805473",
X"81c42983",
X"cb840553",
X"800b8314",
X"34811470",
X"81ff0655",
X"538f7427",
X"e638853d",
X"0d04fe3d",
X"0d747682",
X"113370bf",
X"0681712b",
X"ff055651",
X"51525390",
X"71278338",
X"ff527651",
X"71712383",
X"caf80851",
X"87133390",
X"1234800b",
X"83c0a434",
X"800b83c0",
X"a8348813",
X"338a1433",
X"52527180",
X"2eaa3870",
X"81ff0651",
X"84527083",
X"38705271",
X"83c0a434",
X"8a133370",
X"30708025",
X"842b7088",
X"07515152",
X"537083c0",
X"a8349039",
X"7081ff06",
X"51708338",
X"98527183",
X"c0a83480",
X"0b83c080",
X"0c843d0d",
X"04f13d0d",
X"61656802",
X"8c0580cb",
X"05330290",
X"0580ce05",
X"22029405",
X"80d60522",
X"4240415a",
X"4040fd8b",
X"3f83c080",
X"08a78805",
X"5b807071",
X"5b5b5283",
X"943983ca",
X"f808517d",
X"94123483",
X"c0a43381",
X"07558070",
X"54567f86",
X"2680ea38",
X"7f842981",
X"db9c0583",
X"caf80853",
X"51700804",
X"800b8413",
X"34a13977",
X"33703070",
X"80258371",
X"31515152",
X"53708413",
X"348d3981",
X"0b841334",
X"b839830b",
X"84133481",
X"705456ad",
X"39810b84",
X"1334a239",
X"77337030",
X"70802583",
X"71315151",
X"52537084",
X"13348078",
X"33525270",
X"83388152",
X"71783481",
X"53748807",
X"5583c0a8",
X"3383caf8",
X"08525781",
X"0b81d012",
X"3483caf8",
X"0851810b",
X"81901234",
X"7e802eae",
X"3872802e",
X"a9387eff",
X"1e525470",
X"83ffff06",
X"537283ff",
X"ff2e9738",
X"73708105",
X"553383ca",
X"f8085351",
X"7081c013",
X"34ff1351",
X"de3983ca",
X"f808a811",
X"33535176",
X"88123483",
X"caf80851",
X"74713481",
X"ff529139",
X"83caf808",
X"a0113370",
X"81065152",
X"53708f38",
X"fafd3f7a",
X"83c08008",
X"26e63881",
X"8839810b",
X"a0143483",
X"caf808a8",
X"113380ff",
X"06707807",
X"52535170",
X"802e80ed",
X"3871862a",
X"70810651",
X"5170802e",
X"91388078",
X"33525370",
X"83388153",
X"72783480",
X"e0397184",
X"2a708106",
X"51517080",
X"2e9b3881",
X"197083ff",
X"ff067d30",
X"709f2a51",
X"525a5178",
X"7c2e0981",
X"06af38a4",
X"3971832a",
X"70810651",
X"5170802e",
X"9338811a",
X"7081ff06",
X"5b517983",
X"2e098106",
X"90388a39",
X"71a30651",
X"70802e85",
X"38715192",
X"39f9e43f",
X"7a83c080",
X"0826fce2",
X"387181bf",
X"06517083",
X"c0800c91",
X"3d0d04f6",
X"3d0d02b3",
X"05330284",
X"05b70533",
X"028805ba",
X"05225959",
X"59800b8c",
X"3d348c3d",
X"fc055680",
X"55805476",
X"53775278",
X"51fbf23f",
X"83c08008",
X"81ff0683",
X"c0800c8c",
X"3d0d04f3",
X"3d0d7f62",
X"64028c05",
X"80c20522",
X"72228115",
X"33425f41",
X"5e595980",
X"78237d53",
X"78335281",
X"51ffa03f",
X"83c08008",
X"81ff0656",
X"75802e86",
X"38755481",
X"ad3983ca",
X"f808a811",
X"33821b33",
X"70862a70",
X"81067398",
X"2b535157",
X"5c565779",
X"80258338",
X"81567376",
X"2e873881",
X"f0548182",
X"39818c17",
X"337081ff",
X"0679227d",
X"7131902b",
X"70902c70",
X"09709f2c",
X"72067052",
X"52535153",
X"57575475",
X"74248338",
X"75557484",
X"808029fc",
X"80800570",
X"902c5155",
X"74ff2e94",
X"3883caf8",
X"08818011",
X"33515473",
X"7c708105",
X"5e34db39",
X"77227605",
X"54737823",
X"7909709f",
X"2a708106",
X"821c3381",
X"bf067186",
X"2b075151",
X"51547382",
X"1a347c76",
X"268a3877",
X"22547a74",
X"26febb38",
X"80547383",
X"c0800c8f",
X"3d0d04f9",
X"3d0d7a57",
X"800b893d",
X"23893dfc",
X"05537652",
X"7951f8da",
X"3f83c080",
X"0881ff06",
X"70575574",
X"96387c54",
X"7b53883d",
X"22527651",
X"fde53f83",
X"c0800881",
X"ff065675",
X"83c0800c",
X"893d0d04",
X"f03d0d62",
X"66028805",
X"80ce0522",
X"415d5e80",
X"02840580",
X"d205227f",
X"810533ff",
X"115a5d5a",
X"5d81da58",
X"76bf2680",
X"e9387880",
X"2e80e138",
X"7a58787b",
X"27833878",
X"58821e33",
X"70872a58",
X"5a76923d",
X"34923dfc",
X"05567755",
X"7b547e53",
X"7d335282",
X"51f8de3f",
X"83c08008",
X"81ff065d",
X"800b923d",
X"33585a76",
X"802e8338",
X"815a821e",
X"3380ff06",
X"7a872b07",
X"5776821f",
X"347c9138",
X"78783170",
X"83ffff06",
X"791e5e5a",
X"57ff9b39",
X"7c587783",
X"c0800c92",
X"3d0d04f8",
X"3d0d7b02",
X"8405b205",
X"22585880",
X"0b8a3d23",
X"8a3dfc05",
X"5377527a",
X"51f6f73f",
X"83c08008",
X"81ff0670",
X"57557496",
X"387d5476",
X"53893d22",
X"527751fe",
X"af3f83c0",
X"800881ff",
X"06567583",
X"c0800c8a",
X"3d0d04ec",
X"3d0d666e",
X"02880580",
X"df053302",
X"8c0580e3",
X"05330290",
X"0580e705",
X"33029405",
X"80eb0533",
X"02980580",
X"ee052241",
X"43415f5c",
X"40570280",
X"f2052296",
X"3d23963d",
X"f0055384",
X"17705377",
X"5259f686",
X"3f83c080",
X"0881ff06",
X"587781e5",
X"38777a81",
X"80065840",
X"80772583",
X"38814079",
X"943d347b",
X"02840580",
X"c905347c",
X"02840580",
X"ca05347d",
X"02840580",
X"cb05347a",
X"953d347a",
X"882a5776",
X"02840580",
X"cd053495",
X"3d225776",
X"02840580",
X"ce053476",
X"882a5776",
X"02840580",
X"cf053477",
X"923d3496",
X"3dec1157",
X"578855f4",
X"1754923d",
X"22537752",
X"7751f695",
X"3f83c080",
X"0881ff06",
X"587780ed",
X"387e802e",
X"80cb3892",
X"3d227908",
X"58587f80",
X"2e9c3876",
X"81808007",
X"790c7e54",
X"963dfc05",
X"537783ff",
X"ff065278",
X"51f9fc3f",
X"99397682",
X"80800779",
X"0c7e5495",
X"3d225377",
X"83ffff06",
X"527851fc",
X"8f3f83c0",
X"800881ff",
X"0658779d",
X"38923d22",
X"5380527f",
X"30708025",
X"84713153",
X"5157f987",
X"3f83c080",
X"0881ff06",
X"587783c0",
X"800c963d",
X"0d04f63d",
X"0d7c0284",
X"05b70533",
X"5b5b8058",
X"80578056",
X"80557954",
X"85538052",
X"7a51fda3",
X"3f83c080",
X"0881ff06",
X"59788538",
X"79871c34",
X"7883c080",
X"0c8c3d0d",
X"04f93d0d",
X"02a70533",
X"028405ab",
X"05330288",
X"05af0533",
X"58595780",
X"0b83cb87",
X"33545472",
X"742e9f38",
X"81147081",
X"ff065553",
X"738f2681",
X"b6387381",
X"c42983cb",
X"84058311",
X"33515372",
X"e3387381",
X"c42983cb",
X"80055580",
X"0b871634",
X"76881634",
X"758a1634",
X"77891634",
X"80750c83",
X"caf8088c",
X"160c800b",
X"84163488",
X"0b851634",
X"800b8616",
X"34841508",
X"ffa1ff06",
X"a0800784",
X"160c8114",
X"7081ff06",
X"53537451",
X"febc3f83",
X"c0800881",
X"ff067055",
X"537280cd",
X"388a3973",
X"08750c72",
X"5480c239",
X"7281e1fc",
X"555681e1",
X"fc08802e",
X"b2387584",
X"29147008",
X"76537008",
X"51545472",
X"2d83c080",
X"0881ff06",
X"5372802e",
X"ce388116",
X"7081ff06",
X"81e1fc71",
X"84291153",
X"56575372",
X"08d03880",
X"547383c0",
X"800c893d",
X"0d04f93d",
X"0d795780",
X"0b841808",
X"83caf80c",
X"58f0883f",
X"88170883",
X"c0800827",
X"83ed38ef",
X"fa3f83c0",
X"80088105",
X"88180c83",
X"caf808b8",
X"11337081",
X"ff065151",
X"5473812e",
X"a4387381",
X"24883873",
X"782e8a38",
X"b8397382",
X"2e9538b1",
X"39763381",
X"f0065473",
X"902ea638",
X"917734a1",
X"39735876",
X"3381f006",
X"5473902e",
X"09810691",
X"38efa83f",
X"83c08008",
X"81c8058c",
X"180ca077",
X"34805675",
X"81c42983",
X"cb871133",
X"55557380",
X"2eaa3883",
X"cb801570",
X"08565474",
X"802e9d38",
X"88150880",
X"2e96388c",
X"140883ca",
X"f8082e09",
X"81068938",
X"73518815",
X"0854732d",
X"81167081",
X"ff065754",
X"8f7627ff",
X"ba387633",
X"5473b02e",
X"81993873",
X"b0248f38",
X"73912eab",
X"3873a02e",
X"80f53882",
X"a6397380",
X"d02e81e4",
X"387380d0",
X"248b3873",
X"80c02e81",
X"9938828f",
X"39738180",
X"2e81fb38",
X"82853980",
X"567581c4",
X"2983cb84",
X"11831133",
X"56595573",
X"802ea838",
X"83cb8015",
X"70085654",
X"74802e9b",
X"388c1408",
X"83caf808",
X"2e098106",
X"8e387351",
X"84150854",
X"732d800b",
X"83193481",
X"167081ff",
X"0657548f",
X"7627ffb9",
X"38927734",
X"81b539ed",
X"c23f8c17",
X"0883c080",
X"082781a7",
X"38b07734",
X"81a13983",
X"caf80854",
X"800b8c15",
X"3483caf8",
X"0854840b",
X"88153480",
X"c07734ed",
X"963f83c0",
X"8008b205",
X"8c180c80",
X"fa39ed87",
X"3f8c1708",
X"83c08008",
X"2780ec38",
X"83caf808",
X"54810b8c",
X"153483ca",
X"f8085480",
X"0b881534",
X"83caf808",
X"54880ba0",
X"1534ecdb",
X"3f83c080",
X"0894058c",
X"180c80d0",
X"7734bc39",
X"83caf808",
X"a0113370",
X"832a7081",
X"06515155",
X"5573802e",
X"a638880b",
X"a01634ec",
X"ae3f8c17",
X"0883c080",
X"08279438",
X"ff807734",
X"8e397753",
X"80528051",
X"fa8b3fff",
X"90773483",
X"caf808a0",
X"11337083",
X"2a708106",
X"51515555",
X"73802e86",
X"38880ba0",
X"1634893d",
X"0d04f63d",
X"0d02b305",
X"33028405",
X"b705335b",
X"5b800b83",
X"cb847084",
X"1272745d",
X"59575b58",
X"56831533",
X"5372802e",
X"80f33873",
X"33537a73",
X"2e098106",
X"80e73881",
X"14335379",
X"732e0981",
X"0680da38",
X"80557481",
X"c42983cb",
X"88057033",
X"831b3358",
X"55537376",
X"2e098106",
X"8a388113",
X"33527351",
X"ff9c3f81",
X"157081ff",
X"0656538f",
X"7527d338",
X"800b83cb",
X"80197008",
X"56545573",
X"752e9138",
X"72518414",
X"0853722d",
X"83c08008",
X"81ff0655",
X"800b8318",
X"347453a0",
X"39811681",
X"c41981c4",
X"1781c417",
X"81c41d81",
X"c41c5c5d",
X"57575956",
X"8f7625fe",
X"e8388053",
X"7283c080",
X"0c8c3d0d",
X"04f83d0d",
X"02ae0522",
X"7d595780",
X"56815580",
X"54865381",
X"80527a51",
X"f5953f83",
X"c0800881",
X"ff0683c0",
X"800c8a3d",
X"0d04f73d",
X"0d02b205",
X"22028405",
X"b7053360",
X"5a5b5780",
X"56825579",
X"54865381",
X"80527b51",
X"f4e53f83",
X"c0800881",
X"ff0683c0",
X"800c8b3d",
X"0d04f83d",
X"0d02af05",
X"33598058",
X"80578056",
X"80557854",
X"89538052",
X"7a51f4bb",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8a3d0d04",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002bd9",
X"00002c1a",
X"00002c3c",
X"00002c5e",
X"00002c84",
X"00002c84",
X"00002c84",
X"00002c84",
X"00002cf5",
X"00002d4a",
X"00002d4a",
X"00002d8a",
X"000042ed",
X"00004b31",
X"00004bea",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3f00",
X"0c0c4000",
X"0a0a4100",
X"0b0b4100",
X"07074100",
X"0a0b4300",
X"080b4200",
X"04044500",
X"05054400",
X"06060004",
X"08080004",
X"09090004",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"00005876",
X"00005b7d",
X"00005989",
X"00005b7d",
X"000059c6",
X"00005a17",
X"00005a56",
X"00005a5f",
X"00005b7d",
X"00005b7d",
X"00005b7d",
X"00005b7d",
X"00005a68",
X"00005a70",
X"00005a77",
X"00005c7d",
X"00005d76",
X"00005e8a",
X"00006180",
X"0000619b",
X"00006187",
X"0000619b",
X"000061a2",
X"000061ad",
X"000061b4",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"43505520",
X"54757262",
X"6f3a2564",
X"78000000",
X"44726976",
X"65205475",
X"72626f3a",
X"25730000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"4c6f6164",
X"206d656d",
X"6f727900",
X"53617665",
X"206d656d",
X"6f727920",
X"28666f72",
X"20646562",
X"75676769",
X"6e672900",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"66726565",
X"7a65722e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"4d454d00",
X"5374616e",
X"64617264",
X"00000000",
X"46617374",
X"28362900",
X"46617374",
X"28352900",
X"46617374",
X"28342900",
X"46617374",
X"28332900",
X"46617374",
X"28322900",
X"46617374",
X"28312900",
X"46617374",
X"28302900",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00006df8",
X"00006dfc",
X"00006e04",
X"00006e10",
X"00006e1c",
X"00006e28",
X"00006e34",
X"00006e38",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00000028",
X"00000006",
X"00000005",
X"00000004",
X"00000003",
X"00000002",
X"00000001",
X"00000000",
X"00006f04",
X"00006f10",
X"00006f18",
X"00006f20",
X"00006f28",
X"00006f30",
X"00006f38",
X"00006f40",
X"00006d90",
X"00006be4",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"69383030",
X"00000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
