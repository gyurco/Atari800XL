END; 
