
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81ea",
X"e0738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81f3",
X"cc0c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757580f7",
X"802d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7580f6bf",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80e0ce04",
X"fd3d0d75",
X"705254ae",
X"aa3f83c0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"c0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83c0",
X"8008732e",
X"a13883c0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183c0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83c2d008",
X"248a38b4",
X"fb3fff0b",
X"83c2d00c",
X"800b83c0",
X"800c04ff",
X"3d0d7352",
X"83c0ac08",
X"722e8d38",
X"d93f7151",
X"96a03f71",
X"83c0ac0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"55805681",
X"54bc1508",
X"762e0981",
X"06819138",
X"7451c83f",
X"7958757a",
X"2580f738",
X"83c38008",
X"70892a57",
X"83ff0678",
X"84807231",
X"56565773",
X"78258338",
X"73557583",
X"c2d0082e",
X"8438ff82",
X"3f83c2d0",
X"088025a6",
X"3875892b",
X"5198dc3f",
X"83c38008",
X"8f3dfc11",
X"555c5481",
X"52f81b51",
X"96c63f76",
X"1483c380",
X"0c7583c2",
X"d00c7453",
X"76527851",
X"b3a53f83",
X"c0800883",
X"c3800816",
X"83c3800c",
X"78763176",
X"1b5b5956",
X"778024ff",
X"8b38617a",
X"710c5475",
X"5475802e",
X"83388154",
X"7383c080",
X"0c8e3d0d",
X"04fc3d0d",
X"fe943f76",
X"51fea83f",
X"863dfc05",
X"53785277",
X"5195e93f",
X"7975710c",
X"5483c080",
X"085483c0",
X"8008802e",
X"83388154",
X"7383c080",
X"0c863d0d",
X"04fe3d0d",
X"7583c2d0",
X"08535380",
X"72248938",
X"71732e84",
X"38fdcf3f",
X"7451fde3",
X"3f725197",
X"ae3f83c0",
X"80085283",
X"c0800880",
X"2e833881",
X"527183c0",
X"800c843d",
X"0d04803d",
X"0d7280c0",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"3d0d72bc",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"c40b83c0",
X"800c04fd",
X"3d0d7577",
X"71547053",
X"5553a9fb",
X"3f82c813",
X"08bc150c",
X"82c01308",
X"80c0150c",
X"fce43f73",
X"5193ab3f",
X"7383c0ac",
X"0c83c080",
X"085383c0",
X"8008802e",
X"83388153",
X"7283c080",
X"0c853d0d",
X"04fd3d0d",
X"75775553",
X"fcb83f72",
X"802ea538",
X"bc130852",
X"7351a985",
X"3f83c080",
X"088f3877",
X"527251ff",
X"9a3f83c0",
X"8008538a",
X"3982cc13",
X"0853d839",
X"81537283",
X"c0800c85",
X"3d0d04fe",
X"3d0dff0b",
X"83c2d00c",
X"7483c0b0",
X"0c7583c2",
X"cc0cafd9",
X"3f83c080",
X"0881ff06",
X"52815371",
X"993883c2",
X"e8518e94",
X"3f83c080",
X"085283c0",
X"8008802e",
X"83387252",
X"71537283",
X"c0800c84",
X"3d0d04fa",
X"3d0d787a",
X"82c41208",
X"82c41208",
X"70722459",
X"56565757",
X"73732e09",
X"81069138",
X"80c01652",
X"80c01751",
X"a6f63f83",
X"c0800855",
X"7483c080",
X"0c883d0d",
X"04f63d0d",
X"7c5b807b",
X"715c5457",
X"7a772e8c",
X"38811a82",
X"cc140854",
X"5a72f638",
X"805980d9",
X"397a5481",
X"5780707b",
X"7b315a57",
X"55ff1853",
X"74732580",
X"c13882cc",
X"14085273",
X"51ff8c3f",
X"800b83c0",
X"800825a1",
X"3882cc14",
X"0882cc11",
X"0882cc16",
X"0c7482cc",
X"120c5375",
X"802e8638",
X"7282cc17",
X"0c725480",
X"577382cc",
X"15088117",
X"575556ff",
X"b8398119",
X"59800bff",
X"1b545478",
X"73258338",
X"81547681",
X"32707506",
X"515372ff",
X"90388c3d",
X"0d04f73d",
X"0d7b7d5a",
X"5a82d052",
X"83c2cc08",
X"5180e5bb",
X"3f83c080",
X"0857f9da",
X"3f795283",
X"c2d45195",
X"b73f83c0",
X"80085480",
X"5383c080",
X"08732e09",
X"81068283",
X"3883c0b0",
X"080b0b81",
X"effc5370",
X"5256a6b3",
X"3f0b0b81",
X"effc5280",
X"c01651a6",
X"a63f75bc",
X"170c7382",
X"c0170c81",
X"0b82c417",
X"0c810b82",
X"c8170c73",
X"82cc170c",
X"ff1782d0",
X"17555781",
X"913983c0",
X"bc337082",
X"2a708106",
X"51545572",
X"81803874",
X"812a8106",
X"587780f6",
X"3874842a",
X"810682c4",
X"150c83c0",
X"bc338106",
X"82c8150c",
X"79527351",
X"a5cd3f73",
X"51a5e43f",
X"83c08008",
X"1453af73",
X"70810555",
X"3472bc15",
X"0c83c0bd",
X"527251a5",
X"ae3f83c0",
X"b40882c0",
X"150c83c0",
X"ca5280c0",
X"1451a59b",
X"3f78802e",
X"8d387351",
X"782d83c0",
X"8008802e",
X"99387782",
X"cc150c75",
X"802e8638",
X"7382cc17",
X"0c7382d0",
X"15ff1959",
X"55567680",
X"2e9b3883",
X"c0b45283",
X"c2d45194",
X"ad3f83c0",
X"80088a38",
X"83c0bd33",
X"5372fed2",
X"3878802e",
X"893883c0",
X"b00851fc",
X"b83f83c0",
X"b0085372",
X"83c0800c",
X"8b3d0d04",
X"ff3d0d80",
X"527351fd",
X"b53f833d",
X"0d04f03d",
X"0d627052",
X"54f6893f",
X"83c08008",
X"7453873d",
X"70535555",
X"f6a93ff7",
X"893f7351",
X"d33f6353",
X"745283c0",
X"800851fa",
X"b83f923d",
X"0d047183",
X"c0800c04",
X"80c01283",
X"c0800c04",
X"803d0d72",
X"82c01108",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"7282cc11",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d7282c4",
X"110883c0",
X"800c5182",
X"3d0d04f9",
X"3d0d7983",
X"c0900857",
X"57817727",
X"81963876",
X"88170827",
X"818e3875",
X"33557482",
X"2e893874",
X"832eb338",
X"80fe3974",
X"54761083",
X"fe065376",
X"882a8c17",
X"08055289",
X"3dfc0551",
X"aa873f83",
X"c0800880",
X"df38029d",
X"0533893d",
X"3371882b",
X"07565680",
X"d1398454",
X"76822b83",
X"fc065376",
X"872a8c17",
X"08055289",
X"3dfc0551",
X"a9d73f83",
X"c08008b0",
X"38029f05",
X"33028405",
X"9e053371",
X"982b7190",
X"2b07028c",
X"059d0533",
X"70882b72",
X"078d3d33",
X"7180ffff",
X"fe800607",
X"51525357",
X"58568339",
X"81557483",
X"c0800c89",
X"3d0d04fb",
X"3d0d83c0",
X"9008fe19",
X"881208fe",
X"05555654",
X"80567473",
X"278d3882",
X"14337571",
X"29941608",
X"05575375",
X"83c0800c",
X"873d0d04",
X"fc3d0d76",
X"52800b83",
X"c0900870",
X"33515253",
X"70832e09",
X"81069138",
X"95123394",
X"13337198",
X"2b71902b",
X"07555551",
X"9b12339a",
X"13337188",
X"2b077407",
X"83c0800c",
X"55863d0d",
X"04fc3d0d",
X"7683c090",
X"08555580",
X"75238815",
X"08537281",
X"2e883888",
X"14087326",
X"85388152",
X"b2397290",
X"38733352",
X"71832e09",
X"81068538",
X"90140853",
X"728c160c",
X"72802e8d",
X"387251fe",
X"d63f83c0",
X"80085285",
X"39901408",
X"52719016",
X"0c805271",
X"83c0800c",
X"863d0d04",
X"fa3d0d78",
X"83c09008",
X"71228105",
X"7083ffff",
X"06575457",
X"5573802e",
X"88389015",
X"08537286",
X"38835280",
X"e739738f",
X"06527180",
X"da388113",
X"90160c8c",
X"15085372",
X"9038830b",
X"84172257",
X"52737627",
X"80c638bf",
X"39821633",
X"ff057484",
X"2a065271",
X"b2387251",
X"fcb13f81",
X"527183c0",
X"800827a8",
X"38835283",
X"c0800888",
X"1708279c",
X"3883c080",
X"088c160c",
X"83c08008",
X"51fdbc3f",
X"83c08008",
X"90160c73",
X"75238052",
X"7183c080",
X"0c883d0d",
X"04f23d0d",
X"60626458",
X"5e5b7533",
X"5574a02e",
X"09810688",
X"38811670",
X"4456ef39",
X"62703356",
X"5674af2e",
X"09810684",
X"38811643",
X"800b881c",
X"0c627033",
X"5155749f",
X"2691387a",
X"51fdd23f",
X"83c08008",
X"56807d34",
X"83813993",
X"3d841c08",
X"7058595f",
X"8a55a076",
X"70810558",
X"34ff1555",
X"74ff2e09",
X"8106ef38",
X"80705a5c",
X"887f085f",
X"5a7b811d",
X"7081ff06",
X"60137033",
X"70af3270",
X"30a07327",
X"71802507",
X"5151525b",
X"535e5755",
X"7480e738",
X"76ae2e09",
X"81068338",
X"8155787a",
X"27750755",
X"74802e9f",
X"38798832",
X"703078ae",
X"32703070",
X"73079f2a",
X"53515751",
X"5675bb38",
X"88598b5a",
X"ffab3976",
X"982b5574",
X"80258738",
X"81e9f017",
X"3357ff9f",
X"17557499",
X"268938e0",
X"177081ff",
X"06585578",
X"811a7081",
X"ff06721b",
X"535b5755",
X"767534fe",
X"f8397b1e",
X"7f0c8055",
X"76a02683",
X"38815574",
X"8b19347a",
X"51fc823f",
X"83c08008",
X"80f538a0",
X"547a2270",
X"852b83e0",
X"06545590",
X"1b08527c",
X"51a4923f",
X"83c08008",
X"5783c080",
X"08818138",
X"7c335574",
X"802e80f4",
X"388b1d33",
X"70832a70",
X"81065156",
X"5674b438",
X"8b7d841d",
X"0883c080",
X"08595b5b",
X"58ff1858",
X"77ff2e9a",
X"38797081",
X"055b3379",
X"7081055b",
X"33717131",
X"52565675",
X"802ee238",
X"86397580",
X"2e96387a",
X"51fbe53f",
X"ff863983",
X"c0800856",
X"83c08008",
X"b6388339",
X"7656841b",
X"088b1133",
X"515574a7",
X"388b1d33",
X"70842a70",
X"81065156",
X"56748938",
X"83569439",
X"81569039",
X"7c51fa94",
X"3f83c080",
X"08881c0c",
X"fd813975",
X"83c0800c",
X"903d0d04",
X"f83d0d7a",
X"7c595782",
X"5483fe53",
X"77527651",
X"a2d73f83",
X"5683c080",
X"0880ec38",
X"81173377",
X"3371882b",
X"07565682",
X"567482d4",
X"d52e0981",
X"0680d438",
X"7554b653",
X"77527651",
X"a2ab3f83",
X"c0800898",
X"38811733",
X"77337188",
X"2b0783c0",
X"80085256",
X"56748182",
X"c62eac38",
X"825480d2",
X"53775276",
X"51a2823f",
X"83c08008",
X"98388117",
X"33773371",
X"882b0783",
X"c0800852",
X"56567481",
X"82c62e83",
X"38815675",
X"83c0800c",
X"8a3d0d04",
X"eb3d0d67",
X"5a800b83",
X"c0900ca1",
X"a43f83c0",
X"80088106",
X"55825674",
X"83ef3874",
X"75538f3d",
X"70535759",
X"feca3f83",
X"c0800881",
X"ff065776",
X"812e0981",
X"0680d438",
X"905483be",
X"53745275",
X"51a1963f",
X"83c08008",
X"80c9388f",
X"3d335574",
X"802e80c9",
X"3802bf05",
X"33028405",
X"be053371",
X"982b7190",
X"2b07028c",
X"05bd0533",
X"70882b72",
X"07953d33",
X"71077058",
X"7b575e52",
X"5e575957",
X"fdee3f83",
X"c0800881",
X"ff065776",
X"832e0981",
X"06863881",
X"5682f239",
X"76802e86",
X"38865682",
X"e839a454",
X"8d537852",
X"7551a0ad",
X"3f815683",
X"c0800882",
X"d43802be",
X"05330284",
X"05bd0533",
X"71882b07",
X"595d77ab",
X"380280ce",
X"05330284",
X"0580cd05",
X"3371982b",
X"71902b07",
X"973d3370",
X"882b7207",
X"02940580",
X"cb053371",
X"0754525e",
X"57595602",
X"b7053378",
X"71290288",
X"05b60533",
X"028c05b5",
X"05337188",
X"2b07701d",
X"707f8c05",
X"0c5f5957",
X"595d8e3d",
X"33821b34",
X"02b90533",
X"903d3371",
X"882b075a",
X"5c78841b",
X"2302bb05",
X"33028405",
X"ba053371",
X"882b0756",
X"5c74ab38",
X"0280ca05",
X"33028405",
X"80c90533",
X"71982b71",
X"902b0796",
X"3d337088",
X"2b720702",
X"940580c7",
X"05337107",
X"51525357",
X"5e5c7476",
X"31783179",
X"842a903d",
X"33547171",
X"31535656",
X"80d6a03f",
X"83c08008",
X"82057088",
X"1c0c83c0",
X"8008e08a",
X"05565674",
X"83dffe26",
X"83388257",
X"83fff676",
X"27853883",
X"57893986",
X"5676802e",
X"80db3876",
X"7a347683",
X"2e098106",
X"b0380280",
X"d6053302",
X"840580d5",
X"05337198",
X"2b71902b",
X"07993d33",
X"70882b72",
X"07029405",
X"80d30533",
X"71077f90",
X"050c525e",
X"57585686",
X"39771b90",
X"1b0c841a",
X"228c1b08",
X"1971842a",
X"05941c0c",
X"5d800b81",
X"1b347983",
X"c0900c80",
X"567583c0",
X"800c973d",
X"0d04e93d",
X"0d83c090",
X"08568554",
X"75802e81",
X"8238800b",
X"81173499",
X"3de01146",
X"6a548a3d",
X"705458ec",
X"0551f6e5",
X"3f83c080",
X"085483c0",
X"800880df",
X"38893d33",
X"5473802e",
X"913802ab",
X"05337084",
X"2a810651",
X"5574802e",
X"86388354",
X"80c13976",
X"51f4893f",
X"83c08008",
X"a0170c02",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"9c1c0c52",
X"78981b0c",
X"53565957",
X"810b8117",
X"34745473",
X"83c0800c",
X"993d0d04",
X"f53d0d7d",
X"7f617283",
X"c090085a",
X"5d5d595c",
X"807b0c85",
X"5775802e",
X"81e03881",
X"16338106",
X"55845774",
X"802e81d2",
X"38913974",
X"81173486",
X"39800b81",
X"17348157",
X"81c0399c",
X"16089817",
X"08315574",
X"78278338",
X"74587780",
X"2e81a938",
X"98160870",
X"83ff0656",
X"577480cf",
X"38821633",
X"ff057789",
X"2a067081",
X"ff065a55",
X"78a03876",
X"8738a016",
X"08558d39",
X"a4160851",
X"f0e93f83",
X"c0800855",
X"817527ff",
X"a83874a4",
X"170ca416",
X"0851f283",
X"3f83c080",
X"085583c0",
X"8008802e",
X"ff893883",
X"c0800819",
X"a8170c98",
X"160883ff",
X"06848071",
X"31515577",
X"75278338",
X"77557483",
X"ffff0654",
X"98160883",
X"ff0653a8",
X"16085279",
X"577b8338",
X"7b577651",
X"9ad33f83",
X"c08008fe",
X"d0389816",
X"08159817",
X"0c741a78",
X"76317c08",
X"177d0c59",
X"5afed339",
X"80577683",
X"c0800c8d",
X"3d0d04fa",
X"3d0d7883",
X"c0900855",
X"56855573",
X"802e81e3",
X"38811433",
X"81065384",
X"5572802e",
X"81d5389c",
X"14085372",
X"76278338",
X"72569814",
X"0857800b",
X"98150c75",
X"802e81b9",
X"38821433",
X"70892b56",
X"5376802e",
X"b7387452",
X"ff165180",
X"d1a13f83",
X"c08008ff",
X"18765470",
X"53585380",
X"d1913f83",
X"c0800873",
X"26963874",
X"30707806",
X"7098170c",
X"777131a4",
X"17085258",
X"51538939",
X"a0140870",
X"a4160c53",
X"747627b9",
X"387251ee",
X"d63f83c0",
X"80085381",
X"0b83c080",
X"08278b38",
X"88140883",
X"c0800826",
X"8838800b",
X"811534b0",
X"3983c080",
X"08a4150c",
X"98140815",
X"98150c75",
X"753156c4",
X"39981408",
X"16709816",
X"0c735256",
X"efc53f83",
X"c080088c",
X"3883c080",
X"08811534",
X"81559439",
X"821433ff",
X"0576892a",
X"0683c080",
X"0805a815",
X"0c805574",
X"83c0800c",
X"883d0d04",
X"ef3d0d63",
X"56855583",
X"c0900880",
X"2e80d238",
X"933df405",
X"84170c64",
X"53883d70",
X"53765257",
X"f1cf3f83",
X"c0800855",
X"83c08008",
X"b438883d",
X"33547380",
X"2ea13802",
X"a7053370",
X"842a7081",
X"06515555",
X"83557380",
X"2e973876",
X"51eef53f",
X"83c08008",
X"88170c75",
X"51efa63f",
X"83c08008",
X"557483c0",
X"800c933d",
X"0d04e43d",
X"0d6ea13d",
X"08405e85",
X"5683c090",
X"08802e84",
X"85389e3d",
X"f405841f",
X"0c7e9838",
X"7d51eef5",
X"3f83c080",
X"085683ee",
X"39814181",
X"f6398341",
X"81f13993",
X"3d7f9605",
X"4159807f",
X"8295055e",
X"56756081",
X"ff053483",
X"41901e08",
X"762e81d3",
X"38a0547d",
X"2270852b",
X"83e00654",
X"58901e08",
X"52785196",
X"dc3f83c0",
X"80084183",
X"c08008ff",
X"b8387833",
X"5c7b802e",
X"ffb4388b",
X"193370bf",
X"06718106",
X"52435574",
X"802e80de",
X"387b81bf",
X"0655748f",
X"2480d338",
X"9a193355",
X"7480cb38",
X"f31d7058",
X"5d815675",
X"8b2e0981",
X"0685388e",
X"568b3975",
X"9a2e0981",
X"0683389c",
X"56751970",
X"70810552",
X"33713381",
X"1a821a5f",
X"5b525b55",
X"74863879",
X"77348539",
X"80df7734",
X"777b5757",
X"7aa02e09",
X"8106c038",
X"81567b81",
X"e5327030",
X"709f2a51",
X"51557bae",
X"2e933874",
X"802e8e38",
X"61832a70",
X"81065155",
X"74802e97",
X"387d51ed",
X"df3f83c0",
X"80084183",
X"c0800887",
X"38901e08",
X"feaf3880",
X"60347580",
X"2e88387c",
X"527f518e",
X"823f6080",
X"2e863880",
X"0b901f0c",
X"60566083",
X"2e853860",
X"81d03889",
X"1f57901e",
X"08802e81",
X"a8388056",
X"75197033",
X"515574a0",
X"2ea03874",
X"852e0981",
X"06843881",
X"e5557477",
X"70810559",
X"34811670",
X"81ff0657",
X"55877627",
X"d7388819",
X"335574a0",
X"2ea938ae",
X"77708105",
X"59348856",
X"75197033",
X"515574a0",
X"2e953874",
X"77708105",
X"59348116",
X"7081ff06",
X"57558a76",
X"27e2388b",
X"19337f88",
X"05349f19",
X"339e1a33",
X"71982b71",
X"902b079d",
X"1c337088",
X"2b72079c",
X"1e337107",
X"640c5299",
X"1d33981e",
X"3371882b",
X"07535153",
X"57595674",
X"7f840523",
X"97193396",
X"1a337188",
X"2b075656",
X"747f8605",
X"23807734",
X"7d51ebf0",
X"3f83c080",
X"08833270",
X"30707207",
X"9f2c83c0",
X"80080652",
X"5656961f",
X"3355748a",
X"38891f52",
X"961f518c",
X"8e3f7583",
X"c0800c9e",
X"3d0d04f4",
X"3d0d7e8f",
X"3dec1156",
X"56589053",
X"f0155277",
X"51e0d23f",
X"83c08008",
X"80d63878",
X"902e0981",
X"0680cd38",
X"02ab0533",
X"81f3d40b",
X"81f3d433",
X"5758568c",
X"3974762e",
X"8a388417",
X"70335657",
X"74f33876",
X"33705755",
X"74802eac",
X"38821722",
X"708a2b90",
X"3dec0556",
X"70555656",
X"96800a52",
X"7751e081",
X"3f83c080",
X"08863878",
X"752e8538",
X"80568539",
X"81173356",
X"7583c080",
X"0c8e3d0d",
X"04fc3d0d",
X"76705255",
X"8b953f83",
X"c0800815",
X"ff055473",
X"752e8e38",
X"73335372",
X"ae2e8638",
X"ff1454ef",
X"39775281",
X"14518aad",
X"3f83c080",
X"08307083",
X"c0800807",
X"802583c0",
X"800c5386",
X"3d0d04fc",
X"3d0d7670",
X"5255e6ee",
X"3f83c080",
X"08548153",
X"83c08008",
X"80c13874",
X"51e6b13f",
X"83c08008",
X"81f08c53",
X"83c08008",
X"5253ff91",
X"3f83c080",
X"08a13881",
X"f0905272",
X"51ff823f",
X"83c08008",
X"923881f0",
X"94527251",
X"fef33f83",
X"c0800880",
X"2e833881",
X"54735372",
X"83c0800c",
X"863d0d04",
X"fd3d0d75",
X"705254e6",
X"8d3f8153",
X"83c08008",
X"98387351",
X"e5d63f83",
X"c3980852",
X"83c08008",
X"51feba3f",
X"83c08008",
X"537283c0",
X"800c853d",
X"0d04df3d",
X"0da43d08",
X"70525edb",
X"f43f83c0",
X"80083395",
X"3d565473",
X"963881f7",
X"a4527451",
X"898d3f9a",
X"397d5278",
X"51defc3f",
X"84d0397d",
X"51dbda3f",
X"83c08008",
X"527451db",
X"8a3f8043",
X"80428041",
X"804083c3",
X"a0085294",
X"3d70525d",
X"e1e43f83",
X"c0800859",
X"800b83c0",
X"8008555b",
X"83c08008",
X"7b2e9438",
X"811b7452",
X"5be4e63f",
X"83c08008",
X"5483c080",
X"08ee3880",
X"5aff5f79",
X"09709f2c",
X"7b065b54",
X"7a7a2484",
X"38ff1b5a",
X"f61a7009",
X"709f2c72",
X"067bff12",
X"5a5a5255",
X"55807525",
X"95387651",
X"e4ab3f83",
X"c0800876",
X"ff185855",
X"57738024",
X"ed38747f",
X"2e8638a1",
X"b53f745f",
X"78ff1b70",
X"585d5880",
X"7a259538",
X"7751e481",
X"3f83c080",
X"0876ff18",
X"58555873",
X"8024ed38",
X"800b83c7",
X"d00c800b",
X"83c8880c",
X"81f09851",
X"8d8c3f81",
X"800b83c8",
X"880c81f0",
X"a0518cfe",
X"3fa80b83",
X"c7d00c76",
X"802e80e4",
X"3883c7d0",
X"08777932",
X"70307072",
X"07802570",
X"872b83c8",
X"880c5156",
X"78535656",
X"e3b83f83",
X"c0800880",
X"2e883881",
X"f0a8518c",
X"c53f7651",
X"e2fa3f83",
X"c0800852",
X"81f28851",
X"8cb43f76",
X"51e3823f",
X"83c08008",
X"83c7d008",
X"55577574",
X"258638a8",
X"1656f739",
X"7583c7d0",
X"0c86f076",
X"24ff9838",
X"87980b83",
X"c7d00c77",
X"802eb138",
X"7751e2b8",
X"3f83c080",
X"08785255",
X"e2d83f81",
X"f0b05483",
X"c080088d",
X"38873980",
X"763481d0",
X"3981f0ac",
X"54745373",
X"5281f080",
X"518bd33f",
X"805481f0",
X"88518bca",
X"3f811454",
X"73a82e09",
X"8106ef38",
X"868da051",
X"9da83f80",
X"52903d70",
X"525780c7",
X"8e3f8352",
X"765180c7",
X"863f6281",
X"8f386180",
X"2e80fb38",
X"7b5473ff",
X"2e963878",
X"802e818a",
X"387851e1",
X"dc3f83c0",
X"8008ff15",
X"5559e739",
X"78802e80",
X"f5387851",
X"e1d83f83",
X"c0800880",
X"2efc8e38",
X"7851e1a0",
X"3f83c080",
X"085281ef",
X"fc5183e0",
X"3f83c080",
X"08a3387c",
X"5185983f",
X"83c08008",
X"5574ff16",
X"56548074",
X"25ae3874",
X"1d703355",
X"5673af2e",
X"fecd38e9",
X"397851e0",
X"e13f83c0",
X"8008527c",
X"5184d03f",
X"8f397f88",
X"29601005",
X"7a056105",
X"5afc9039",
X"62802efb",
X"d1388052",
X"765180c5",
X"e63fa33d",
X"0d04803d",
X"0d9088b8",
X"337081ff",
X"0670842a",
X"81327081",
X"06515151",
X"5170802e",
X"8d38a80b",
X"9088b834",
X"b80b9088",
X"b8347083",
X"c0800c82",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067085",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d3898",
X"0b9088b8",
X"34b80b90",
X"88b83470",
X"83c0800c",
X"823d0d04",
X"930b9088",
X"bc34ff0b",
X"9088a834",
X"04ff3d0d",
X"028f0533",
X"52800b90",
X"88bc348a",
X"519aef3f",
X"df3f80f8",
X"0b9088a0",
X"34800b90",
X"888834fa",
X"12527190",
X"88803480",
X"0b908898",
X"34719088",
X"90349088",
X"b8528072",
X"34b87234",
X"833d0d04",
X"803d0d02",
X"8b053351",
X"709088b4",
X"34febf3f",
X"83c08008",
X"802ef638",
X"823d0d04",
X"803d0d84",
X"39a8de3f",
X"fed93f83",
X"c0800880",
X"2ef33890",
X"88b43370",
X"81ff0683",
X"c0800c51",
X"823d0d04",
X"803d0da3",
X"0b9088bc",
X"34ff0b90",
X"88a83490",
X"88b851a8",
X"7134b871",
X"34823d0d",
X"04803d0d",
X"9088bc33",
X"70982b70",
X"802583c0",
X"800c5151",
X"823d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"832a8132",
X"70810651",
X"51515170",
X"802ee838",
X"b00b9088",
X"b834b80b",
X"9088b834",
X"823d0d04",
X"803d0d90",
X"80ac0881",
X"0683c080",
X"0c823d0d",
X"04fd3d0d",
X"75775454",
X"80732594",
X"38737081",
X"05553352",
X"81f0b451",
X"87843fff",
X"1353e939",
X"853d0d04",
X"fd3d0d75",
X"77535473",
X"33517089",
X"38713351",
X"70802ea1",
X"38733372",
X"33525372",
X"71278538",
X"ff519439",
X"70732785",
X"3881518b",
X"39811481",
X"135354d3",
X"39805170",
X"83c0800c",
X"853d0d04",
X"fd3d0d75",
X"77545472",
X"337081ff",
X"06525270",
X"802ea338",
X"7181ff06",
X"8114ffbf",
X"12535452",
X"70992689",
X"38a01270",
X"81ff0653",
X"51717470",
X"81055634",
X"d2398074",
X"34853d0d",
X"04ffbd3d",
X"0d80c63d",
X"0852a53d",
X"705254ff",
X"b33f80c7",
X"3d085285",
X"3d705253",
X"ffa63f72",
X"527351fe",
X"df3f80c5",
X"3d0d04fe",
X"3d0d7476",
X"53537170",
X"81055333",
X"51707370",
X"81055534",
X"70f03884",
X"3d0d04fe",
X"3d0d7452",
X"80723352",
X"5370732e",
X"8d388112",
X"81147133",
X"53545270",
X"f5387283",
X"c0800c84",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"bdf93f83",
X"c080087a",
X"27ee3874",
X"802e80dd",
X"38745275",
X"51bde43f",
X"83c08008",
X"75537652",
X"54bde83f",
X"83c08008",
X"7a537552",
X"56bdcc3f",
X"83c08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"c08008c5",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9f",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fc813f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd53f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbb13f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83c0940c",
X"7183c098",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383c094",
X"085283c0",
X"980851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"bdbe5351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fc3d",
X"0d765574",
X"83c3ac08",
X"2eaf3880",
X"53745187",
X"c13f83c0",
X"800881ff",
X"06ff1470",
X"81ff0672",
X"30709f2a",
X"51525553",
X"5472802e",
X"843871dd",
X"3873fe38",
X"7483c3ac",
X"0c863d0d",
X"04ff3d0d",
X"ff0b83c3",
X"ac0c84a5",
X"3f815187",
X"853f83c0",
X"800881ff",
X"065271ee",
X"3881d33f",
X"7183c080",
X"0c833d0d",
X"04fc3d0d",
X"76028405",
X"a2052202",
X"8805a605",
X"227a5455",
X"5555ff82",
X"3f72802e",
X"a03883c3",
X"c0143375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552dd",
X"39800b83",
X"c0800c86",
X"3d0d04fc",
X"3d0d7678",
X"7a115653",
X"55805371",
X"742e9338",
X"72155170",
X"3383c3c0",
X"13348112",
X"81145452",
X"ea39800b",
X"83c0800c",
X"863d0d04",
X"fd3d0d90",
X"5483c3ac",
X"085186f4",
X"3f83c080",
X"0881ff06",
X"ff157130",
X"71307073",
X"079f2a72",
X"9f2a0652",
X"55525553",
X"72db3885",
X"3d0d0480",
X"3d0d83c3",
X"b8081083",
X"c3b00807",
X"9080a80c",
X"823d0d04",
X"800b83c3",
X"b80ce43f",
X"04810b83",
X"c3b80cdb",
X"3f04ed3f",
X"047183c3",
X"b40c0480",
X"3d0d8051",
X"f43f810b",
X"83c3b80c",
X"810b83c3",
X"b00cffbb",
X"3f823d0d",
X"04803d0d",
X"72307074",
X"07802583",
X"c3b00c51",
X"ffa53f82",
X"3d0d0480",
X"3d0d028b",
X"05339080",
X"a40c9080",
X"a8087081",
X"06515170",
X"f5389080",
X"a4087081",
X"ff0683c0",
X"800c5182",
X"3d0d0480",
X"3d0d81ff",
X"51d13f83",
X"c0800881",
X"ff0683c0",
X"800c823d",
X"0d04803d",
X"0d73902b",
X"73079080",
X"b40c823d",
X"0d0404fb",
X"3d0d7802",
X"84059f05",
X"3370982b",
X"55575572",
X"80259b38",
X"7580ff06",
X"56805280",
X"f751e03f",
X"83c08008",
X"81ff0654",
X"73812680",
X"ff388051",
X"fee73fff",
X"a23f8151",
X"fedf3fff",
X"9a3f7551",
X"feed3f74",
X"982a51fe",
X"e63f7490",
X"2a7081ff",
X"065253fe",
X"da3f7488",
X"2a7081ff",
X"065253fe",
X"ce3f7481",
X"ff0651fe",
X"c63f8155",
X"7580c02e",
X"09810686",
X"38819555",
X"8d397580",
X"c82e0981",
X"06843881",
X"87557451",
X"fea53f8a",
X"55fec83f",
X"83c08008",
X"81ff0670",
X"982b5454",
X"7280258c",
X"38ff1570",
X"81ff0656",
X"5374e238",
X"7383c080",
X"0c873d0d",
X"04fa3d0d",
X"fdc53f80",
X"51fdda3f",
X"8a54fe93",
X"3fff1470",
X"81ff0655",
X"5373f338",
X"73745355",
X"80c051fe",
X"a63f83c0",
X"800881ff",
X"06547381",
X"2e098106",
X"829f3883",
X"aa5280c8",
X"51fe8c3f",
X"83c08008",
X"81ff0653",
X"72812e09",
X"810681a8",
X"38745487",
X"3d741154",
X"56fdc83f",
X"83c08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e53802",
X"9a053353",
X"72812e09",
X"810681d9",
X"38029b05",
X"335380ce",
X"90547281",
X"aa2e8d38",
X"81c73980",
X"e4518b9a",
X"3fff1454",
X"73802e81",
X"b838820a",
X"5281e951",
X"fda53f83",
X"c0800881",
X"ff065372",
X"de387252",
X"80fa51fd",
X"923f83c0",
X"800881ff",
X"06537281",
X"90387254",
X"731653fc",
X"d63f83c0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e8",
X"38873d33",
X"70862a70",
X"81065154",
X"548c5572",
X"80e33884",
X"5580de39",
X"745281e9",
X"51fccc3f",
X"83c08008",
X"81ff0653",
X"825581e9",
X"56817327",
X"86387355",
X"80c15680",
X"ce90548a",
X"3980e451",
X"8a8c3fff",
X"14547380",
X"2ea93880",
X"527551fc",
X"9a3f83c0",
X"800881ff",
X"065372e1",
X"38848052",
X"80d051fc",
X"863f83c0",
X"800881ff",
X"06537280",
X"2e833880",
X"557483c3",
X"bc348051",
X"fb873ffb",
X"c23f883d",
X"0d04fb3d",
X"0d775480",
X"0b83c3bc",
X"3370832a",
X"70810651",
X"55575572",
X"752e0981",
X"06853873",
X"892b5473",
X"5280d151",
X"fbbd3f83",
X"c0800881",
X"ff065372",
X"bd3882b8",
X"c054fb83",
X"3f83c080",
X"0881ff06",
X"537281ff",
X"2e098106",
X"8938ff14",
X"5473e738",
X"9f397281",
X"fe2e0981",
X"06963883",
X"c7c05283",
X"c3c051fa",
X"ed3ffad3",
X"3ffad03f",
X"83398155",
X"8051fa89",
X"3ffac43f",
X"7481ff06",
X"83c0800c",
X"873d0d04",
X"fb3d0d77",
X"83c3c056",
X"548151f9",
X"ec3f83c3",
X"bc337083",
X"2a708106",
X"51545672",
X"85387389",
X"2b547352",
X"80d851fa",
X"b63f83c0",
X"800881ff",
X"06537280",
X"e43881ff",
X"51f9d43f",
X"81fe51f9",
X"ce3f8480",
X"53747081",
X"05563351",
X"f9c13fff",
X"137083ff",
X"ff065153",
X"72eb3872",
X"51f9b03f",
X"7251f9ab",
X"3ff9d03f",
X"83c08008",
X"9f0653a7",
X"88547285",
X"2e8c3899",
X"3980e451",
X"87c43fff",
X"1454f9b3",
X"3f83c080",
X"0881ff2e",
X"843873e9",
X"388051f8",
X"e43ff99f",
X"3f800b83",
X"c0800c87",
X"3d0d0471",
X"83c7c40c",
X"8880800b",
X"83c7c00c",
X"8480800b",
X"83c7c80c",
X"04fd3d0d",
X"77701755",
X"7705ff1a",
X"535371ff",
X"2e943873",
X"70810555",
X"33517073",
X"70810555",
X"34ff1252",
X"e939853d",
X"0d04fb3d",
X"0d87a681",
X"0b83c7c4",
X"08565675",
X"3383a680",
X"1634a054",
X"83a08053",
X"83c7c408",
X"5283c7c0",
X"0851ffb1",
X"3fa05483",
X"a4805383",
X"c7c40852",
X"83c7c008",
X"51ff9e3f",
X"905483a8",
X"805383c7",
X"c4085283",
X"c7c00851",
X"ff8b3fa0",
X"53805283",
X"c7c80883",
X"a0800551",
X"86953fa0",
X"53805283",
X"c7c80883",
X"a4800551",
X"86853f90",
X"53805283",
X"c7c80883",
X"a8800551",
X"85f53fff",
X"763483a0",
X"80548053",
X"83c7c408",
X"5283c7c8",
X"0851fec5",
X"3f80d080",
X"5483b080",
X"5383c7c4",
X"085283c7",
X"c80851fe",
X"b03f87ba",
X"3fa25480",
X"5383c7c8",
X"088c8005",
X"5281f4c8",
X"51fe9a3f",
X"860b87a8",
X"8334800b",
X"87a88234",
X"800b87a0",
X"9a34af0b",
X"87a09634",
X"bf0b87a0",
X"9734800b",
X"87a09834",
X"9f0b87a0",
X"9934800b",
X"87a09b34",
X"e00b87a8",
X"8934a20b",
X"87a88034",
X"830b87a4",
X"8f34820b",
X"87a88134",
X"873d0d04",
X"fc3d0d83",
X"a0805480",
X"5383c7c8",
X"085283c7",
X"c40851fd",
X"b83f80d0",
X"805483b0",
X"805383c7",
X"c8085283",
X"c7c40851",
X"fda33fa0",
X"5483a080",
X"5383c7c8",
X"085283c7",
X"c40851fd",
X"903fa054",
X"83a48053",
X"83c7c808",
X"5283c7c4",
X"0851fcfd",
X"3f905483",
X"a8805383",
X"c7c80852",
X"83c7c408",
X"51fcea3f",
X"83c7c408",
X"5583a680",
X"153387a6",
X"8134863d",
X"0d04fa3d",
X"0d787052",
X"55c1e33f",
X"83ffff0b",
X"83c08008",
X"25a93874",
X"51c1e43f",
X"83c08008",
X"9e3883c0",
X"80085788",
X"3dfc0554",
X"84808053",
X"83c7c408",
X"527451ff",
X"bf963fff",
X"bedc3f88",
X"3d0d04fa",
X"3d0d7870",
X"5255c1a2",
X"3f83ffff",
X"0b83c080",
X"08259638",
X"8057883d",
X"fc055484",
X"80805383",
X"c7c40852",
X"7451c095",
X"3f883d0d",
X"04803d0d",
X"90809008",
X"810683c0",
X"800c823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087081",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fd0676",
X"1007720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870822c",
X"bf0683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe830676",
X"822b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087088",
X"2c870683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f1ff06",
X"76882b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"912cbf06",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fc87",
X"ffff0676",
X"912b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087099",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70ffbf0a",
X"0676992b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90808008",
X"70882c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"0870892c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708a",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8b2c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708c2cbf",
X"0683c080",
X"0c51823d",
X"0d04fe3d",
X"0d7481e6",
X"29872a90",
X"80a00c84",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70810554",
X"34ff1151",
X"f039843d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"8405540c",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"84808053",
X"80528880",
X"0a51ffb3",
X"3f818080",
X"53805282",
X"800a51c6",
X"3f843d0d",
X"04803d0d",
X"8151fcaa",
X"3f72802e",
X"90388051",
X"fdfe3fcd",
X"3f83c7cc",
X"3351fdf4",
X"3f8151fc",
X"bb3f8051",
X"fcb63f80",
X"51fc873f",
X"823d0d04",
X"fd3d0d75",
X"52805480",
X"ff722588",
X"38810bff",
X"80135354",
X"ffbf1251",
X"70992686",
X"38e01252",
X"b039ff9f",
X"12519971",
X"27a738d0",
X"12e01354",
X"51708926",
X"85387252",
X"9839728f",
X"26853872",
X"528f3971",
X"ba2e0981",
X"0685389a",
X"52833980",
X"5273802e",
X"85388180",
X"12527181",
X"ff0683c0",
X"800c853d",
X"0d04803d",
X"0d84d8c0",
X"51807170",
X"81055334",
X"7084e0c0",
X"2e098106",
X"f038823d",
X"0d04fe3d",
X"0d029705",
X"3351fef4",
X"3f83c080",
X"0881ff06",
X"83c7d008",
X"54528073",
X"249b3883",
X"c8840813",
X"7283c888",
X"08075353",
X"71733483",
X"c7d00881",
X"0583c7d0",
X"0c843d0d",
X"04fa3d0d",
X"82800a1b",
X"55805788",
X"3dfc0554",
X"79537452",
X"7851ffba",
X"ac3f883d",
X"0d04fe3d",
X"0d83c7e8",
X"08527451",
X"c1903f83",
X"c080088c",
X"38765375",
X"5283c7e8",
X"0851c63f",
X"843d0d04",
X"fe3d0d83",
X"c7e80853",
X"75527451",
X"ffbbce3f",
X"83c08008",
X"8d387753",
X"765283c7",
X"e80851ff",
X"a03f843d",
X"0d04f73d",
X"0daa8f3f",
X"83c08008",
X"81ff06ff",
X"05577683",
X"38815780",
X"fed13f83",
X"c0800883",
X"c0800856",
X"5a871533",
X"5473802e",
X"80df3874",
X"0881ec9c",
X"2e098106",
X"80d33880",
X"0b911633",
X"55597379",
X"2e80c638",
X"74569a16",
X"33547383",
X"2e098106",
X"a438a416",
X"70335558",
X"80527351",
X"a7f93f80",
X"53805273",
X"51a8993f",
X"81145476",
X"74258338",
X"80547378",
X"34811980",
X"d8179117",
X"33565759",
X"78742e09",
X"8106ffbe",
X"3881c415",
X"98c01b55",
X"5574742e",
X"098106ff",
X"88388b3d",
X"0d04f63d",
X"0d80fdc3",
X"3f83c080",
X"087d83c0",
X"80085859",
X"5b7783c7",
X"d00c8716",
X"33557480",
X"2e81a738",
X"75085473",
X"81efd42e",
X"09810693",
X"38901633",
X"53871633",
X"5281f0bc",
X"51e8f33f",
X"81883973",
X"81ec9c2e",
X"09810680",
X"fd387452",
X"81f0d051",
X"e8dc3f80",
X"70911833",
X"565b5973",
X"792e80e6",
X"38a41657",
X"f6173355",
X"79802e91",
X"38ff1554",
X"73822689",
X"38a81870",
X"83c7d00c",
X"5874812e",
X"09810687",
X"3881f0d8",
X"518d3974",
X"822e0981",
X"068a3881",
X"f0e051e8",
X"953f9539",
X"74832e09",
X"81068f38",
X"76338105",
X"5281f0ec",
X"51e7ff3f",
X"815a8119",
X"80d81891",
X"18335658",
X"5978742e",
X"098106ff",
X"9f38a818",
X"81c41798",
X"c01d5657",
X"5875742e",
X"098106fe",
X"b8388c3d",
X"0d04fe3d",
X"0d83c7e8",
X"0851ffb7",
X"c13f83c0",
X"80088180",
X"802e0981",
X"06883883",
X"c1808053",
X"9c3983c7",
X"e80851ff",
X"b7a43f83",
X"c0800880",
X"d0802e09",
X"81069338",
X"83c1b080",
X"5383c080",
X"085283c7",
X"e80851fb",
X"d43f843d",
X"0d04803d",
X"0df6fc3f",
X"83c08008",
X"842981f4",
X"ec057008",
X"83c0800c",
X"51823d0d",
X"04ed3d0d",
X"80448043",
X"80428041",
X"80705a5b",
X"facc3f80",
X"0b83c7d0",
X"0c800b83",
X"c8880c81",
X"f1c051e6",
X"c53f8180",
X"0b83c888",
X"0c81f1c4",
X"51e6b73f",
X"80d00b83",
X"c7d00c78",
X"30707a07",
X"80257087",
X"2b83c888",
X"0c5155f5",
X"ed3f83c0",
X"80085281",
X"f1cc51e6",
X"913f80f8",
X"0b83c7d0",
X"0c788132",
X"70307072",
X"07802570",
X"872b83c8",
X"880c5156",
X"569e8a3f",
X"83c08008",
X"5281f1dc",
X"51e5e73f",
X"81a00b83",
X"c7d00c78",
X"82327030",
X"70720780",
X"2570872b",
X"83c8880c",
X"515656fe",
X"c53f83c0",
X"80085281",
X"f1ec51e5",
X"bd3f81c8",
X"0b83c7d0",
X"0c788332",
X"70307072",
X"07802570",
X"872b83c8",
X"880c5156",
X"83c7e808",
X"5256ffb2",
X"983f83c0",
X"80085281",
X"f1f451e5",
X"8d3f8298",
X"0b83c7d0",
X"0c810b83",
X"c7d45b58",
X"83c7d008",
X"83197a32",
X"70307072",
X"07802570",
X"872b83c8",
X"880c5157",
X"8e3d7055",
X"ff1b5457",
X"57579bcc",
X"3f797084",
X"055b0851",
X"ffb1ce3f",
X"745483c0",
X"80085377",
X"5281f1fc",
X"51e4bf3f",
X"a81783c7",
X"d00c8118",
X"5877852e",
X"098106ff",
X"af3883b8",
X"0b83c7d0",
X"0c788832",
X"70307072",
X"07802570",
X"872b83c8",
X"880c5156",
X"56f4b93f",
X"81f28c55",
X"83c08008",
X"802e8f38",
X"83c7e408",
X"51ffb0f9",
X"3f83c080",
X"08557452",
X"81f29451",
X"e3ec3f83",
X"e00b83c7",
X"d00c7889",
X"32703070",
X"72078025",
X"70872b83",
X"c8880c51",
X"5681f2a0",
X"5256e3ca",
X"3f84b00b",
X"83c7d00c",
X"788a3270",
X"30707207",
X"80257087",
X"2b83c888",
X"0c515681",
X"f2b85256",
X"e3a83f80",
X"0b83c888",
X"0c858051",
X"f9ec3f86",
X"8da051f5",
X"853f8052",
X"913d7052",
X"559eec3f",
X"83527451",
X"9ee53f63",
X"557483a6",
X"38611959",
X"78802585",
X"38745990",
X"398a7925",
X"85388a59",
X"8739788a",
X"26838538",
X"78822b55",
X"81ebf015",
X"0804f2a6",
X"3f83c080",
X"08615755",
X"75812e09",
X"81068938",
X"83c08008",
X"10559039",
X"75ff2e09",
X"81068838",
X"83c08008",
X"812c5590",
X"75258538",
X"90558839",
X"74802483",
X"38815574",
X"51f2803f",
X"82ba399a",
X"a33f83c0",
X"80086105",
X"55748025",
X"85388055",
X"88398775",
X"25833887",
X"5574518e",
X"863f8298",
X"39f1f03f",
X"83c08008",
X"61055574",
X"80258538",
X"80558839",
X"86752583",
X"38865574",
X"51f1e93f",
X"81f63960",
X"87386280",
X"2e81ed38",
X"83c39c08",
X"83c3980c",
X"adec0b83",
X"c3a00c83",
X"c7e80851",
X"d2b43ff9",
X"e13f81d0",
X"39605680",
X"76259838",
X"ad8b0b83",
X"c3a00c83",
X"c7c41570",
X"085255d2",
X"953f7408",
X"52923975",
X"80259238",
X"83c7c415",
X"0851ffae",
X"923f8052",
X"fc1951b8",
X"3962802e",
X"81963883",
X"c7c41570",
X"0883c7d4",
X"08720c83",
X"c7d40cfc",
X"1a705351",
X"558cd33f",
X"83c08008",
X"5680518c",
X"c93f83c0",
X"80085274",
X"5188e23f",
X"75528051",
X"88db3f80",
X"df396055",
X"807525b6",
X"3883c3a8",
X"0883c398",
X"0cadec0b",
X"83c3a00c",
X"83c7e408",
X"51d19f3f",
X"83c7e408",
X"51cec03f",
X"83c08008",
X"81ff0670",
X"5255f0c9",
X"3f74802e",
X"a7388155",
X"ab397480",
X"259e3883",
X"c7e40851",
X"ffad843f",
X"8051f0ad",
X"3f8e3962",
X"802e8938",
X"f5943f84",
X"39628738",
X"7a802ef8",
X"ff388055",
X"7483c080",
X"0c953d0d",
X"04fe3d0d",
X"83c7f451",
X"8183a93f",
X"f0c73f83",
X"c0800880",
X"2e863880",
X"51818a39",
X"f0cc3f83",
X"c0800880",
X"fe38f0ec",
X"3f83c080",
X"08802eb9",
X"388151ee",
X"a93f8051",
X"f0823fea",
X"a13f800b",
X"83c7d00c",
X"f89f3f83",
X"c0800853",
X"ff0b83c7",
X"d00cec94",
X"3f7280cb",
X"3883c7cc",
X"3351efdc",
X"3f7251ed",
X"f93f80c0",
X"39f0943f",
X"83c08008",
X"802eb538",
X"8151ede6",
X"3f8051ef",
X"bf3fe9de",
X"3fad8b0b",
X"83c3a00c",
X"83c7d408",
X"51cfbf3f",
X"ff0b83c7",
X"d00cebd0",
X"3f83c7d4",
X"08528051",
X"86c73f81",
X"51f1863f",
X"843d0d04",
X"fb3d0d80",
X"5283c7f4",
X"5180f2b8",
X"3f800b83",
X"c7cc3490",
X"80805286",
X"84808051",
X"ffafa83f",
X"83c08008",
X"81a03883",
X"c7f00851",
X"8188ee3f",
X"8a993f81",
X"f78c51ff",
X"b3de3f83",
X"c0800855",
X"9c800a54",
X"80c08053",
X"81f2c052",
X"83c08008",
X"51f2d93f",
X"83c7e808",
X"5381f2d0",
X"527451ff",
X"aea73f83",
X"c0800884",
X"38f5e73f",
X"83c7ec08",
X"5381f2dc",
X"527451ff",
X"ae8f3f83",
X"c08008b6",
X"38873dfc",
X"05548480",
X"805386a8",
X"80805283",
X"c7ec0851",
X"ffac9a3f",
X"83c08008",
X"93387584",
X"80802e09",
X"81068938",
X"810b83c7",
X"cc348739",
X"800b83c7",
X"cc3483c7",
X"cc3351ed",
X"d33f8151",
X"efbf3f93",
X"ca3f8151",
X"efb73f81",
X"51fd863f",
X"fa3983c0",
X"8c080283",
X"c08c0cfb",
X"3d0d0281",
X"f2e80b83",
X"c39c0c81",
X"f2ec0b83",
X"c3940c81",
X"f2f00b83",
X"c3a80c81",
X"f2f40b83",
X"c3a40c83",
X"c08c08fc",
X"050c800b",
X"83c7d40b",
X"83c08c08",
X"f8050c83",
X"c08c08f4",
X"050cffac",
X"a23f83c0",
X"80088605",
X"fc0683c0",
X"8c08f005",
X"0c0283c0",
X"8c08f005",
X"08310d83",
X"3d7083c0",
X"8c08f805",
X"08708405",
X"83c08c08",
X"f8050c0c",
X"51ffa8e3",
X"3f83c08c",
X"08f40508",
X"810583c0",
X"8c08f405",
X"0c83c08c",
X"08f40508",
X"882e0981",
X"06ffab38",
X"86948080",
X"51e5fc3f",
X"ff0b83c7",
X"d00c800b",
X"83c8880c",
X"84d8c00b",
X"83c8840c",
X"8151eaa2",
X"3f8151ea",
X"c73f8051",
X"eac23f81",
X"51eae83f",
X"8251eb90",
X"3f8051eb",
X"b83f8051",
X"ebe23f80",
X"d1ae5280",
X"51dae03f",
X"fcc63f83",
X"c08c08fc",
X"05080d80",
X"0b83c080",
X"0c873d0d",
X"83c08c0c",
X"04803d0d",
X"81ff5180",
X"0b83c898",
X"1234ff11",
X"5170f438",
X"823d0d04",
X"ff3d0d73",
X"70335351",
X"81113371",
X"34718112",
X"34833d0d",
X"04ff3d0d",
X"83cab408",
X"a82e0981",
X"068b3883",
X"cacc0883",
X"cab40c87",
X"39a80b83",
X"cab40c83",
X"cab40886",
X"057081ff",
X"065252d0",
X"e83f833d",
X"0d04fb3d",
X"0d777956",
X"56807071",
X"55555271",
X"7525ac38",
X"72167033",
X"70147081",
X"ff065551",
X"51517174",
X"27893881",
X"127081ff",
X"06535171",
X"81147083",
X"ffff0655",
X"52547473",
X"24d63871",
X"83c0800c",
X"873d0d04",
X"fb3d0d77",
X"568939f9",
X"d83f8351",
X"eb903fd1",
X"ef3f83c0",
X"8008802e",
X"ee3883ca",
X"b4088605",
X"7081ff06",
X"5253cff5",
X"3f810b90",
X"88d434f9",
X"b03f8351",
X"eae83f90",
X"88d43370",
X"81ff0655",
X"5373802e",
X"ea387386",
X"2a708106",
X"515372ff",
X"be387398",
X"2b538073",
X"2480de38",
X"d0df3f83",
X"c0800855",
X"83c08008",
X"80cf3874",
X"1675822b",
X"54549088",
X"c0133374",
X"34811555",
X"74852e09",
X"8106e838",
X"753383c8",
X"98348116",
X"3383c899",
X"34821633",
X"83c89a34",
X"83163383",
X"c89b3484",
X"5283c898",
X"51fe933f",
X"83c08008",
X"81ff0684",
X"17335553",
X"72742e87",
X"38fdce3f",
X"fed13980",
X"e451e9da",
X"3f873d0d",
X"04f43d0d",
X"7e605955",
X"805d8075",
X"822b7183",
X"cab8120c",
X"83cad017",
X"5b5b5776",
X"79347777",
X"2e83b738",
X"76527751",
X"ffa6fe3f",
X"8e3dfc05",
X"54905383",
X"caa05277",
X"51ffa6b9",
X"3f7c5675",
X"902e0981",
X"06839338",
X"83caa051",
X"fcde3f83",
X"caa251fc",
X"d73f83ca",
X"a451fcd0",
X"3f7683ca",
X"b00c7751",
X"ffa3fe3f",
X"81f09052",
X"83c08008",
X"51c69e3f",
X"83c08008",
X"812e0981",
X"0680d438",
X"7683cac8",
X"0c820b83",
X"caa034ff",
X"960b83ca",
X"a1347751",
X"ffa6cb3f",
X"83c08008",
X"5583c080",
X"08772588",
X"3883c080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"caa23474",
X"83caa334",
X"7683caa4",
X"34ff800b",
X"83caa534",
X"81903983",
X"caa03383",
X"caa13371",
X"882b0756",
X"5b7483ff",
X"ff2e0981",
X"0680e838",
X"fe800b83",
X"cac80c81",
X"0b83cab0",
X"0cff0b83",
X"caa034ff",
X"0b83caa1",
X"347751ff",
X"a5d83f83",
X"c0800883",
X"cad40c83",
X"c0800855",
X"83c08008",
X"80258838",
X"83c08008",
X"8f055574",
X"842c7083",
X"ffff0670",
X"882a5851",
X"557583ca",
X"a2347483",
X"caa33476",
X"83caa434",
X"ff800b83",
X"caa53481",
X"0b83caaf",
X"34a53974",
X"85962e09",
X"810680fe",
X"387583ca",
X"c80c7751",
X"ffa58c3f",
X"83caaf33",
X"83c08008",
X"07557483",
X"caaf3483",
X"caaf3381",
X"06557480",
X"2e833884",
X"5783caa4",
X"3383caa5",
X"3371882b",
X"07565c74",
X"81802e09",
X"8106a138",
X"83caa233",
X"83caa333",
X"71882b07",
X"565bad80",
X"75278738",
X"76820757",
X"9c397681",
X"07579639",
X"7482802e",
X"09810687",
X"38768307",
X"57873974",
X"81ff268a",
X"387783ca",
X"b81b0c76",
X"79348e3d",
X"0d04803d",
X"0d728429",
X"83cab805",
X"700883c0",
X"800c5182",
X"3d0d0480",
X"3d0d7270",
X"83c8900c",
X"70842981",
X"f6c00570",
X"0883cacc",
X"0c515182",
X"3d0d04fe",
X"3d0d8151",
X"de3f800b",
X"83ca9c0c",
X"800b83ca",
X"980cff0b",
X"83c8940c",
X"a80b83ca",
X"b40cae51",
X"caa33f80",
X"0b83cab8",
X"54528073",
X"70840555",
X"0c811252",
X"71842e09",
X"8106ef38",
X"843d0d04",
X"fe3d0d74",
X"02840596",
X"05225353",
X"71802e96",
X"38727081",
X"05543351",
X"caae3fff",
X"127083ff",
X"ff065152",
X"e739843d",
X"0d04fe3d",
X"0d029205",
X"225382ac",
X"51e4cf3f",
X"80c351ca",
X"8b3f8196",
X"51e4c33f",
X"725283c8",
X"9851ffb4",
X"3f725283",
X"c89851f8",
X"cd3f83c0",
X"800881ff",
X"0651c9e8",
X"3f843d0d",
X"04ffb13d",
X"0d80d13d",
X"f80551f8",
X"f73f83ca",
X"9c088105",
X"83ca9c0c",
X"80cf3d33",
X"cf117081",
X"ff065156",
X"56748326",
X"88e63875",
X"8f06ff05",
X"567583c8",
X"94082e9b",
X"38758326",
X"96387583",
X"c8940c75",
X"842983ca",
X"b8057008",
X"53557551",
X"f9fb3f80",
X"762488c2",
X"38758429",
X"83cab805",
X"55740880",
X"2e88b338",
X"83c89408",
X"842983ca",
X"b8057008",
X"02880582",
X"b9053352",
X"5b557480",
X"d22e84b0",
X"387480d2",
X"24903874",
X"bf2e9c38",
X"7480d02e",
X"81d53887",
X"f2397480",
X"d32e80d3",
X"387480d7",
X"2e81c438",
X"87e13902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"5656c8e4",
X"3f80c151",
X"c89e3ff6",
X"983f83ca",
X"cf3383c8",
X"98348152",
X"83c89851",
X"c9bb3f81",
X"51fde73f",
X"748b3883",
X"cacc0883",
X"cab40c87",
X"39a80b83",
X"cab40cc8",
X"af3f80c1",
X"51c7e93f",
X"f5e33f90",
X"0b83caaf",
X"33810656",
X"5674802e",
X"83389856",
X"83caa433",
X"83caa533",
X"71882b07",
X"56597481",
X"802e0981",
X"069c3883",
X"caa23383",
X"caa33371",
X"882b0756",
X"57ad8075",
X"278c3875",
X"81800756",
X"853975a0",
X"07567583",
X"c89834ff",
X"0b83c899",
X"34e00b83",
X"c89a3480",
X"0b83c89b",
X"34845283",
X"c89851c8",
X"b03f8451",
X"869b3902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"5659c7a4",
X"3f7951ff",
X"9fb93f83",
X"c0800880",
X"2e8a3880",
X"ce51c6d0",
X"3f85f139",
X"80c151c6",
X"c73fc7b8",
X"3fc5f13f",
X"83cac808",
X"58837525",
X"9b3883ca",
X"a43383ca",
X"a5337188",
X"2b07fc17",
X"71297a05",
X"8380055a",
X"51578d39",
X"74818029",
X"18ff8005",
X"58818057",
X"80567676",
X"2e9238c6",
X"a33f83c0",
X"800883c8",
X"98173481",
X"1656eb39",
X"c6923f83",
X"c0800881",
X"ff067753",
X"83c89852",
X"56f4bf3f",
X"83c08008",
X"81ff0655",
X"75752e09",
X"81068195",
X"389451e0",
X"8d3fc68c",
X"3f80c151",
X"c5c63fc6",
X"b73f7752",
X"7951ff9d",
X"cc3f805e",
X"80d13dfd",
X"f4055476",
X"5383c898",
X"527951ff",
X"9bd23f02",
X"82b90533",
X"55815974",
X"80d72e09",
X"810680c5",
X"38775279",
X"51ff9d9d",
X"3f80d13d",
X"fdf00554",
X"76538f3d",
X"70537a52",
X"58ff9cd5",
X"3f805676",
X"762ea238",
X"751883c8",
X"98173371",
X"33707232",
X"70307080",
X"2570307f",
X"06811d5d",
X"5f515151",
X"525b55db",
X"3982ac51",
X"df883f78",
X"802e8638",
X"80c35184",
X"3980ce51",
X"c4ba3fc5",
X"ab3fc3e4",
X"3f83d839",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"05595580",
X"705d5980",
X"e451ded2",
X"3fc4d13f",
X"80c151c4",
X"8b3f83ca",
X"b008792e",
X"82d63883",
X"cad40880",
X"fc055580",
X"fd527451",
X"85c13f83",
X"c080085b",
X"778224b2",
X"38ff1870",
X"872b83ff",
X"ff800681",
X"f58c0583",
X"c8985957",
X"55818055",
X"75708105",
X"57337770",
X"81055934",
X"ff157081",
X"ff065155",
X"74ea3882",
X"85397782",
X"e82e81a3",
X"387782e9",
X"2e098106",
X"81aa3878",
X"58778732",
X"70307072",
X"0780257a",
X"8a327030",
X"70720780",
X"25730753",
X"545a5157",
X"5575802e",
X"97387878",
X"269238a0",
X"0b83c898",
X"1a348119",
X"7081ff06",
X"5a55eb39",
X"81187081",
X"ff065955",
X"8a7827ff",
X"bc388f58",
X"83c89318",
X"3383c898",
X"1934ff18",
X"7081ff06",
X"59557784",
X"26ea3890",
X"58800b83",
X"c8981934",
X"81187081",
X"ff067098",
X"2b525955",
X"748025e9",
X"3880c655",
X"7a858f24",
X"843880c2",
X"557483c8",
X"983480f1",
X"0b83c89b",
X"34810b83",
X"c89c347a",
X"83c89934",
X"7a882c55",
X"7483c89a",
X"3480cb39",
X"82f07825",
X"80c43877",
X"80fd29fd",
X"97d30552",
X"7951ff99",
X"f83f80d1",
X"3dfdec05",
X"5480fd53",
X"83c89852",
X"7951ff99",
X"b03f7b81",
X"19595675",
X"80fc2483",
X"38785877",
X"882c5574",
X"83c99534",
X"7783c996",
X"347583c9",
X"97348180",
X"5980cc39",
X"83cac808",
X"57837825",
X"9b3883ca",
X"a43383ca",
X"a5337188",
X"2b07fc1a",
X"71297905",
X"83800559",
X"51598d39",
X"77818029",
X"17ff8005",
X"57818059",
X"76527951",
X"ff99863f",
X"80d13dfd",
X"ec055478",
X"5383c898",
X"527951ff",
X"98bf3f78",
X"51f6bf3f",
X"c1ce3fc0",
X"873f8b39",
X"83ca9808",
X"810583ca",
X"980c80d1",
X"3d0d04f6",
X"e03ffc39",
X"fc3d0d76",
X"78718429",
X"83cab805",
X"70085153",
X"5353709e",
X"3880ce72",
X"3480cf0b",
X"81133480",
X"ce0b8213",
X"3480c50b",
X"83133470",
X"84133480",
X"e73983ca",
X"d0133354",
X"80d27234",
X"73822a70",
X"81065151",
X"80cf5370",
X"843880d7",
X"53728113",
X"34a00b82",
X"13347383",
X"06517081",
X"2e9e3870",
X"81248838",
X"70802e8f",
X"389f3970",
X"822e9238",
X"70832e92",
X"38933980",
X"d8558e39",
X"80d35589",
X"3980cd55",
X"843980c4",
X"55748313",
X"3480c40b",
X"84133480",
X"0b851334",
X"863d0d04",
X"83c89008",
X"83c0800c",
X"04803d0d",
X"83c89008",
X"842981f6",
X"e0057008",
X"83c0800c",
X"51823d0d",
X"04fc3d0d",
X"76785354",
X"81538055",
X"87397110",
X"73105452",
X"73722651",
X"72802ea7",
X"3870802e",
X"86387180",
X"25e83872",
X"802e9838",
X"71742689",
X"38737231",
X"75740756",
X"5472812a",
X"72812a53",
X"53e53973",
X"51788338",
X"74517083",
X"c0800c86",
X"3d0d04fe",
X"3d0d8053",
X"75527451",
X"ffa33f84",
X"3d0d04fe",
X"3d0d8153",
X"75527451",
X"ff933f84",
X"3d0d04fb",
X"3d0d7779",
X"55558056",
X"74762586",
X"38743055",
X"81567380",
X"25883873",
X"30768132",
X"57548053",
X"73527451",
X"fee73f83",
X"c0800854",
X"75802e87",
X"3883c080",
X"08305473",
X"83c0800c",
X"873d0d04",
X"fa3d0d78",
X"7a575580",
X"57747725",
X"86387430",
X"55815775",
X"9f2c5481",
X"53757432",
X"74315274",
X"51feaa3f",
X"83c08008",
X"5476802e",
X"873883c0",
X"80083054",
X"7383c080",
X"0c883d0d",
X"04fc3d0d",
X"76558075",
X"0c800b84",
X"160c800b",
X"88160c80",
X"0b8c160c",
X"83c7f451",
X"80e9a93f",
X"87a68033",
X"7081ff06",
X"7071842a",
X"06515152",
X"d78b3f71",
X"812a8132",
X"72813271",
X"81067181",
X"06318418",
X"0c545471",
X"832a8132",
X"72822a81",
X"32708106",
X"72713178",
X"0c515353",
X"87a09033",
X"87a09133",
X"7081ff06",
X"70730681",
X"32810688",
X"190c5153",
X"5383c080",
X"08802e80",
X"c23883c0",
X"8008812a",
X"70810683",
X"c0800881",
X"06318417",
X"0c5283c0",
X"8008832a",
X"83c08008",
X"822a7181",
X"06718106",
X"31770c53",
X"5383c080",
X"08842a81",
X"0688160c",
X"83c08008",
X"852a8106",
X"8c160c86",
X"3d0d04fe",
X"3d0d7476",
X"54527151",
X"feb33f72",
X"812ea238",
X"8173268d",
X"3872822e",
X"a8387283",
X"2e9c38e6",
X"397108e2",
X"38841208",
X"dd388812",
X"08d838a5",
X"39881208",
X"812e9e38",
X"91398812",
X"08812e95",
X"38710891",
X"38841208",
X"8c388c12",
X"08812e09",
X"8106ffb2",
X"38843d0d",
X"04fb3d0d",
X"78028405",
X"9f053355",
X"56800b81",
X"ee885653",
X"81732b74",
X"06527180",
X"2e833881",
X"52747082",
X"05562270",
X"73902b07",
X"90809c0c",
X"51811353",
X"72882e09",
X"8106d938",
X"805383ca",
X"dc133351",
X"7081ff2e",
X"b2387010",
X"81eca805",
X"70225551",
X"80731770",
X"33701081",
X"eca80570",
X"22515151",
X"52527371",
X"2e913881",
X"12527186",
X"2e098106",
X"f1387390",
X"809c0c81",
X"13537286",
X"2e098106",
X"ffb83880",
X"53721670",
X"33515170",
X"81ff2e94",
X"38701081",
X"eca80570",
X"22708480",
X"80079080",
X"9c0c5151",
X"81135372",
X"862e0981",
X"06d73880",
X"53721651",
X"703383ca",
X"dc143481",
X"13537286",
X"2e098106",
X"ec38873d",
X"0d0404fe",
X"3d0d7502",
X"84059305",
X"33810652",
X"52708838",
X"71908094",
X"0c8e3970",
X"812e0981",
X"06863871",
X"9080980c",
X"843d0d04",
X"fb3d0d78",
X"982b7098",
X"2c7b982b",
X"70982c02",
X"90059f05",
X"33810683",
X"caf81170",
X"3370982b",
X"70982c51",
X"585c5a56",
X"51555154",
X"70742e09",
X"81069438",
X"83cad812",
X"3370982b",
X"70982c51",
X"52567073",
X"2eb13873",
X"75347283",
X"cad81334",
X"83cad933",
X"83caf933",
X"71982b71",
X"902b0783",
X"cad83370",
X"882b7207",
X"83caf833",
X"71079080",
X"b80c5259",
X"53545287",
X"3d0d04fe",
X"3d0d7481",
X"11337133",
X"71882b07",
X"83c0800c",
X"5351843d",
X"0d0483ca",
X"e43383c0",
X"800c04f5",
X"3d0d02bb",
X"05330284",
X"05bf0533",
X"02880580",
X"c3053302",
X"8c0580c6",
X"0522665c",
X"5a5e5c56",
X"7a557b54",
X"8953a152",
X"7d5180df",
X"843f83c0",
X"800881ff",
X"0683c080",
X"0c8d3d0d",
X"0483c08c",
X"080283c0",
X"8c0cf53d",
X"0d83c08c",
X"08880508",
X"83c08c08",
X"8f053383",
X"c08c0892",
X"0522028c",
X"05739005",
X"83c08c08",
X"e8050c83",
X"c08c08f8",
X"050c83c0",
X"8c08f005",
X"0c83c08c",
X"08ec050c",
X"83c08c08",
X"f4050c80",
X"0b83c08c",
X"08f00508",
X"83c08c08",
X"e0050c83",
X"c08c08fc",
X"050c83c0",
X"8c08f005",
X"0889278a",
X"38890b83",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08860587",
X"fffc0683",
X"c08c08e0",
X"050c0283",
X"c08c08e0",
X"0508310d",
X"853d7055",
X"83c08c08",
X"ec050854",
X"83c08c08",
X"f0050853",
X"83c08c08",
X"f4050852",
X"83c08c08",
X"e4050c80",
X"e8dd3f83",
X"c0800881",
X"ff0683c0",
X"8c08e405",
X"0883c08c",
X"08ec050c",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508802e",
X"8c3883c0",
X"8c08f805",
X"080d89c8",
X"3983c08c",
X"08f00508",
X"802e89a6",
X"3883c08c",
X"08ec0508",
X"81053383",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08842ea9",
X"38840b83",
X"c08c08e0",
X"05082588",
X"c73883c0",
X"8c08e005",
X"08852e85",
X"9b3883c0",
X"8c08e005",
X"08a12e87",
X"ad3888ac",
X"39800b83",
X"c08c08ec",
X"05088505",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"fc050c83",
X"c08c08e0",
X"0508832e",
X"09810688",
X"833883c0",
X"8c08e805",
X"08810533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"05088126",
X"87e63881",
X"0b83c08c",
X"08e00508",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08fc05",
X"0c83c08c",
X"08ec0508",
X"82053383",
X"c08c08e0",
X"05088705",
X"3483c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c800b83",
X"c08c08e0",
X"05088b05",
X"3483c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08f405",
X"0c800b83",
X"c08c08e0",
X"05088c05",
X"3483c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c800b83",
X"c08c08e0",
X"05088d05",
X"3483c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08f405",
X"0c800b83",
X"c08c08e0",
X"05088e05",
X"2383c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c800b83",
X"c08c08e0",
X"05088a05",
X"3483c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080570",
X"940508fc",
X"ffff0671",
X"94050c83",
X"c08c08e0",
X"050c83c0",
X"8c08ec05",
X"08860533",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c83c0",
X"8c08e005",
X"0883c08c",
X"08fc0508",
X"2e098106",
X"b63883c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c83c0",
X"8c08fc05",
X"0883c08c",
X"08e00508",
X"8b053483",
X"c08c08ec",
X"05088705",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e0050881",
X"2e8f3883",
X"c08c08e0",
X"0508822e",
X"b738848c",
X"3983c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08f405",
X"0c820b83",
X"c08c08e0",
X"05088a05",
X"3483d939",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"83c08c08",
X"fc050883",
X"c08c08e0",
X"05088a05",
X"3483a139",
X"83c08c08",
X"fc050880",
X"2e839538",
X"83c08c08",
X"ec050883",
X"05338306",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508832e",
X"09810682",
X"f33883c0",
X"8c08ec05",
X"08820533",
X"70982b83",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08e00508",
X"802582cc",
X"3883c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08f405",
X"0c83c08c",
X"08ec0508",
X"86053383",
X"c08c08e0",
X"050880d6",
X"053483c0",
X"8c08e005",
X"08840583",
X"c08c08ec",
X"05088205",
X"338f0683",
X"c08c08e4",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08e40508",
X"83c08c08",
X"e0050834",
X"83c08c08",
X"ec050884",
X"053383c0",
X"8c08e005",
X"08810534",
X"800b83c0",
X"8c08e005",
X"08820534",
X"83c08c08",
X"e0050808",
X"ff83ff06",
X"82800783",
X"c08c08e0",
X"05080c83",
X"c08c08e8",
X"05088105",
X"33810583",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"0883c08c",
X"08e80508",
X"81053481",
X"833983c0",
X"8c08fc05",
X"08802e80",
X"f73883c0",
X"8c08ec05",
X"08860533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508a22e",
X"09810680",
X"d73883c0",
X"8c08ec05",
X"08880533",
X"83c08c08",
X"ec050887",
X"05337182",
X"80290583",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"5283c08c",
X"08e4050c",
X"83c08c08",
X"f4050c83",
X"c08c08e4",
X"050883c0",
X"8c08e005",
X"08880523",
X"83c08c08",
X"ec050833",
X"83c08c08",
X"f0050871",
X"317083ff",
X"ff0683c0",
X"8c08f005",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"ec050805",
X"83c08c08",
X"ec050cf6",
X"d03983c0",
X"8c08f805",
X"080d83c0",
X"8c08f005",
X"0883c08c",
X"08e0050c",
X"83c08c08",
X"f805080d",
X"83c08c08",
X"e0050883",
X"c0800c8d",
X"3d0d83c0",
X"8c0c0483",
X"c08c0802",
X"83c08c0c",
X"e73d0d83",
X"c08c0888",
X"05080284",
X"0583c08c",
X"08e8050c",
X"83c08c08",
X"d4050c80",
X"0b83cb80",
X"3483c08c",
X"08d40508",
X"900583c0",
X"8c08c405",
X"0c800b83",
X"c08c08c4",
X"05083480",
X"0b83c08c",
X"08c40508",
X"81053480",
X"0b83c08c",
X"08c8050c",
X"83c08c08",
X"c8050880",
X"d82983c0",
X"8c08c405",
X"080583c0",
X"8c08ffb8",
X"050c800b",
X"83c08c08",
X"ffb80508",
X"80d8050c",
X"83c08c08",
X"ffb80508",
X"840583c0",
X"8c08ffb8",
X"050c83c0",
X"8c08c805",
X"0883c08c",
X"08ffb805",
X"0834880b",
X"83c08c08",
X"ffb80508",
X"81053480",
X"0b83c08c",
X"08ffb805",
X"08820534",
X"83c08c08",
X"ffb80508",
X"08ffa1ff",
X"06a08007",
X"83c08c08",
X"ffb80508",
X"0c83c08c",
X"08c80508",
X"81057081",
X"ff0683c0",
X"8c08c805",
X"0c83c08c",
X"08ffb805",
X"0c810b83",
X"c08c08c8",
X"050827fe",
X"db3883c0",
X"8c08ec05",
X"705483c0",
X"8c08cc05",
X"0c925283",
X"c08c08d4",
X"05085180",
X"dc843f83",
X"c0800881",
X"ff067083",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"bc050891",
X"c63883c0",
X"8c08f405",
X"51f18c3f",
X"83c08008",
X"83ffff06",
X"83c08c08",
X"f6055283",
X"c08c08e0",
X"050cf0f3",
X"3f83c080",
X"0883ffff",
X"0683c08c",
X"08fd0533",
X"83c08c08",
X"ffbc0508",
X"83c08c08",
X"c8050c83",
X"c08c08c0",
X"050c83c0",
X"8c08dc05",
X"0c83c08c",
X"08c80508",
X"83c08c08",
X"c0050827",
X"80fe3883",
X"c08c08cc",
X"05085483",
X"c08c08c8",
X"05085389",
X"5283c08c",
X"08d40508",
X"5180db8b",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffbc0508",
X"83eb3883",
X"c08c08ee",
X"0551eff3",
X"3f83c080",
X"0883ffff",
X"065383c0",
X"8c08c805",
X"085283c0",
X"8c08d405",
X"0851f0b5",
X"3f83c08c",
X"08c80508",
X"81057081",
X"ff0683c0",
X"8c08c805",
X"0c83c08c",
X"08ffb805",
X"0cfef239",
X"83c08c08",
X"c4050881",
X"053383c0",
X"8c08c005",
X"0c83c08c",
X"08c00508",
X"839e3883",
X"c08c08c0",
X"050883c0",
X"8c08ffb8",
X"050c83c0",
X"8c08e005",
X"0888de2e",
X"0981068b",
X"38810b83",
X"c08c08ff",
X"b8050c83",
X"c08c08dc",
X"0508858e",
X"2e098106",
X"82c53881",
X"7083c08c",
X"08ffb805",
X"080683c0",
X"8c08ffb8",
X"050c83c0",
X"8c08c805",
X"0c83c08c",
X"08ffb805",
X"08802e82",
X"9e3883c0",
X"8c08c805",
X"0883c08c",
X"08c40508",
X"81053483",
X"c08c08c0",
X"050883c0",
X"8c08c405",
X"08870534",
X"83c08c08",
X"c0050883",
X"c08c08c4",
X"05088b05",
X"3483c08c",
X"08c00508",
X"83c08c08",
X"c405088c",
X"0534830b",
X"83c08c08",
X"c405088d",
X"053483c0",
X"8c08c005",
X"0883c08c",
X"08c40508",
X"8e052383",
X"0b83c08c",
X"08c40508",
X"8a053483",
X"c08c08c4",
X"05089405",
X"08838080",
X"0783c08c",
X"08c40508",
X"94050c83",
X"cae43370",
X"83c08c08",
X"c8050805",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb80508",
X"83cae434",
X"83c08c08",
X"ffbc0508",
X"83c08c08",
X"c4050894",
X"053483c0",
X"8c08c805",
X"0883c08c",
X"08c40508",
X"80d60534",
X"83c08c08",
X"c8050883",
X"c08c08c4",
X"05088405",
X"348e0b83",
X"c08c08c4",
X"05088505",
X"3483c08c",
X"08c00508",
X"83c08c08",
X"c4050886",
X"053483c0",
X"8c08c405",
X"08840508",
X"ff83ff06",
X"82800783",
X"c08c08c4",
X"05088405",
X"0ca23981",
X"db0b83c0",
X"8c08ffb8",
X"050c8cc3",
X"3983c08c",
X"08ffbc05",
X"0883c08c",
X"08ffb805",
X"0c8cb039",
X"83c08c08",
X"f1053352",
X"83c08c08",
X"d4050851",
X"80d7903f",
X"800b83c0",
X"8c08c405",
X"08810533",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"c8050c83",
X"c08c08c8",
X"050883c0",
X"8c08ffb8",
X"0508278a",
X"cb3883c0",
X"8c08c805",
X"0880d829",
X"7083c08c",
X"08c40508",
X"05708805",
X"70830533",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"cc050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08d8",
X"050c83c0",
X"8c08ffb8",
X"05088889",
X"3883c08c",
X"08ffbc05",
X"088d0533",
X"83c08c08",
X"d0050c83",
X"c08c08d0",
X"050887ed",
X"3883c08c",
X"08cc0508",
X"22028405",
X"71860587",
X"fffc0683",
X"c08c08ff",
X"b8050c83",
X"c08c08e4",
X"050c83c0",
X"8c08c005",
X"0c0283c0",
X"8c08ffb8",
X"0508310d",
X"893d7059",
X"83c08c08",
X"c0050858",
X"83c08c08",
X"ffbc0508",
X"87053357",
X"83c08c08",
X"ffb8050c",
X"a25583c0",
X"8c08d005",
X"08548653",
X"81815283",
X"c08c08d4",
X"05085180",
X"c9c33f83",
X"c0800881",
X"ff0683c0",
X"8c08d005",
X"0c83c08c",
X"08d00508",
X"81c03883",
X"c08c08ff",
X"bc050896",
X"055383c0",
X"8c08c005",
X"085283c0",
X"8c08ffb8",
X"050851ac",
X"f73f83c0",
X"800881ff",
X"0683c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"08802e81",
X"853883c0",
X"8c08ffbc",
X"05089405",
X"83c08c08",
X"ffbc0508",
X"96053370",
X"862a83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08c005",
X"0c83c08c",
X"08ffb805",
X"08832e09",
X"810680c6",
X"3883c08c",
X"08ffb805",
X"0883c08c",
X"08cc0508",
X"82053483",
X"cae43370",
X"810583c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb8",
X"050883ca",
X"e43483c0",
X"8c08ffbc",
X"050883c0",
X"8c08c005",
X"083483c0",
X"8c08e405",
X"080d83c0",
X"8c08d005",
X"0881ff06",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffbc0508",
X"fbe33883",
X"c08c08d8",
X"050883c0",
X"8c08c405",
X"08058805",
X"70820533",
X"5183c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"08832e09",
X"810680e3",
X"3883c08c",
X"08ffbc05",
X"0883c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"08810570",
X"81ff0651",
X"83c08c08",
X"ffb8050c",
X"810b83c0",
X"8c08ffb8",
X"050827dd",
X"38800b83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b8050881",
X"057081ff",
X"065183c0",
X"8c08ffb8",
X"050c970b",
X"83c08c08",
X"ffb80508",
X"27dd3883",
X"c08c08e0",
X"050880f9",
X"32703070",
X"80255151",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"dc050891",
X"2e098106",
X"80f93883",
X"c08c08ff",
X"b8050880",
X"2e80ec38",
X"83c08c08",
X"c8050880",
X"e238850b",
X"83c08c08",
X"c40508a6",
X"0534a00b",
X"83c08c08",
X"c40508a7",
X"0534850b",
X"83c08c08",
X"c40508a8",
X"053480c0",
X"0b83c08c",
X"08c40508",
X"a9053486",
X"0b83c08c",
X"08c40508",
X"aa053490",
X"0b83c08c",
X"08c40508",
X"ab053486",
X"0b83c08c",
X"08c40508",
X"ac0534a0",
X"0b83c08c",
X"08c40508",
X"ad053483",
X"c08c08e0",
X"050889d8",
X"32703070",
X"80255151",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"dc050883",
X"edec2e09",
X"810680f6",
X"38817083",
X"c08c08ff",
X"b8050806",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb80508",
X"802e80ce",
X"3883c08c",
X"08c80508",
X"80c43884",
X"0b83c08c",
X"08c40508",
X"aa053480",
X"c00b83c0",
X"8c08c405",
X"08ab0534",
X"840b83c0",
X"8c08c405",
X"08ac0534",
X"900b83c0",
X"8c08c405",
X"08ad0534",
X"83c08c08",
X"ffbc0508",
X"83c08c08",
X"c405088c",
X"053483c0",
X"8c08e005",
X"0880f932",
X"70307080",
X"25515183",
X"c08c08ff",
X"b8050c83",
X"c08c08dc",
X"0508862e",
X"09810680",
X"c3388170",
X"83c08c08",
X"ffb80508",
X"0683c08c",
X"08ffb805",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffb805",
X"08802e9c",
X"3883c08c",
X"08c80508",
X"933883c0",
X"8c08ffbc",
X"050883c0",
X"8c08c405",
X"088d0534",
X"83c08c08",
X"e00508b4",
X"b4327030",
X"70802551",
X"5183c08c",
X"08ffb805",
X"0c83c08c",
X"08dc0508",
X"90892e09",
X"8106a238",
X"83c08c08",
X"ffb80508",
X"802e9638",
X"83c08c08",
X"c805088d",
X"38820b83",
X"c08c08c4",
X"05088d05",
X"3483c08c",
X"08c80508",
X"80d82983",
X"c08c08c4",
X"05080570",
X"84057083",
X"053383c0",
X"8c08ffb8",
X"050c83c0",
X"8c08cc05",
X"0c83c08c",
X"08c0050c",
X"80588057",
X"83c08c08",
X"ffb80508",
X"56805580",
X"548a53a1",
X"5283c08c",
X"08d40508",
X"5180c1f5",
X"3f83c080",
X"0881ff06",
X"7030709f",
X"2a5183c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffbc",
X"0508a02e",
X"8c3883c0",
X"8c08ffb8",
X"0508f5dd",
X"3883c08c",
X"08c00508",
X"8b053383",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b8050880",
X"2eb43883",
X"c08c08cc",
X"05088305",
X"3383c08c",
X"08ffb805",
X"0c805880",
X"5783c08c",
X"08ffb805",
X"08568055",
X"80548b53",
X"a15283c0",
X"8c08d405",
X"085180c0",
X"f03f83c0",
X"8c08c805",
X"08810570",
X"81ff0683",
X"c08c08c4",
X"05088105",
X"335283c0",
X"8c08c805",
X"0c83c08c",
X"08ffb805",
X"0cf5a439",
X"800b83c0",
X"8c08c805",
X"0c83c08c",
X"08c80508",
X"80d82983",
X"c08c08d4",
X"05080570",
X"9a053383",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"b8050882",
X"2e098106",
X"a93883cb",
X"80568155",
X"805483c0",
X"8c08ffb8",
X"05085383",
X"c08c08ff",
X"bc050897",
X"05335283",
X"c08c08d4",
X"050851e0",
X"ae3f83c0",
X"8c08c805",
X"08810570",
X"81ff0683",
X"c08c08c8",
X"050c83c0",
X"8c08ffb8",
X"050c810b",
X"83c08c08",
X"c8050827",
X"fefb3881",
X"0b83c08c",
X"08c40508",
X"34800b83",
X"c08c08ff",
X"b8050c83",
X"c08c08e8",
X"05080d83",
X"c08c08ff",
X"b8050883",
X"c0800c9b",
X"3d0d83c0",
X"8c0c04f4",
X"3d0d901f",
X"59800b81",
X"1a33555b",
X"7a742781",
X"ad387a80",
X"d829198a",
X"11335555",
X"73832e09",
X"81068188",
X"38941533",
X"57805276",
X"51dde03f",
X"80538052",
X"7651de80",
X"3fb3e43f",
X"83c08008",
X"5c805877",
X"81c4291c",
X"87113355",
X"5573802e",
X"80c03874",
X"0881ec9c",
X"2e098106",
X"b5388075",
X"5b567580",
X"d8291a9a",
X"11335555",
X"73832e09",
X"81069238",
X"a4157033",
X"55557674",
X"278738ff",
X"14547375",
X"34811670",
X"81ff0657",
X"54817627",
X"d1388118",
X"7081ff06",
X"59548f78",
X"27ffa438",
X"83cae433",
X"ff055473",
X"83cae434",
X"811b7081",
X"ff06811b",
X"335f5c54",
X"7c7b26fe",
X"d538800b",
X"83c0800c",
X"8e3d0d04",
X"83c08c08",
X"0283c08c",
X"0ce63d0d",
X"83c08c08",
X"88050802",
X"84057190",
X"05703370",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"cc050c83",
X"c08c08dc",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08ffa405",
X"08802e9f",
X"8c38800b",
X"83c08c08",
X"cc050881",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08d405",
X"0c83c08c",
X"08d40508",
X"83c08c08",
X"ffa40508",
X"259ed438",
X"83c08c08",
X"d4050880",
X"d82983c0",
X"8c08cc05",
X"08058405",
X"70860533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffa40508",
X"802e9de0",
X"38b18a3f",
X"83c08c08",
X"ffbc0508",
X"80d40508",
X"83c08008",
X"269dc938",
X"0283c08c",
X"08ffbc05",
X"08810533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"d8050c83",
X"c08c08ff",
X"a4050883",
X"c08c08fc",
X"052383c0",
X"8c08ffa4",
X"05088605",
X"83fc0683",
X"c08c08ff",
X"a4050c02",
X"83c08c08",
X"ffa40508",
X"310d853d",
X"705583c0",
X"8c08fc05",
X"5483c08c",
X"08ffbc05",
X"085383c0",
X"8c08e005",
X"085283c0",
X"8c08c005",
X"0cb8e23f",
X"83c08008",
X"81ff0683",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a405089c",
X"923883c0",
X"8c08ffbc",
X"05088705",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e80",
X"d53883c0",
X"8c08ffbc",
X"05088605",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08822e09",
X"8106b338",
X"83c08c08",
X"fc052283",
X"c08c08ff",
X"a4050c87",
X"0b83c08c",
X"08ffa405",
X"08279738",
X"83c08c08",
X"c0050882",
X"055283c0",
X"8c08c005",
X"083351d7",
X"b43f83c0",
X"8c08ffbc",
X"05088605",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08832e09",
X"81069afb",
X"3883c08c",
X"08ffbc05",
X"08920583",
X"c08c08ff",
X"bc050889",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08c405",
X"0c83c08c",
X"08ffa405",
X"08832eb6",
X"3883c08c",
X"08c40508",
X"82053383",
X"c08c08fc",
X"052283c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa8",
X"050883c0",
X"8c08ffac",
X"0508269a",
X"9638800b",
X"83c08c08",
X"e4050c80",
X"0b83c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa405",
X"08832e09",
X"810688c1",
X"3883c08c",
X"08c00508",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffb005",
X"082e0981",
X"0687fa38",
X"83c08c08",
X"c0050881",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508942e",
X"09810687",
X"d83883c0",
X"8c08c005",
X"08820533",
X"70810683",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"b005082e",
X"8a38880b",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"a8050881",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e91",
X"3883c08c",
X"08e40508",
X"840783c0",
X"8c08e405",
X"0c83c08c",
X"08ffa805",
X"08822a70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e913883",
X"c08c08e4",
X"05088207",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"a8050883",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e91",
X"3883c08c",
X"08e40508",
X"810783c0",
X"8c08e405",
X"0c83c08c",
X"08c00508",
X"83053370",
X"982b83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"05088025",
X"913883c0",
X"8c08e405",
X"08900783",
X"c08c08e4",
X"050c83c0",
X"8c08ffa8",
X"050881ff",
X"0670852a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa40508",
X"802e9138",
X"83c08c08",
X"e40508a0",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"ffa80508",
X"842a7081",
X"065183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"923883c0",
X"8c08e405",
X"0880c007",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"a8050886",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e92",
X"3883c08c",
X"08e40508",
X"81800783",
X"c08c08e4",
X"050c83c0",
X"8c08ffa8",
X"05088106",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9238",
X"83c08c08",
X"e4050882",
X"800783c0",
X"8c08e405",
X"0c83c08c",
X"08ffa805",
X"08812a70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e923883",
X"c08c08e4",
X"05088480",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"c0050884",
X"05337098",
X"2b83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa405",
X"08802592",
X"3883c08c",
X"08e40508",
X"88800783",
X"c08c08e4",
X"050c83c0",
X"8c08c005",
X"08850533",
X"70982b83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050880",
X"25923883",
X"c08c08e4",
X"05089080",
X"0783c08c",
X"08e4050c",
X"83c08c08",
X"c0050882",
X"05337081",
X"ff067085",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa405",
X"08802e92",
X"3883c08c",
X"08e40508",
X"a0800783",
X"c08c08e4",
X"050c83c0",
X"8c08ffa8",
X"0508842a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9338",
X"83c08c08",
X"e4050880",
X"c0800783",
X"c08c08e4",
X"050c83c0",
X"8c08ffa8",
X"0508862a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9338",
X"83c08c08",
X"e4050881",
X"80800783",
X"c08c08e4",
X"050c83c0",
X"8c08ffac",
X"0508982b",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"80259338",
X"83c08c08",
X"e4050882",
X"80800783",
X"c08c08e4",
X"050c83c0",
X"8c08c005",
X"08870533",
X"70982b83",
X"c08c08c0",
X"05088905",
X"3370982b",
X"70982c73",
X"982c8180",
X"05545153",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa80508",
X"83c08c08",
X"f8052380",
X"ff0b83c0",
X"8c08ffa4",
X"05083183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08fa",
X"052384d9",
X"39800b83",
X"c08c08e4",
X"050c8180",
X"0b83c08c",
X"08f80523",
X"81800b83",
X"c08c08fa",
X"052384b9",
X"3983c08c",
X"08ffb005",
X"081083c0",
X"8c0805f8",
X"0583c08c",
X"08ffb005",
X"08842983",
X"c08c08ff",
X"b0050810",
X"0583c08c",
X"08c40508",
X"05708405",
X"703383c0",
X"8c08c005",
X"08057033",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffb80508",
X"2383c08c",
X"08ffa805",
X"08810533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"902e0981",
X"06be3883",
X"c08c08ff",
X"a8050833",
X"83c08c08",
X"c0050805",
X"81057033",
X"70828029",
X"83c08c08",
X"ffb40508",
X"05515183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"b8050823",
X"83c08c08",
X"ffac0508",
X"86052283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a80508a2",
X"3883c08c",
X"08ffac05",
X"08880522",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"81ff2e80",
X"e53883c0",
X"8c08ffb8",
X"05082270",
X"83c08c08",
X"ffa80508",
X"31708280",
X"29713183",
X"c08c08ff",
X"ac050888",
X"05227083",
X"c08c08ff",
X"a8050831",
X"70733553",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffb805",
X"082383c0",
X"8c08ffb0",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa4050c",
X"810b83c0",
X"8c08ffb0",
X"050827fc",
X"e038800b",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffb00508",
X"1083c08c",
X"08c40508",
X"05709005",
X"703383c0",
X"8c08c005",
X"08057033",
X"72810533",
X"70720651",
X"535183c0",
X"8c08ffa8",
X"050c5183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e9b3890",
X"0b83c08c",
X"08ffb005",
X"082b83c0",
X"8c08e405",
X"080783c0",
X"8c08e405",
X"0c83c08c",
X"08ffb005",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a4050c97",
X"0b83c08c",
X"08ffb005",
X"0827fef4",
X"3883c08c",
X"08f80522",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"bf269138",
X"83c08c08",
X"e4050882",
X"0783c08c",
X"08e4050c",
X"81c00b83",
X"c08c08ff",
X"a4050827",
X"913883c0",
X"8c08e405",
X"08810783",
X"c08c08e4",
X"050c83c0",
X"8c08fa05",
X"2283c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08bf2691",
X"3883c08c",
X"08e40508",
X"880783c0",
X"8c08e405",
X"0c81c00b",
X"83c08c08",
X"ffa40508",
X"27913883",
X"c08c08e4",
X"05088407",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"bc050890",
X"053383c0",
X"8c08e405",
X"0883c08c",
X"08ffa405",
X"0c83c08c",
X"08c4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffbc0508",
X"8c05082e",
X"85e03883",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"bc05088c",
X"050c83c0",
X"8c08ffbc",
X"05088905",
X"3383c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa805",
X"08802e85",
X"9a3883c0",
X"8c08e405",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffa40508",
X"8f0683c0",
X"8c08e405",
X"0c83c08c",
X"08ffb005",
X"0c83c08c",
X"08d0050c",
X"83c08c08",
X"ffa80508",
X"822e0981",
X"0681c238",
X"800b83c0",
X"8c08ffa4",
X"0508862a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffa80508",
X"2e8c3881",
X"c00b83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffb0",
X"0508872a",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9438",
X"83c08c08",
X"ffa80508",
X"81903283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"b0050884",
X"2a708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e94",
X"3883c08c",
X"08ffa805",
X"0880d032",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffb00508",
X"83c08c08",
X"ffa80508",
X"3283c08c",
X"08ffb005",
X"0c800b83",
X"c08c08f0",
X"050c800b",
X"83c08c08",
X"f4052380",
X"0b81ee98",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffb805",
X"082e82d3",
X"3883c08c",
X"08f00581",
X"ee980b83",
X"c08c08ff",
X"ac050c83",
X"c08c08c8",
X"050c83c0",
X"8c08ffac",
X"05083383",
X"c08c08ff",
X"ac050881",
X"05338172",
X"2b81722b",
X"077083c0",
X"8c08ffb0",
X"05080652",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffa80508",
X"2e098106",
X"81be3883",
X"c08c08ff",
X"b8050885",
X"2680f638",
X"83c08c08",
X"ffac0508",
X"82053370",
X"81ff0683",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050880",
X"2e80ca38",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"ffb80508",
X"81057081",
X"ff0683c0",
X"8c08c805",
X"08730553",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffa40508",
X"3483c08c",
X"08ffac05",
X"08830533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e9d38",
X"810b83c0",
X"8c08ffa4",
X"05082b83",
X"c08c08d0",
X"05080807",
X"83c08c08",
X"d005080c",
X"83c08c08",
X"ffac0508",
X"84057033",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa40508",
X"fdc83883",
X"c08c08f0",
X"05528051",
X"c1fb3f83",
X"c08c08e4",
X"05085283",
X"c08c08c4",
X"050851c3",
X"b63f83c0",
X"8c08fb05",
X"33708180",
X"0a29810a",
X"0570982c",
X"5583c08c",
X"08ffa405",
X"0c83c08c",
X"08f90533",
X"7081800a",
X"29810a05",
X"70982c55",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"c4050853",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa8050c",
X"c38e3f83",
X"c08c08ff",
X"bc050888",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"84e13883",
X"c08c08ff",
X"bc050890",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"05088126",
X"84c13880",
X"7081eed8",
X"0b81eed8",
X"0b810533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffb40508",
X"2e81ae38",
X"83c08c08",
X"ffac0508",
X"842983c0",
X"8c08ffa8",
X"05080570",
X"3383c08c",
X"08c00508",
X"05703372",
X"81053370",
X"72065153",
X"5183c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802eaa",
X"38810b83",
X"c08c08ff",
X"ac05082b",
X"83c08c08",
X"ffb40508",
X"077083ff",
X"ff0683c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffac",
X"05088105",
X"7081ff06",
X"81eed871",
X"84297105",
X"70810533",
X"515383c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508fed4",
X"3883c08c",
X"08ffbc05",
X"088a0522",
X"83c08c08",
X"c0050c83",
X"c08c08ff",
X"b4050883",
X"c08c08c0",
X"05082e82",
X"ae38800b",
X"83c08c08",
X"e8050c80",
X"0b83c08c",
X"08ec0523",
X"807083c0",
X"8c08e805",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffb0050c",
X"81af3983",
X"c08c08ff",
X"b4050883",
X"c08c08ff",
X"ac05082c",
X"70810651",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e80e7",
X"3883c08c",
X"08ffb005",
X"0883c08c",
X"08ffb005",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"b8050873",
X"0583c08c",
X"08ffbc05",
X"08900533",
X"83c08c08",
X"ffac0508",
X"84290553",
X"5383c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa805",
X"0881eeda",
X"053383c0",
X"8c08ffa4",
X"05083483",
X"c08c08ff",
X"ac050881",
X"057081ff",
X"0683c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa405",
X"0c8f0b83",
X"c08c08ff",
X"ac050827",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb00508",
X"85268c38",
X"83c08c08",
X"ffa40508",
X"fea93883",
X"c08c08e8",
X"05528051",
X"ffbcaa3f",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffbc0508",
X"8a052383",
X"c08c08ff",
X"bc050880",
X"d2053383",
X"c08c08ff",
X"bc050880",
X"d4050805",
X"83c08c08",
X"ffbc0508",
X"80d4050c",
X"83c08c08",
X"d805080d",
X"83c08c08",
X"d4050881",
X"800a2981",
X"800a0570",
X"982c83c0",
X"8c08cc05",
X"08810533",
X"83c08c08",
X"ffa8050c",
X"5183c08c",
X"08d4050c",
X"83c08c08",
X"ffa80508",
X"83c08c08",
X"d4050824",
X"e1ae3880",
X"0b83c08c",
X"08ffa805",
X"0c83c08c",
X"08dc0508",
X"0d83c08c",
X"08ffa805",
X"0883c080",
X"0c9c3d0d",
X"83c08c0c",
X"04f33d0d",
X"02bf0533",
X"02840580",
X"c3053383",
X"cb80335a",
X"5b597980",
X"2e8d3878",
X"78065776",
X"802e8e38",
X"818a3978",
X"78065776",
X"802e8180",
X"3883cb80",
X"33707a07",
X"58587988",
X"38780970",
X"79065157",
X"7683cb80",
X"3492983f",
X"83c08008",
X"5e805c8f",
X"5d7d1c87",
X"11335858",
X"76802e80",
X"c2387708",
X"81ec9c2e",
X"098106b7",
X"38805b81",
X"5a7d1c70",
X"1c9a1133",
X"59595976",
X"822e0981",
X"06953883",
X"cb805681",
X"55805476",
X"53971833",
X"527851ff",
X"bd813fff",
X"1a80d81c",
X"5c5a7980",
X"25cf38ff",
X"1d81c41d",
X"5d5d7c80",
X"25ffa638",
X"8f3d0d04",
X"e93d0d69",
X"6c028805",
X"80ea0522",
X"5c5a5b80",
X"7071415e",
X"58ff7879",
X"7a7b7c7d",
X"464c4a45",
X"405d4362",
X"993d3462",
X"02840580",
X"dd053477",
X"792280ff",
X"ff065445",
X"72792379",
X"782e8887",
X"387a7081",
X"055c3370",
X"842a718c",
X"0670822a",
X"5a565683",
X"06ff1b70",
X"83ffff06",
X"5c545680",
X"5475742e",
X"91387a70",
X"81055c33",
X"ff1b7083",
X"ffff065c",
X"54548176",
X"279b3873",
X"81ff067b",
X"7081055d",
X"33557482",
X"802905ff",
X"1b7083ff",
X"ff065c54",
X"54827627",
X"aa387383",
X"ffff067b",
X"7081055d",
X"3370902b",
X"72077d70",
X"81055f33",
X"70982b72",
X"07fe1f70",
X"83ffff06",
X"40525252",
X"5254547e",
X"802e80c4",
X"387686f7",
X"38748a2e",
X"09810694",
X"38811f70",
X"81ff0681",
X"1e7081ff",
X"065f5240",
X"5386dc39",
X"748c2e09",
X"810686d3",
X"38ff1f70",
X"81ff06ff",
X"1e7081ff",
X"065f5240",
X"537b6325",
X"86bd38ff",
X"4386b839",
X"76812e83",
X"bb387681",
X"24893876",
X"802e8d38",
X"86a53976",
X"822e84a6",
X"38869c39",
X"f8155372",
X"84268495",
X"38728429",
X"81ef9805",
X"53720804",
X"64802e80",
X"cd387822",
X"83808006",
X"53728380",
X"802e0981",
X"06bc3880",
X"56756427",
X"a438751e",
X"7083ffff",
X"0677101b",
X"90117283",
X"2a585157",
X"51537375",
X"34728706",
X"81712b51",
X"53728116",
X"34811670",
X"81ff0657",
X"53977627",
X"cc387f84",
X"0740800b",
X"993d4356",
X"61167033",
X"70982b70",
X"982c5151",
X"51538073",
X"2480fb38",
X"6073291e",
X"7083ffff",
X"067a2283",
X"80800652",
X"58537283",
X"80802e09",
X"810680de",
X"38608832",
X"70307072",
X"07802563",
X"90327030",
X"70720780",
X"25730753",
X"54585155",
X"5373802e",
X"bd387687",
X"065372b6",
X"38758429",
X"76100579",
X"11841179",
X"832a5757",
X"51537375",
X"34608116",
X"34658614",
X"23668814",
X"23758738",
X"7f810740",
X"8d397581",
X"2e098106",
X"85387f82",
X"07408116",
X"7081ff06",
X"57538176",
X"27fee538",
X"6361291e",
X"7083ffff",
X"065f5380",
X"704642ff",
X"02840580",
X"dd0534ff",
X"0b993d34",
X"83f53981",
X"1c7081ff",
X"065d5380",
X"4273812e",
X"0981068e",
X"38778180",
X"0a298180",
X"0a055880",
X"d3397380",
X"2e893873",
X"822e0981",
X"068d387c",
X"81800a29",
X"81800a05",
X"5da43981",
X"5f83b839",
X"ff1c7081",
X"ff065d53",
X"7b632583",
X"38ff437c",
X"802e9238",
X"7c81800a",
X"2981ff0a",
X"055d7c98",
X"2c5d8393",
X"3977802e",
X"92387781",
X"800a2981",
X"ff0a0558",
X"77982c58",
X"82fd3977",
X"53839e39",
X"74892680",
X"f4387484",
X"2981efac",
X"05537208",
X"0473872e",
X"82e13873",
X"852e82db",
X"3873882e",
X"82d53873",
X"8c2e82cf",
X"3873892e",
X"09810686",
X"38814582",
X"c2397381",
X"2e098106",
X"82b93862",
X"802582b3",
X"387b982b",
X"70982c51",
X"4382a839",
X"7383ffff",
X"0646829f",
X"397383ff",
X"ff064782",
X"96397381",
X"ff064182",
X"8e397381",
X"1a348287",
X"397381ff",
X"064481ff",
X"397e5382",
X"a0397481",
X"2e81e338",
X"74812489",
X"3874802e",
X"8d3881e7",
X"3974822e",
X"81d83881",
X"de397456",
X"7b833881",
X"56745373",
X"862e0981",
X"06973875",
X"81065372",
X"802e8e38",
X"782282ff",
X"ff06fe80",
X"800753b6",
X"397b8338",
X"81537382",
X"2e098106",
X"97387281",
X"06537280",
X"2e8e3878",
X"2281ffff",
X"06818080",
X"07539339",
X"7b9638fc",
X"14537281",
X"268e3878",
X"22ff8080",
X"07537279",
X"2380e539",
X"80557381",
X"2e098106",
X"83387355",
X"77537780",
X"2e893874",
X"81065372",
X"80ca3872",
X"d0155455",
X"72812683",
X"38815577",
X"802eb938",
X"74810653",
X"72802eb0",
X"38782283",
X"80800653",
X"72838080",
X"2e098106",
X"9f3873b0",
X"2e098106",
X"87386199",
X"3d349139",
X"73b12e09",
X"81068938",
X"61028405",
X"80dd0534",
X"61810553",
X"8c396174",
X"31810553",
X"84396114",
X"537283ff",
X"ff064279",
X"f7fb387d",
X"832a5372",
X"821a3478",
X"22838080",
X"06537283",
X"80802e09",
X"81068838",
X"81537f87",
X"2e833880",
X"537283c0",
X"800c993d",
X"0d04fd3d",
X"0d758311",
X"33821233",
X"71982b71",
X"902b0781",
X"14337088",
X"2b720775",
X"33710783",
X"c0800c52",
X"53545654",
X"52853d0d",
X"04f63d0d",
X"02b70533",
X"028405bb",
X"05330288",
X"05bf0533",
X"5b5b5b80",
X"58805778",
X"882b7a07",
X"5680557a",
X"548153a3",
X"527c5192",
X"cc3f83c0",
X"800881ff",
X"0683c080",
X"0c8c3d0d",
X"04f63d0d",
X"02b70533",
X"028405bb",
X"05330288",
X"05bf0533",
X"5b5b5b80",
X"58805778",
X"882b7a07",
X"5680557a",
X"548353a3",
X"527c5192",
X"903f83c0",
X"800881ff",
X"0683c080",
X"0c8c3d0d",
X"04f73d0d",
X"02b30533",
X"028405b6",
X"0522605a",
X"58568055",
X"80548053",
X"81a3527b",
X"5191e23f",
X"83c08008",
X"81ff0683",
X"c0800c8b",
X"3d0d04ee",
X"3d0d6490",
X"115c5c80",
X"7b34800b",
X"841c0c80",
X"0b881c34",
X"810b891c",
X"34880b8a",
X"1c34800b",
X"8b1c3488",
X"1b08c106",
X"8107881c",
X"0c8f3d70",
X"545d8852",
X"7b519c92",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"81a93890",
X"3d335e81",
X"db5a7d89",
X"2e098106",
X"8199387c",
X"5392527b",
X"519beb3f",
X"83c08008",
X"81ff0670",
X"5b597881",
X"82387c58",
X"88577856",
X"a9557854",
X"865381a0",
X"527b5190",
X"d03f83c0",
X"800881ff",
X"06705b59",
X"7880e038",
X"02ba0533",
X"7b347c54",
X"78537d52",
X"7b519bd3",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"80c13802",
X"bd053352",
X"7b519beb",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"aa38817b",
X"335a5a79",
X"79269938",
X"80547953",
X"88527b51",
X"fdbb3f81",
X"1a7081ff",
X"067c3352",
X"5b59e439",
X"810b881c",
X"34805a79",
X"83c0800c",
X"943d0d04",
X"800b83c0",
X"800c04f9",
X"3d0d7902",
X"8405ab05",
X"338e3d70",
X"54585858",
X"ffafec3f",
X"8a3d8a05",
X"51ffafe3",
X"3f7551fc",
X"8d3f83c0",
X"80088486",
X"812ebe38",
X"83c08008",
X"84868126",
X"993883c0",
X"80088482",
X"802e80e6",
X"3883c080",
X"08848281",
X"2e9f3881",
X"b43983c0",
X"800880c0",
X"82832e80",
X"f43883c0",
X"800880c0",
X"86832e80",
X"e8388199",
X"3983c09c",
X"33558056",
X"74762e09",
X"8106818b",
X"38745476",
X"53915277",
X"51fbd63f",
X"74547653",
X"90527751",
X"fbcb3f74",
X"54765384",
X"527751fb",
X"fc3f810b",
X"83c09c34",
X"81b15680",
X"de398054",
X"76539152",
X"7751fba9",
X"3f805476",
X"53905277",
X"51fb9e3f",
X"800b83c0",
X"9c347652",
X"87183351",
X"97963fb5",
X"39805476",
X"53945277",
X"51fb823f",
X"80547653",
X"90527751",
X"faf73f75",
X"51ffae97",
X"3f83c080",
X"08892a81",
X"06537652",
X"87183351",
X"90cd3f80",
X"0b83c09c",
X"34805675",
X"83c0800c",
X"893d0d04",
X"f23d0d60",
X"90115a58",
X"800b881a",
X"33715956",
X"5674762e",
X"82a53882",
X"ac3f8419",
X"0883c080",
X"08268295",
X"3878335a",
X"810b8e3d",
X"23903df8",
X"1155f405",
X"53991852",
X"77518ae5",
X"3f83c080",
X"0881ff06",
X"70575574",
X"772e0981",
X"0681d938",
X"86397456",
X"81d23981",
X"5682578e",
X"3d337706",
X"5574802e",
X"bb38800b",
X"8d3d3490",
X"3df00554",
X"84537552",
X"7751facd",
X"3f83c080",
X"0881ff06",
X"55749d38",
X"7b537552",
X"7751fce7",
X"3f83c080",
X"0881ff06",
X"557481b1",
X"2e818b38",
X"74ffb338",
X"761081fc",
X"06811770",
X"81ff0658",
X"56578776",
X"27ffa838",
X"8156757a",
X"2680eb38",
X"800b8d3d",
X"348c3d70",
X"55578453",
X"75527751",
X"f9f73f83",
X"c0800881",
X"ff065574",
X"80c13876",
X"51ffac93",
X"3f83c080",
X"08828706",
X"55748281",
X"2e098106",
X"aa3802ae",
X"05338107",
X"55740284",
X"05ae0534",
X"7b537552",
X"7751fbeb",
X"3f83c080",
X"0881ff06",
X"557481b1",
X"2e903874",
X"feb83881",
X"167081ff",
X"065755ff",
X"91398056",
X"7581ff06",
X"56973f83",
X"c080088f",
X"d005841a",
X"0c755776",
X"83c0800c",
X"903d0d04",
X"049080a0",
X"0883c080",
X"0c04ff3d",
X"0d7387e8",
X"2951fefd",
X"dd3f833d",
X"0d040483",
X"cb840b83",
X"c0800c04",
X"fd3d0d75",
X"77545480",
X"0b83cae4",
X"34728a38",
X"9090800b",
X"84150c90",
X"3972812e",
X"09810688",
X"38909880",
X"0b84150c",
X"84140883",
X"cafc0c80",
X"0b88150c",
X"800b8c15",
X"0c83cafc",
X"0853820b",
X"87801434",
X"8151ff9e",
X"3f83cafc",
X"0853800b",
X"88143483",
X"cafc0853",
X"810b8780",
X"143483ca",
X"fc085380",
X"0b8c1434",
X"83cafc08",
X"53800ba4",
X"14349174",
X"34800b83",
X"c0a03480",
X"0b83c0a4",
X"34800b83",
X"c0a83480",
X"547381c4",
X"2983cb88",
X"0553800b",
X"83143481",
X"147081ff",
X"0655538f",
X"7427e638",
X"853d0d04",
X"fe3d0d74",
X"76821133",
X"70bf0681",
X"712bff05",
X"56515152",
X"53907127",
X"8338ff52",
X"76517171",
X"2383cafc",
X"08518713",
X"33901234",
X"800b83c0",
X"a434800b",
X"83c0a834",
X"8813338a",
X"14335252",
X"71802eaa",
X"387081ff",
X"06518452",
X"70833870",
X"527183c0",
X"a4348a13",
X"33703070",
X"8025842b",
X"70880751",
X"51525370",
X"83c0a834",
X"90397081",
X"ff065170",
X"83389852",
X"7183c0a8",
X"34800b83",
X"c0800c84",
X"3d0d04f1",
X"3d0d6165",
X"68028c05",
X"80cb0533",
X"02900580",
X"ce052202",
X"940580d6",
X"05224240",
X"415a4040",
X"fd8b3f83",
X"c08008a7",
X"88055b80",
X"70715b5b",
X"52839439",
X"83cafc08",
X"517d9412",
X"3483c0a4",
X"33810755",
X"80705456",
X"7f862680",
X"ea387f84",
X"2981efe0",
X"0583cafc",
X"08535170",
X"0804800b",
X"841334a1",
X"39773370",
X"30708025",
X"83713151",
X"51525370",
X"8413348d",
X"39810b84",
X"1334b839",
X"830b8413",
X"34817054",
X"56ad3981",
X"0b841334",
X"a2397733",
X"70307080",
X"25837131",
X"51515253",
X"70841334",
X"80783352",
X"52708338",
X"81527178",
X"34815374",
X"88075583",
X"c0a83383",
X"cafc0852",
X"57810b81",
X"d0123483",
X"cafc0851",
X"810b8190",
X"12347e80",
X"2eae3872",
X"802ea938",
X"7eff1e52",
X"547083ff",
X"ff065372",
X"83ffff2e",
X"97387370",
X"81055533",
X"83cafc08",
X"53517081",
X"c01334ff",
X"1351de39",
X"83cafc08",
X"a8113353",
X"51768812",
X"3483cafc",
X"08517471",
X"3481ff52",
X"913983ca",
X"fc08a011",
X"33708106",
X"51525370",
X"8f38fafd",
X"3f7a83c0",
X"800826e6",
X"38818839",
X"810ba014",
X"3483cafc",
X"08a81133",
X"80ff0670",
X"78075253",
X"5170802e",
X"80ed3871",
X"862a7081",
X"06515170",
X"802e9138",
X"80783352",
X"53708338",
X"81537278",
X"3480e039",
X"71842a70",
X"81065151",
X"70802e9b",
X"38811970",
X"83ffff06",
X"7d30709f",
X"2a51525a",
X"51787c2e",
X"098106af",
X"38a43971",
X"832a7081",
X"06515170",
X"802e9338",
X"811a7081",
X"ff065b51",
X"79832e09",
X"81069038",
X"8a3971a3",
X"06517080",
X"2e853871",
X"519239f9",
X"e43f7a83",
X"c0800826",
X"fce23871",
X"81bf0651",
X"7083c080",
X"0c913d0d",
X"04f63d0d",
X"02b30533",
X"028405b7",
X"05330288",
X"05ba0522",
X"59595980",
X"0b8c3d34",
X"8c3dfc05",
X"56805580",
X"54765377",
X"527851fb",
X"f23f83c0",
X"800881ff",
X"0683c080",
X"0c8c3d0d",
X"04f33d0d",
X"7f626402",
X"8c0580c2",
X"05227222",
X"81153342",
X"5f415e59",
X"59807823",
X"7d537833",
X"528151ff",
X"a03f83c0",
X"800881ff",
X"06567580",
X"2e863875",
X"5481ad39",
X"83cafc08",
X"a8113382",
X"1b337086",
X"2a708106",
X"73982b53",
X"51575c56",
X"57798025",
X"83388156",
X"73762e87",
X"3881f054",
X"81823981",
X"8c173370",
X"81ff0679",
X"227d7131",
X"902b7090",
X"2c700970",
X"9f2c7206",
X"70525253",
X"51535757",
X"54757424",
X"83387555",
X"74848080",
X"29fc8080",
X"0570902c",
X"515574ff",
X"2e943883",
X"cafc0881",
X"80113351",
X"54737c70",
X"81055e34",
X"db397722",
X"76055473",
X"78237909",
X"709f2a70",
X"8106821c",
X"3381bf06",
X"71862b07",
X"51515154",
X"73821a34",
X"7c76268a",
X"38772254",
X"7a7426fe",
X"bb388054",
X"7383c080",
X"0c8f3d0d",
X"04f93d0d",
X"7a57800b",
X"893d2389",
X"3dfc0553",
X"76527951",
X"f8da3f83",
X"c0800881",
X"ff067057",
X"55749638",
X"7c547b53",
X"883d2252",
X"7651fde5",
X"3f83c080",
X"0881ff06",
X"567583c0",
X"800c893d",
X"0d04f03d",
X"0d626602",
X"880580ce",
X"0522415d",
X"5e800284",
X"0580d205",
X"227f8105",
X"33ff115a",
X"5d5a5d81",
X"da5876bf",
X"2680e938",
X"78802e80",
X"e1387a58",
X"787b2783",
X"38785882",
X"1e337087",
X"2a585a76",
X"923d3492",
X"3dfc0556",
X"77557b54",
X"7e537d33",
X"528251f8",
X"de3f83c0",
X"800881ff",
X"065d800b",
X"923d3358",
X"5a76802e",
X"8338815a",
X"821e3380",
X"ff067a87",
X"2b075776",
X"821f347c",
X"91387878",
X"317083ff",
X"ff06791e",
X"5e5a57ff",
X"9b397c58",
X"7783c080",
X"0c923d0d",
X"04f83d0d",
X"7b028405",
X"b2052258",
X"58800b8a",
X"3d238a3d",
X"fc055377",
X"527a51f6",
X"f73f83c0",
X"800881ff",
X"06705755",
X"7496387d",
X"54765389",
X"3d225277",
X"51feaf3f",
X"83c08008",
X"81ff0656",
X"7583c080",
X"0c8a3d0d",
X"04ec3d0d",
X"666e0288",
X"0580df05",
X"33028c05",
X"80e30533",
X"02900580",
X"e7053302",
X"940580eb",
X"05330298",
X"0580ee05",
X"22414341",
X"5f5c4057",
X"0280f205",
X"22963d23",
X"963df005",
X"53841770",
X"53775259",
X"f6863f83",
X"c0800881",
X"ff065877",
X"81e53877",
X"7a818006",
X"58408077",
X"25833881",
X"4079943d",
X"347b0284",
X"0580c905",
X"347c0284",
X"0580ca05",
X"347d0284",
X"0580cb05",
X"347a953d",
X"347a882a",
X"57760284",
X"0580cd05",
X"34953d22",
X"57760284",
X"0580ce05",
X"3476882a",
X"57760284",
X"0580cf05",
X"3477923d",
X"34963dec",
X"11575788",
X"55f41754",
X"923d2253",
X"77527751",
X"f6953f83",
X"c0800881",
X"ff065877",
X"80ed387e",
X"802e80cb",
X"38923d22",
X"79085858",
X"7f802e9c",
X"38768180",
X"8007790c",
X"7e54963d",
X"fc055377",
X"83ffff06",
X"527851f9",
X"fc3f9939",
X"76828080",
X"07790c7e",
X"54953d22",
X"537783ff",
X"ff065278",
X"51fc8f3f",
X"83c08008",
X"81ff0658",
X"779d3892",
X"3d225380",
X"527f3070",
X"80258471",
X"31535157",
X"f9873f83",
X"c0800881",
X"ff065877",
X"83c0800c",
X"963d0d04",
X"f63d0d7c",
X"028405b7",
X"05335b5b",
X"80588057",
X"80568055",
X"79548553",
X"80527a51",
X"fda33f83",
X"c0800881",
X"ff065978",
X"85387987",
X"1c347883",
X"c0800c8c",
X"3d0d04f9",
X"3d0d02a7",
X"05330284",
X"05ab0533",
X"028805af",
X"05335859",
X"57800b83",
X"cb8b3354",
X"5472742e",
X"9f388114",
X"7081ff06",
X"5553738f",
X"2681b638",
X"7381c429",
X"83cb8805",
X"83113351",
X"5372e338",
X"7381c429",
X"83cb8405",
X"55800b87",
X"16347688",
X"1634758a",
X"16347789",
X"16348075",
X"0c83cafc",
X"088c160c",
X"800b8416",
X"34880b85",
X"1634800b",
X"86163484",
X"1508ffa1",
X"ff06a080",
X"0784160c",
X"81147081",
X"ff065353",
X"7451febc",
X"3f83c080",
X"0881ff06",
X"70555372",
X"80cd388a",
X"39730875",
X"0c725480",
X"c2397281",
X"f7805556",
X"81f78008",
X"802eb238",
X"75842914",
X"70087653",
X"70085154",
X"54722d83",
X"c0800881",
X"ff065372",
X"802ece38",
X"81167081",
X"ff0681f7",
X"80718429",
X"11535657",
X"537208d0",
X"38805473",
X"83c0800c",
X"893d0d04",
X"f93d0d79",
X"57800b84",
X"180883ca",
X"fc0c58f0",
X"883f8817",
X"0883c080",
X"082783ed",
X"38effa3f",
X"83c08008",
X"81058818",
X"0c83cafc",
X"08b81133",
X"7081ff06",
X"51515473",
X"812ea438",
X"73812488",
X"3873782e",
X"8a38b839",
X"73822e95",
X"38b13976",
X"3381f006",
X"5473902e",
X"a6389177",
X"34a13973",
X"58763381",
X"f0065473",
X"902e0981",
X"069138ef",
X"a83f83c0",
X"800881c8",
X"058c180c",
X"a0773480",
X"567581c4",
X"2983cb8b",
X"11335555",
X"73802eaa",
X"3883cb84",
X"15700856",
X"5474802e",
X"9d388815",
X"08802e96",
X"388c1408",
X"83cafc08",
X"2e098106",
X"89387351",
X"88150854",
X"732d8116",
X"7081ff06",
X"57548f76",
X"27ffba38",
X"76335473",
X"b02e8199",
X"3873b024",
X"8f387391",
X"2eab3873",
X"a02e80f5",
X"3882a639",
X"7380d02e",
X"81e43873",
X"80d0248b",
X"387380c0",
X"2e819938",
X"828f3973",
X"81802e81",
X"fb388285",
X"39805675",
X"81c42983",
X"cb881183",
X"11335659",
X"5573802e",
X"a83883cb",
X"84157008",
X"56547480",
X"2e9b388c",
X"140883ca",
X"fc082e09",
X"81068e38",
X"73518415",
X"0854732d",
X"800b8319",
X"34811670",
X"81ff0657",
X"548f7627",
X"ffb93892",
X"773481b5",
X"39edc23f",
X"8c170883",
X"c0800827",
X"81a738b0",
X"773481a1",
X"3983cafc",
X"0854800b",
X"8c153483",
X"cafc0854",
X"840b8815",
X"3480c077",
X"34ed963f",
X"83c08008",
X"b2058c18",
X"0c80fa39",
X"ed873f8c",
X"170883c0",
X"80082780",
X"ec3883ca",
X"fc085481",
X"0b8c1534",
X"83cafc08",
X"54800b88",
X"153483ca",
X"fc085488",
X"0ba01534",
X"ecdb3f83",
X"c0800894",
X"058c180c",
X"80d07734",
X"bc3983ca",
X"fc08a011",
X"3370832a",
X"70810651",
X"51555573",
X"802ea638",
X"880ba016",
X"34ecae3f",
X"8c170883",
X"c0800827",
X"9438ff80",
X"77348e39",
X"77538052",
X"8051fa8b",
X"3fff9077",
X"3483cafc",
X"08a01133",
X"70832a70",
X"81065151",
X"55557380",
X"2e863888",
X"0ba01634",
X"893d0d04",
X"f43d0d02",
X"bb053302",
X"8405bf05",
X"335d5d80",
X"0b83cb88",
X"0b83cb84",
X"0b8c1172",
X"71881475",
X"5c5a5b5f",
X"5c595b58",
X"83153353",
X"72802e81",
X"88387333",
X"537c732e",
X"09810680",
X"fc388114",
X"33537b73",
X"2e098106",
X"80ef3875",
X"0883cafc",
X"082e0981",
X"0680e238",
X"80567581",
X"c42983cb",
X"8c117033",
X"831e335b",
X"57555374",
X"782e0981",
X"06973883",
X"cb901308",
X"79082e09",
X"81068a38",
X"81143352",
X"7451fef8",
X"3f811670",
X"81ff0657",
X"538f7627",
X"c5388077",
X"08545472",
X"742e9138",
X"76518413",
X"0853722d",
X"83c08008",
X"81ff0654",
X"800b831b",
X"347353a9",
X"39811881",
X"c41681c4",
X"1681c419",
X"81c41f81",
X"c41e81c4",
X"1d6081c4",
X"05415d5e",
X"5f595656",
X"588f7825",
X"feca3880",
X"537283c0",
X"800c8e3d",
X"0d04f83d",
X"0d02ae05",
X"227d5957",
X"80568155",
X"80548653",
X"8180527a",
X"51f4ee3f",
X"83c08008",
X"81ff0683",
X"c0800c8a",
X"3d0d04f7",
X"3d0d02b2",
X"05220284",
X"05b70533",
X"605a5b57",
X"80568255",
X"79548653",
X"8180527b",
X"51f4be3f",
X"83c08008",
X"81ff0683",
X"c0800c8b",
X"3d0d04f8",
X"3d0d02af",
X"05335980",
X"58805780",
X"56805578",
X"54895380",
X"527a51f4",
X"943f83c0",
X"800881ff",
X"0683c080",
X"0c8a3d0d",
X"04ffb83d",
X"0d80cb3d",
X"08705381",
X"f3bc5256",
X"feaaf73f",
X"83c08008",
X"80f33875",
X"51fea4e2",
X"3f83ffff",
X"0b83c080",
X"082580e1",
X"387551fe",
X"a4e13f83",
X"c0800855",
X"83c08008",
X"80cf3882",
X"805383c0",
X"8008528a",
X"3d705257",
X"fee6b83f",
X"74527551",
X"fea3f23f",
X"805980ca",
X"3dfdfc05",
X"54828053",
X"76527551",
X"fea1f93f",
X"81155574",
X"88802e09",
X"8106e138",
X"80527551",
X"fea3ca3f",
X"800b83e3",
X"c80c7583",
X"e3c40c87",
X"39800b83",
X"e3c40c80",
X"ca3d0d04",
X"ff3d0d73",
X"70085351",
X"02930533",
X"72347008",
X"8105710c",
X"833d0d04",
X"ffb83d0d",
X"80cb3d70",
X"70840552",
X"08585683",
X"e3c40880",
X"2e80fa38",
X"8a3d705a",
X"76557754",
X"81e9b053",
X"80cb3dfd",
X"fc055255",
X"fed0883f",
X"805280ca",
X"3dfdfc05",
X"51ffad3f",
X"83e3c808",
X"5283e3c4",
X"0851fea2",
X"d03f8058",
X"7451fecd",
X"ce3f80ca",
X"3dfdf805",
X"5483c080",
X"08537452",
X"83e3c408",
X"51fea0cc",
X"3f83e3c8",
X"081883e3",
X"c80c80ca",
X"3dfdf805",
X"54815381",
X"f3c85283",
X"e3c40851",
X"fea0ad3f",
X"83e3c808",
X"1883e3c8",
X"0c80ca3d",
X"0d040000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002d46",
X"00002d87",
X"00002da9",
X"00002dcb",
X"00002df1",
X"00002df1",
X"00002df1",
X"00002df1",
X"00002e62",
X"00002eb3",
X"00002ebd",
X"00004477",
X"00004e97",
X"00004f60",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3f00",
X"0c0c4000",
X"0a0a4100",
X"0b0b4100",
X"07074100",
X"0a0b4300",
X"080b4200",
X"06060004",
X"04044500",
X"05054400",
X"0e0f2900",
X"08080004",
X"09090004",
X"0a0f4300",
X"090f4200",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"00006144",
X"0000644b",
X"00006257",
X"0000644b",
X"00006294",
X"000062e5",
X"00006324",
X"0000632d",
X"0000644b",
X"0000644b",
X"0000644b",
X"0000644b",
X"00006336",
X"0000633e",
X"00006345",
X"0000654b",
X"00006644",
X"00006758",
X"00006a4e",
X"00006a69",
X"00006a55",
X"00006a69",
X"00006a70",
X"00006a7b",
X"00006a82",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"25782e48",
X"75622e20",
X"25642070",
X"6f727473",
X"00000000",
X"25782e48",
X"49440000",
X"204d6f75",
X"73650000",
X"204b6579",
X"626f6172",
X"64000000",
X"204a6f79",
X"73746963",
X"6b3a2564",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"43505520",
X"54757262",
X"6f3a2564",
X"78000000",
X"44726976",
X"65205475",
X"72626f3a",
X"25730000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"526f7461",
X"74652055",
X"5342206a",
X"6f797374",
X"69636b73",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"66726565",
X"7a65722e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"4d454d00",
X"5374616e",
X"64617264",
X"00000000",
X"46617374",
X"28362900",
X"46617374",
X"28352900",
X"46617374",
X"28342900",
X"46617374",
X"28332900",
X"46617374",
X"28322900",
X"46617374",
X"28312900",
X"46617374",
X"28302900",
X"2f757362",
X"2e6c6f67",
X"00000000",
X"0a000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"0000787c",
X"00007880",
X"00007888",
X"00007894",
X"000078a0",
X"000078ac",
X"000078b8",
X"000078bc",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00000028",
X"00000006",
X"00000005",
X"00000004",
X"00000003",
X"00000002",
X"00000001",
X"00000000",
X"00007978",
X"00007984",
X"0000798c",
X"00007994",
X"0000799c",
X"000079a4",
X"000079ac",
X"000079b4",
X"000077d4",
X"0000761c",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"69383030",
X"00000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
