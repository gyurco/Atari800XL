-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 12.1 Build 243 01/31/2013 Service Pack 1.33 SJ Web Edition"
-- CREATED		"Tue Dec 31 22:21:48 2013"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 
use IEEE.STD_LOGIC_MISC.all;
use ieee.numeric_std.all;

LIBRARY work;

ENTITY atari800core IS 
	PORT
	(
		CLK :  IN  STD_LOGIC;
		PLL_LOCKED: IN STD_LOGIC;

		VGA_VS :  OUT  STD_LOGIC;
		VGA_HS :  OUT  STD_LOGIC;
		VGA_B :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		VGA_G :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		VGA_R :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		
		JOY1_n :  IN  STD_LOGIC_VECTOR(5 DOWNTO 0);
		JOY2_n :  IN  STD_LOGIC_VECTOR(5 DOWNTO 0);

		matrix_out : in std_logic_vector(15 downto 0);
		matrix_in : out std_logic_vector(7 downto 0);
		static_keys : in std_logic_vector(6 downto 0);
		pause_key : in std_logic;
		
		AUDIO_L : OUT std_logic_vector(15 downto 0);
		AUDIO_R : OUT std_logic_vector(15 downto 0);

		SDRAM_REQUEST : OUT std_logic;
		SDRAM_REQUEST_COMPLETE : IN std_logic;
		SDRAM_READ_ENABLE : out STD_LOGIC;
		SDRAM_WRITE_ENABLE : out std_logic;
		SDRAM_DI : out std_logic_vector(31 downto 0);
		SDRAM_ADDR : out STD_LOGIC_VECTOR(22 DOWNTO 0);
		SDRAM_DO : in STD_LOGIC_VECTOR(31 DOWNTO 0);
		SDRAM_WIDTH_8bit_ACCESS : out std_logic;
		SDRAM_WIDTH_16bit_ACCESS : out std_logic;
		SDRAM_WIDTH_32bit_ACCESS : out std_logic;

		SIO_RXD : in std_logic;
		SIO_TXD : out std_logic;
		SIO_COMMAND_TX : out std_logic;

   		ram_select : in std_logic_vector(2 downto 0);
    		rom_select : in std_logic_vector(5 downto 0);

		halt : in std_logic
	);
END atari800core;

ARCHITECTURE bdf_type OF atari800core IS 
component synchronizer IS
PORT 
( 
	CLK : IN STD_LOGIC;
	RAW : IN STD_LOGIC;
	SYNC : OUT STD_LOGIC
);
END component;

COMPONENT complete_address_decoder IS
generic (width : natural := 1);
PORT 
( 
	addr_in : in std_logic_vector(width-1 downto 0);			
	addr_decoded : out std_logic_vector((2**width)-1 downto 0)
);
END component;

COMPONENT cpu
	PORT(CLK : IN STD_LOGIC;
		 RESET : IN STD_LOGIC;
		 ENABLE : IN STD_LOGIC;
		 IRQ_n : IN STD_LOGIC;
		 NMI_n : IN STD_LOGIC;
		 MEMORY_READY : IN STD_LOGIC;
		 THROTTLE : IN STD_LOGIC;
		 RDY : IN STD_LOGIC;
		 DI : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 R_W_n : OUT STD_LOGIC;
		 CPU_FETCH : OUT STD_LOGIC;
		 A : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 DO : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

component internalromram IS
  PORT(
    clock   : IN     STD_LOGIC;                             --system clock
    reset_n : IN     STD_LOGIC;                             --asynchronous reset

	ROM_ADDR : in STD_LOGIC_VECTOR(21 downto 0);
	ROM_REQUEST_COMPLETE : out STD_LOGIC;
	ROM_REQUEST : in std_logic;
	ROM_DATA : out std_logic_vector(7 downto 0);
	
	RAM_ADDR : in STD_LOGIC_VECTOR(18 downto 0);
	RAM_WR_ENABLE : in std_logic;
	RAM_DATA_IN : in STD_LOGIC_VECTOR(7 downto 0);
	RAM_REQUEST_COMPLETE : out STD_LOGIC;
	RAM_REQUEST : in std_logic;
	RAM_DATA : out std_logic_vector(7 downto 0)
	);
	
END component;

COMPONENT antic
	PORT(CLK : IN STD_LOGIC;
		 WR_EN : IN STD_LOGIC;
		 RESET_N : IN STD_LOGIC;
		 MEMORY_READY_ANTIC : IN STD_LOGIC;
		 MEMORY_READY_CPU : IN STD_LOGIC;
		 ANTIC_ENABLE_179 : IN STD_LOGIC;
		 PAL : IN STD_LOGIC;
		 lightpen : IN STD_LOGIC;
		 ADDR : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 CPU_DATA_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 MEMORY_DATA_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 NMI_N_OUT : OUT STD_LOGIC;
		 ANTIC_READY : OUT STD_LOGIC;
		 COLOUR_CLOCK_ORIGINAL_OUT : OUT STD_LOGIC;
		 COLOUR_CLOCK_OUT : OUT STD_LOGIC;
		 HIGHRES_COLOUR_CLOCK_OUT : OUT STD_LOGIC;
		 dma_fetch_out : OUT STD_LOGIC;
		 refresh_out : OUT STD_LOGIC;
		 dma_clock_out : OUT STD_LOGIC;
		 hcount_out : out std_logic_vector(7 downto 0);
		 vcount_out : out std_logic_vector(8 downto 0);
		 AN : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 DATA_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 dma_address_out : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT pokey_mixer
	PORT(CLK : IN STD_LOGIC;
		 GTIA_SOUND : IN STD_LOGIC;
		 CHANNEL_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 CHANNEL_1 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 CHANNEL_2 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 CHANNEL_3 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 COVOX_CHANNEL_0 : IN STD_LOGIC_VECTOR(7 downto 0);
		 COVOX_CHANNEL_1 : IN STD_LOGIC_VECTOR(7 downto 0);
		 CHANNEL_ENABLE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 VOLUME_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT zpu_glue
	PORT(CLK : IN STD_LOGIC;
		 RESET : IN STD_LOGIC;
		 PAUSE : IN STD_LOGIC;
		 MEMORY_READY : IN STD_LOGIC;
		 ZPU_CONFIG_DI : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 ZPU_DI : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 ZPU_RAM_DI : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 ZPU_ROM_DI : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 ZPU_SECTOR_DI : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 MEMORY_FETCH : OUT STD_LOGIC;
		 ZPU_READ_ENABLE : OUT STD_LOGIC;
		 ZPU_32BIT_WRITE_ENABLE : OUT STD_LOGIC;
		 ZPU_16BIT_WRITE_ENABLE : OUT STD_LOGIC;
		 ZPU_8BIT_WRITE_ENABLE : OUT STD_LOGIC;
		 ZPU_CONFIG_WRITE : OUT STD_LOGIC;
		 ZPU_ADDR_FETCH : OUT STD_LOGIC_VECTOR(23 DOWNTO 0);
		 ZPU_ADDR_ROM_RAM : OUT STD_LOGIC_VECTOR(23 DOWNTO 0);
		 ZPU_DO : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 ZPU_STACK_WRITE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT pokey
	PORT(CLK : IN STD_LOGIC;
		 CPU_MEMORY_READY : IN STD_LOGIC;
		 ANTIC_MEMORY_READY : IN STD_LOGIC;
		 WR_EN : IN STD_LOGIC;
		 RESET_N : IN STD_LOGIC;
		 SIO_IN1 : IN STD_LOGIC;
		 SIO_IN2 : IN STD_LOGIC;
		 SIO_IN3 : IN STD_LOGIC;
		 SIO_CLOCK : INOUT STD_LOGIC;
		 ADDR : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 DATA_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 keyboard_response : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 POT_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 IRQ_N_OUT : OUT STD_LOGIC;
		 SIO_OUT1 : OUT STD_LOGIC;
		 SIO_OUT2 : OUT STD_LOGIC;
		 SIO_OUT3 : OUT STD_LOGIC;
		 POT_RESET : OUT STD_LOGIC;
		 CHANNEL_0_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 CHANNEL_1_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 CHANNEL_2_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 CHANNEL_3_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 DATA_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 keyboard_scan : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END COMPONENT;

COMPONENT pia
	PORT(	CLK : IN STD_LOGIC;
	ADDR : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
	CPU_DATA_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	EN : IN STD_LOGIC;
	WR_EN : IN STD_LOGIC;
	
	RESET_N : IN STD_LOGIC;
	
	CA1 : IN STD_LOGIC;
	CB1 : IN STD_LOGIC;		
	
	CA2_DIR_OUT : OUT std_logic;
	CA2_OUT : OUT std_logic;
	CA2_IN : IN STD_LOGIC;

	CB2_DIR_OUT : OUT std_logic;
	CB2_OUT : OUT std_logic;
	CB2_IN : IN STD_LOGIC;
	
	-- remember these two are different if connecting to gpio (push pull vs pull up - check 6520 data sheet...)
	-- pull up - i.e. 0 driven only
	PORTA_DIR_OUT : OUT STD_LOGIC_VECTOR(7 downto 0); -- set bit to 1 to enable output mode
	PORTA_OUT : OUT STD_LOGIC_VECTOR(7 downto 0); 
	PORTA_IN : IN STD_LOGIC_VECTOR(7 downto 0);
	
	PORTB_DIR_OUT : OUT STD_LOGIC_VECTOR(7 downto 0);
	PORTB_OUT : OUT STD_LOGIC_VECTOR(7 downto 0); -- push pull
	PORTB_IN : IN STD_LOGIC_VECTOR(7 downto 0); -- push pull
	
	-- CPU interface
	DATA_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		
	IRQA_N : OUT STD_LOGIC;
	IRQB_N : OUT STD_LOGIC	);
END COMPONENT;

COMPONENT shared_enable
	PORT(CLK : IN STD_LOGIC;
		 RESET_N : IN STD_LOGIC;
		 MEMORY_READY_CPU : IN STD_LOGIC;
		 MEMORY_READY_ANTIC : IN STD_LOGIC;
		 PAUSE_6502 : IN STD_LOGIC;
		 THROTTLE_COUNT_6502 : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		 POKEY_ENABLE_179 : OUT STD_LOGIC;
		 ANTIC_ENABLE_179 : OUT STD_LOGIC;
		 oldcpu_enable : OUT STD_LOGIC;
		 CPU_ENABLE_OUT : OUT STD_LOGIC;
		 SCANDOUBLER_ENABLE_LOW : OUT STD_LOGIC;
		 SCANDOUBLER_ENABLE_HIGH : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT address_decoder
	PORT(CLK : IN STD_LOGIC;
		 CPU_FETCH : IN STD_LOGIC;
		 CPU_WRITE_N : IN STD_LOGIC;
		 ANTIC_FETCH : IN STD_LOGIC;
		 antic_refresh : IN STD_LOGIC;
		 ZPU_FETCH : IN STD_LOGIC;
		 ZPU_READ_ENABLE : IN STD_LOGIC;
		 ZPU_32BIT_WRITE_ENABLE : IN STD_LOGIC;
		 ZPU_16BIT_WRITE_ENABLE : IN STD_LOGIC;
		 ZPU_8BIT_WRITE_ENABLE : IN STD_LOGIC;
		 RAM_REQUEST_COMPLETE : IN STD_LOGIC;
		 ROM_REQUEST_COMPLETE : IN STD_LOGIC;
		 CART_REQUEST_COMPLETE : IN STD_LOGIC;
		 reset_n : IN STD_LOGIC;
		 CART_RD4 : IN STD_LOGIC;
		 CART_RD5 : IN STD_LOGIC;
		 use_sdram : IN STD_LOGIC;
		 SDRAM_REQUEST_COMPLETE : IN STD_LOGIC;
		 ANTIC_ADDR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 ANTIC_DATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 CACHE_ANTIC_DATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 CART_ROM_DATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 CPU_ADDR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 CPU_WRITE_DATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 GTIA_DATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 CACHE_GTIA_DATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 PIA_DATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 POKEY2_DATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 CACHE_POKEY2_DATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 POKEY_DATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 CACHE_POKEY_DATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 PORTB : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 RAM_DATA : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 ram_select : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 ROM_DATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 rom_select : in std_logic_vector(5 downto 0);
		 cart_select : in std_logic_vector(6 downto 0);
		 cart_activate : in std_logic;
		 SDRAM_DATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 ZPU_ADDR : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
		 ZPU_WRITE_DATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 MEMORY_READY_ANTIC : OUT STD_LOGIC;
		 MEMORY_READY_ZPU : OUT STD_LOGIC;
		 MEMORY_READY_CPU : OUT STD_LOGIC;
		 GTIA_WR_ENABLE : OUT STD_LOGIC;
		 POKEY_WR_ENABLE : OUT STD_LOGIC;
		 POKEY2_WR_ENABLE : OUT STD_LOGIC;
		 ANTIC_WR_ENABLE : OUT STD_LOGIC;
		 PIA_WR_ENABLE : OUT STD_LOGIC;
		 PIA_RD_ENABLE : OUT STD_LOGIC;
		 RAM_WR_ENABLE : OUT STD_LOGIC;
		 PBI_WR_ENABLE : OUT STD_LOGIC;
		 RAM_REQUEST : OUT STD_LOGIC;
		 ROM_REQUEST : OUT STD_LOGIC;
		 CART_REQUEST : OUT STD_LOGIC;
		 CART_S4_n : OUT STD_LOGIC;
		 CART_S5_n : OUT STD_LOGIC;
		 CART_CCTL_n : OUT STD_LOGIC;
		 WIDTH_8bit_ACCESS : OUT STD_LOGIC;
		 WIDTH_16bit_ACCESS : OUT STD_LOGIC;
		 WIDTH_32bit_ACCESS : OUT STD_LOGIC;
		 SDRAM_READ_EN : OUT STD_LOGIC;
		 SDRAM_WRITE_EN : OUT STD_LOGIC;
		 SDRAM_REQUEST : OUT STD_LOGIC;
		 SDRAM_REFRESH : OUT STD_LOGIC;
		 MEMORY_DATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 PBI_ADDR : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 RAM_ADDR : OUT STD_LOGIC_VECTOR(18 DOWNTO 0);
		 ROM_ADDR : OUT STD_LOGIC_VECTOR(21 DOWNTO 0);
		 SDRAM_ADDR : OUT STD_LOGIC_VECTOR(22 DOWNTO 0);
		 WRITE_DATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 D6_WR_ENABLE : out std_logic
	);
END COMPONENT;

COMPONENT zpu_rom
	PORT(clock : IN STD_LOGIC;
		 address : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

--COMPONENT zpu_ram
--	PORT(wren : IN STD_LOGIC;
--		 clock : IN STD_LOGIC;
--		 address : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
--		 data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
--		 q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
--	);
--END COMPONENT;

component generic_ram_infer IS
        generic
        (
                ADDRESS_WIDTH : natural := 9;
                SPACE : natural := 512;
                DATA_WIDTH : natural := 8
        );
   PORT
   (
      clock: IN   std_logic;
      data:  IN   std_logic_vector (data_width-1 DOWNTO 0);
      address:  IN   std_logic_vector(address_width-1 downto 0);
      we:    IN   std_logic;
      q:     OUT  std_logic_vector (data_width-1 DOWNTO 0)
   );
END component;

COMPONENT zpu_config_regs
	PORT(CLK : IN STD_LOGIC;
		 ENABLE_179 : IN STD_LOGIC;
		 WR_EN : IN STD_LOGIC;
		 SDCARD_DAT : IN STD_LOGIC;
		 SIO_COMMAND_OUT : IN STD_LOGIC;
		 SIO_DATA_OUT : IN STD_LOGIC;
		 PLL_LOCKED : IN STD_LOGIC;
		 REQUEST_RESET_ZPU : IN STD_LOGIC;
		 ADDR : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 CPU_DATA_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 KEY : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 SWITCH : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		 SDCARD_CLK : OUT STD_LOGIC;
		 SDCARD_CMD : OUT STD_LOGIC;
		 SDCARD_DAT3 : OUT STD_LOGIC;
		 SIO_DATA_IN : OUT STD_LOGIC;
		 PAUSE_ZPU : OUT STD_LOGIC;
		 PAL : OUT STD_LOGIC;
		 USE_SDRAM : OUT STD_LOGIC;
		 VGA : OUT STD_LOGIC;
		 COMPOSITE_ON_HSYNC : OUT STD_LOGIC;
		 GPIO_ENABLE : OUT STD_LOGIC;
		 RESET_6502 : OUT STD_LOGIC;
		 RESET_ZPU : OUT STD_LOGIC;
		 RESET_N : OUT STD_LOGIC;
		 PAUSE_6502 : OUT STD_LOGIC;
		 DATA_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 LEDG : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 LEDR : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		 RAM_SELECT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 ROM_SELECT : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		 THROTTLE_COUNT_6502 : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		 ZPU_HEX : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 sector : out std_logic_vector(31 downto 0);
		 sector_request : out std_logic;
		 sector_ready : in std_logic
	);
END COMPONENT;

COMPONENT gtia_palette IS
PORT 
( 
	ATARI_COLOUR : IN STD_LOGIC_VECTOR(7 downto 0);
	
	R_next : OUT STD_LOGIC_VECTOR(7 downto 0);
	G_next : OUT STD_LOGIC_VECTOR(7 downto 0);
	B_next : OUT STD_LOGIC_VECTOR(7 downto 0)
);
END component;

COMPONENT gtia
	PORT(CLK : IN STD_LOGIC;
		 WR_EN : IN STD_LOGIC;
		 CPU_MEMORY_READY : IN STD_LOGIC;
		 ANTIC_MEMORY_READY : IN STD_LOGIC;
		 ANTIC_FETCH : IN STD_LOGIC;
		 CPU_ENABLE_ORIGINAL : IN STD_LOGIC;
		 RESET_N : IN STD_LOGIC;
		 PAL : IN STD_LOGIC;
		 COLOUR_CLOCK_ORIGINAL : IN STD_LOGIC;
		 COLOUR_CLOCK : IN STD_LOGIC;
		 COLOUR_CLOCK_HIGHRES : IN STD_LOGIC;
		 CONSOL_START : IN STD_LOGIC;
		 CONSOL_SELECT : IN STD_LOGIC;
		 CONSOL_OPTION : IN STD_LOGIC;
		 TRIG0 : IN STD_LOGIC;
		 TRIG1 : IN STD_LOGIC;
		 TRIG2 : IN STD_LOGIC;
		 TRIG3 : IN STD_LOGIC;
		 ADDR : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 AN : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 CPU_DATA_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 MEMORY_DATA_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 VSYNC : OUT STD_LOGIC;
		 HSYNC : OUT STD_LOGIC;
		 BLANK : OUT STD_LOGIC;
		 sound : OUT STD_LOGIC;
		 COLOUR_out : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 DATA_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT irq_glue
	PORT(pokey_irq : IN STD_LOGIC;
		 pia_irqa : IN STD_LOGIC;
		 pia_irqb : IN STD_LOGIC;
		 combined_irq : OUT STD_LOGIC
	);
END COMPONENT;

component reg_file IS
generic
(
	BYTES : natural := 1;
	WIDTH : natural := 1
);
PORT 
( 
	CLK : IN STD_LOGIC;
	ADDR : IN STD_LOGIC_VECTOR(width-1 DOWNTO 0);
	DATA_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	WR_EN : IN STD_LOGIC;
	
	DATA_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END component;

component covox IS
PORT 
( 
	CLK : IN STD_LOGIC;
	ADDR : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
	DATA_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	WR_EN : IN STD_LOGIC;
	
	covox_channel0 : out std_logic_vector(7 downto 0);
	covox_channel1 : out std_logic_vector(7 downto 0);
	covox_channel2 : out std_logic_vector(7 downto 0);
	covox_channel3 : out std_logic_vector(7 downto 0)
);
END component;



SIGNAL	ANTIC_ADDR :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	ANTIC_AN :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	ANTIC_COLOUR_CLOCK_OUT :  STD_LOGIC;
SIGNAL	ANTIC_DO :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	CACHE_ANTIC_DO :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	ANTIC_ENABLE_179 :  STD_LOGIC;
SIGNAL	ANTIC_FETCH :  STD_LOGIC;
SIGNAL	ANTIC_HIGHRES_COLOUR_CLOCK_OUT :  STD_LOGIC;
SIGNAL	ANTIC_ORIGINAL_COLOUR_CLOCK_OUT :  STD_LOGIC;
SIGNAL	ANTIC_RDY :  STD_LOGIC;
SIGNAL	ANTIC_REFRESH :  STD_LOGIC;
SIGNAL	ANTIC_WRITE_ENABLE :  STD_LOGIC;
SIGNAL	BREAK_PRESSED :  STD_LOGIC;

SIGNAL	CART_RD4 :  STD_LOGIC;
SIGNAL	CART_RD5 :  STD_LOGIC;
SIGNAL	CART_REQUEST :  STD_LOGIC;
SIGNAL	CART_REQUEST_COMPLETE :  STD_LOGIC;
SIGNAL	CART_ROM_DO :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	CART_S4_n :  STD_LOGIC;
SIGNAL	CART_S5_N :  STD_LOGIC;
signal CART_CCTL_N : std_logic;
SIGNAL	CA2_OUT :  STD_LOGIC;
SIGNAL	CA2_DIR_OUT:  STD_LOGIC;
SIGNAL	CB2_OUT :  STD_LOGIC;
SIGNAL	CB2_DIR_OUT:  STD_LOGIC;
SIGNAL	COMPOSITE_ON_HSYNC :  STD_LOGIC;
SIGNAL	CONSOL_OPTION :  STD_LOGIC;
SIGNAL	CONSOL_SELECT :  STD_LOGIC;
SIGNAL	CONSOL_START :  STD_LOGIC;
SIGNAL	CPU_6502_RESET :  STD_LOGIC;
SIGNAL	CPU_ADDR :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	CPU_DO :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	CPU_FETCH :  STD_LOGIC;
SIGNAL	CPU_SHARED_ENABLE :  STD_LOGIC;
SIGNAL	ENABLE_179_MEMWAIT :  STD_LOGIC;
SIGNAL   GPIO_0_IN : STD_LOGIC_VECTOR(35 downto 0);
SIGNAL   GPIO_0_OUT : STD_LOGIC_VECTOR(35 downto 0);
SIGNAL   GPIO_0_DIR_OUT : STD_LOGIC_VECTOR(35 downto 0);
SIGNAL   GPIO_1_IN : STD_LOGIC_VECTOR(35 downto 0);
SIGNAL   GPIO_1_OUT : STD_LOGIC_VECTOR(35 downto 0);
SIGNAL   GPIO_1_DIR_OUT : STD_LOGIC_VECTOR(35 downto 0);
SIGNAL	GPIO_CA2_IN:  STD_LOGIC;
SIGNAL	GPIO_CB2_IN:  STD_LOGIC;
SIGNAL	GPIO_ENABLE :  STD_LOGIC;
SIGNAL	GPIO_PORTA_IN :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	GPIO_PORTB_IN :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL   GPIO_SIO_IN : STD_LOGIC;
SIGNAL   GPIO_SIO_OUT : STD_LOGIC;
SIGNAL	GREEN_LEDS :  STD_LOGIC_VECTOR(1 TO 1);
SIGNAL	GREREN_LEDS :  STD_LOGIC_VECTOR(0 TO 0);
SIGNAL	GTIA_DO :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	CACHE_GTIA_DO :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	GTIA_SOUND :  STD_LOGIC;
SIGNAL	GTIA_WRITE_ENABLE :  STD_LOGIC;
SIGNAL	IRQ_n :  STD_LOGIC;
SIGNAL	KBCODE :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	KEY_HELD :  STD_LOGIC;
SIGNAL	KEY_INTERRUPT :  STD_LOGIC;
SIGNAL	KEYBOARD_RESPONSE :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	KEYBOARD_SCAN :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	LIGHTPEN :  STD_LOGIC;
SIGNAL	MEMORY_DATA :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	MEMORY_READY_ANTIC :  STD_LOGIC;
SIGNAL	MEMORY_READY_CPU :  STD_LOGIC;
SIGNAL	MEMORY_READY_ZPU :  STD_LOGIC;
SIGNAL	NMI_n :  STD_LOGIC;
SIGNAL	PAL :  STD_LOGIC;
SIGNAL	PAUSE_6502 :  STD_LOGIC;
SIGNAL	HALT_OR_PAUSE_6502 :  STD_LOGIC;
SIGNAL	PBI_ADDR :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	PBI_WRITE_ENABLE :  STD_LOGIC;
SIGNAL	PIA_DO :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	PIA_IRQA :  STD_LOGIC;
SIGNAL	PIA_IRQB :  STD_LOGIC;
SIGNAL	PIA_READ_ENABLE :  STD_LOGIC;
SIGNAL	PIA_WRITE_ENABLE :  STD_LOGIC;
SIGNAL	POKEY2_DO :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	CACHE_POKEY2_DO :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	POKEY2_WRITE_ENABLE :  STD_LOGIC;
SIGNAL	POKEY_DO :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	CACHE_POKEY_DO :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	POKEY_ENABLE_179 :  STD_LOGIC;
SIGNAL	POKEY_IRQ :  STD_LOGIC;
SIGNAL	POKEY_WRITE_ENABLE :  STD_LOGIC;
SIGNAL	PORTA_OUT :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	PORTA_DIR_OUT :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	PORTB_OUT :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	PORTB_DIR_OUT :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	POT_IN :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	POT_RESET :  STD_LOGIC;
SIGNAL	R_W_N :  STD_LOGIC;
SIGNAL	RAM_ADDR :  STD_LOGIC_VECTOR(18 DOWNTO 0);
SIGNAL	RAM_DO :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	RAM_REQUEST :  STD_LOGIC;
SIGNAL	RAM_REQUEST_COMPLETE :  STD_LOGIC;
SIGNAL	RAM_SELECT_dummy :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	RAM_WRITE_ENABLE :  STD_LOGIC;
SIGNAL	RESET_N :  STD_LOGIC;
SIGNAL	ROM_ADDR :  STD_LOGIC_VECTOR(21 DOWNTO 0);
SIGNAL	ROM_DO :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	ROM_REQUEST :  STD_LOGIC;
SIGNAL	ROM_REQUEST_COMPLETE :  STD_LOGIC;
SIGNAL	ROM_SELECT_dummy :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	SCANDOUBLER_SHARED_ENABLE_HIGH :  STD_LOGIC;
SIGNAL	SCANDOUBLER_SHARED_ENABLE_LOW :  STD_LOGIC;
SIGNAL	SDRAM_REFRESH :  STD_LOGIC;
--SIGNAL	SDRAM_REPLY :  STD_LOGIC;
SIGNAL	SHIFT_PRESSED :  STD_LOGIC;
SIGNAL	SIO_COMMAND_OUT :  STD_LOGIC;
SIGNAL	SIO_DATA_IN :  STD_LOGIC;
SIGNAL	SIO_DATA_OUT :  STD_LOGIC;
SIGNAL	SYNC_KEYS :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNC_SWITCHES :  STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL	SYSTEM_RESET_REQUEST :  STD_LOGIC;
SIGNAL	THROTTLE_COUNT_6502 :  STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL	TRIGGERS :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	USE_SDRAM :  STD_LOGIC;
SIGNAL	VGA :  STD_LOGIC;
SIGNAL	VIRTUAL_STICKS :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	VIRTUAL_TRIGGERS :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	VIRTUAL_KEYS :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	WIDTH_16BIT_ACCESS :  STD_LOGIC;
SIGNAL	WIDTH_32BIT_ACCESS :  STD_LOGIC;
SIGNAL	WIDTH_8BIT_ACCESS :  STD_LOGIC;
SIGNAL	WRITE_DATA :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	ZPU_16BIT_WRITE_ENABLE :  STD_LOGIC;
SIGNAL	ZPU_32BIT_WRITE_ENABLE :  STD_LOGIC;
SIGNAL	ZPU_8BIT_WRITE_ENABLE :  STD_LOGIC;
SIGNAL	ZPU_ADDR_FETCH :  STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL	ZPU_ADDR_ROM_RAM :  STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL	ZPU_CONFIG_DO :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	ZPU_CONFIG_WRITE_ENABLE :  STD_LOGIC;
SIGNAL	ZPU_DO :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	ZPU_FETCH :  STD_LOGIC;
SIGNAL	ZPU_HEX :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	ZPU_PAUSE :  STD_LOGIC;
SIGNAL	ZPU_RAM_DATA :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	ZPU_READ_ENABLE :  STD_LOGIC;
SIGNAL	ZPU_RESET :  STD_LOGIC;
SIGNAL	ZPU_ROM_DATA :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	ZPU_SECTOR_DATA :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	ZPU_STACK_WRITE :  STD_LOGIC_VECTOR(3 DOWNTO 0);

SIGNAL	LEDR_dummy :  STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL	LEDG_dummy :  STD_LOGIC_VECTOR(7 DOWNTO 0);
signal UART_TXD_dummy : std_logic;

SIGNAL		SD_DAT0 :  STD_LOGIC;
SIGNAL		SD_CLK :  STD_LOGIC;
SIGNAL		SD_CMD :  STD_LOGIC;
SIGNAL		SD_DAT3 :  STD_LOGIC;

signal mist_buttons : std_logic_vector(1 downto 0);
signal mist_switches : std_logic_vector(1 downto 0);

SIGNAL	SHIFT_PRESSED_DUMMY :  STD_LOGIC;
SIGNAL	BREAK_PRESSED_DUMMY :  STD_LOGIC;
SIGNAL	CONTROL_PRESSED :  STD_LOGIC;

signal dummy_sector_request : std_logic;
signal dummy_sector : std_logic_vector(31 downto 0);

signal COLOUR : std_logic_vector(7 downto 0);

signal POKEY1_CHANNEL0 : std_logic_vector(3 downto 0);
signal POKEY1_CHANNEL1 : std_logic_vector(3 downto 0);
signal POKEY1_CHANNEL2 : std_logic_vector(3 downto 0);
signal POKEY1_CHANNEL3 : std_logic_vector(3 downto 0);

signal POKEY2_CHANNEL0 : std_logic_vector(3 downto 0);
signal POKEY2_CHANNEL1 : std_logic_vector(3 downto 0);
signal POKEY2_CHANNEL2 : std_logic_vector(3 downto 0);
signal POKEY2_CHANNEL3 : std_logic_vector(3 downto 0);

signal hcount_temp : std_logic_vector(7 downto 0);
signal vcount_temp : std_logic_vector(8 downto 0);
signal VGA_G_dummy : std_logic_vector(7 downto 0);
signal VGA_B_dummy : std_logic_vector(7 downto 0);

signal matrix_out_match : std_logic_vector(7 downto 0);

signal keyboard_scan_inv : std_logic_vector(5 downto 0);

signal covox_write_enable : std_logic;
signal covox_channel0 : std_logic_vector(7 downto 0);
signal covox_channel1 : std_logic_vector(7 downto 0);
signal covox_channel2 : std_logic_vector(7 downto 0);
signal covox_channel3 : std_logic_vector(7 downto 0);

signal gtia_blank : std_logic;

BEGIN 

cpu6502 : cpu
PORT MAP(CLK => CLK,
		 RESET => CPU_6502_RESET,
		 ENABLE => RESET_N,
		 IRQ_n => IRQ_n,
		 NMI_n => NMI_n,
		 MEMORY_READY => MEMORY_READY_CPU,
		 THROTTLE => CPU_SHARED_ENABLE,
		 RDY => ANTIC_RDY,
		 DI => MEMORY_DATA(7 DOWNTO 0),
		 R_W_n => R_W_N,
		 CPU_FETCH => CPU_FETCH,
		 A => CPU_ADDR,
		 DO => CPU_DO);

LIGHTPEN <= '1';
antic1 : antic
PORT MAP(CLK => CLK,
		 WR_EN => ANTIC_WRITE_ENABLE,
		 RESET_N => RESET_N,
		 MEMORY_READY_ANTIC => MEMORY_READY_ANTIC,
		 MEMORY_READY_CPU => MEMORY_READY_CPU,
		 ANTIC_ENABLE_179 => ANTIC_ENABLE_179,
		 PAL => PAL,
		 lightpen => LIGHTPEN,
		 ADDR => PBI_ADDR(3 DOWNTO 0),
		 CPU_DATA_IN => WRITE_DATA(7 DOWNTO 0),
		 MEMORY_DATA_IN => MEMORY_DATA(7 DOWNTO 0),
		 NMI_N_OUT => NMI_n,
		 ANTIC_READY => ANTIC_RDY,
		 COLOUR_CLOCK_ORIGINAL_OUT => ANTIC_ORIGINAL_COLOUR_CLOCK_OUT,
		 COLOUR_CLOCK_OUT => ANTIC_COLOUR_CLOCK_OUT,
		 HIGHRES_COLOUR_CLOCK_OUT => ANTIC_HIGHRES_COLOUR_CLOCK_OUT,
		 dma_fetch_out => ANTIC_FETCH,
		 hcount_out => hcount_temp,
		 vcount_out => vcount_temp,
		 refresh_out => ANTIC_REFRESH,
		 AN => ANTIC_AN,
		 DATA_OUT => ANTIC_DO,
		 dma_address_out => ANTIC_ADDR);

pokey_mixer_l : pokey_mixer
PORT MAP(CLK => CLK,
		 GTIA_SOUND => GTIA_SOUND,
		 CHANNEL_0 => POKEY1_CHANNEL0,
		 CHANNEL_1 => POKEY1_CHANNEL1,
		 CHANNEL_2 => POKEY1_CHANNEL2,
		 CHANNEL_3 => POKEY1_CHANNEL3,
		 CHANNEL_ENABLE => "1111",
		 COVOX_CHANNEL_0 => covox_channel0,
		 COVOX_CHANNEL_1 => covox_channel1,
		 VOLUME_OUT => AUDIO_L);
		 
zpu_glue1 : zpu_glue
PORT MAP(CLK => CLK,
		 RESET => ZPU_RESET,
		 PAUSE => ZPU_PAUSE,
		 MEMORY_READY => MEMORY_READY_ZPU,
		 ZPU_CONFIG_DI => ZPU_CONFIG_DO,
		 ZPU_DI => MEMORY_DATA,
		 ZPU_RAM_DI => ZPU_RAM_DATA,
		 ZPU_ROM_DI => ZPU_ROM_DATA,
		 ZPU_SECTOR_DI => zpu_sector_data,
		 MEMORY_FETCH => ZPU_FETCH,
		 ZPU_READ_ENABLE => ZPU_READ_ENABLE,
		 ZPU_32BIT_WRITE_ENABLE => ZPU_32BIT_WRITE_ENABLE,
		 ZPU_16BIT_WRITE_ENABLE => ZPU_16BIT_WRITE_ENABLE,
		 ZPU_8BIT_WRITE_ENABLE => ZPU_8BIT_WRITE_ENABLE,
		 ZPU_CONFIG_WRITE => ZPU_CONFIG_WRITE_ENABLE,
		 ZPU_ADDR_FETCH => ZPU_ADDR_FETCH,
		 ZPU_ADDR_ROM_RAM => ZPU_ADDR_ROM_RAM,
		 ZPU_DO => ZPU_DO,
		 ZPU_STACK_WRITE => ZPU_STACK_WRITE);


pokey_mixer_r : pokey_mixer
PORT MAP(CLK => CLK,
		 GTIA_SOUND => GTIA_SOUND,
		 CHANNEL_0 => POKEY2_CHANNEL0,
		 CHANNEL_1 => POKEY2_CHANNEL1,
		 CHANNEL_2 => POKEY2_CHANNEL2,
		 CHANNEL_3 => POKEY2_CHANNEL3,
		 COVOX_CHANNEL_0 => covox_channel2,
		 COVOX_CHANNEL_1 => covox_channel3,
		 CHANNEL_ENABLE => "1111",
		 VOLUME_OUT => AUDIO_R);


pokey2 : pokey
PORT MAP(CLK => CLK,
		 CPU_MEMORY_READY => MEMORY_READY_CPU,
		 ANTIC_MEMORY_READY => MEMORY_READY_ANTIC,
		 WR_EN => POKEY2_WRITE_ENABLE,
		 RESET_N => RESET_N,
		 ADDR => PBI_ADDR(3 DOWNTO 0),
		 DATA_IN => WRITE_DATA(7 DOWNTO 0),
		 CHANNEL_0_OUT => POKEY2_CHANNEL0,
		 CHANNEL_1_OUT => POKEY2_CHANNEL1,
		 CHANNEL_2_OUT => POKEY2_CHANNEL2,
		 CHANNEL_3_OUT => POKEY2_CHANNEL3,
		 DATA_OUT => POKEY2_DO,
		 SIO_IN1 => '1',
		 SIO_IN2 => '1',
		 SIO_IN3 => '1',
		 keyboard_response => "00",
		 pot_in=>"00000000");


-- PIA
--GPIO_0[0] <= CA2_OUT when CA2_DIR_OUT='1' else 'Z';
--CA2_IN <= GPIO_0[0];

--GPIO_O[1] <= CB2_OUT when CB2_DIR_OUT='1' else 'Z';
--CB2_IN <= GPIO_O[1];
SIO_COMMAND_OUT <= CB2_OUT; -- we generate command frame, use internal rather than from pin
SIO_COMMAND_TX <= SIO_COMMAND_OUT;
-- TODO - sioto gpio!
GPIO_PORTB_IN <= PORTB_OUT;
GPIO_CA2_IN <= CA2_OUT when CA2_DIR_OUT='1' else '1';
GPIO_CB2_IN <= CB2_OUT when CB2_DIR_OUT='1' else '1';
GPIO_PORTA_IN <= ((JOY1_n(3)&JOY1_n(2)&JOY1_n(1)&JOY1_n(0)&JOY2_n(3)&JOY2_n(2)&JOY2_n(1)&JOY2_n(0)) and not (porta_dir_out)) or (porta_dir_out and porta_out);

pia1 : pia
PORT MAP(CLK => CLK,
		 EN => PIA_READ_ENABLE,
		 WR_EN => PIA_WRITE_ENABLE,
		 RESET_N => RESET_N,
		 CA1 => '1', --todo - high/low?
		 CB1 => '1',
		 CA2_DIR_OUT => CA2_DIR_OUT,
		 CA2_IN => GPIO_CA2_IN,
		 CA2_OUT => CA2_OUT,
		 CB2_DIR_OUT => CB2_DIR_OUT,
		 CB2_IN => GPIO_CB2_IN,
		 CB2_OUT => CB2_OUT,
		 ADDR => PBI_ADDR(1 DOWNTO 0),
		 CPU_DATA_IN => WRITE_DATA(7 DOWNTO 0),
		 IRQA_N => PIA_IRQA,
		 IRQB_N => PIA_IRQB,
		 DATA_OUT => PIA_DO,
		 PORTA_IN => GPIO_PORTA_IN,
		 PORTA_DIR_OUT => PORTA_DIR_OUT,
		 PORTA_OUT => PORTA_OUT,
		 PORTB_IN => GPIO_PORTB_IN,
		 PORTB_DIR_OUT => PORTB_DIR_OUT,
		 PORTB_OUT => PORTB_OUT);

HALT_OR_PAUSE_6502 <= HALT or PAUSE_6502;
enables : shared_enable
PORT MAP(CLK => CLK,
		 RESET_N => RESET_N,
		 MEMORY_READY_CPU => MEMORY_READY_CPU,
		 MEMORY_READY_ANTIC => MEMORY_READY_ANTIC,
		 PAUSE_6502 => HALT_OR_PAUSE_6502,
		 THROTTLE_COUNT_6502 => THROTTLE_COUNT_6502,
		 POKEY_ENABLE_179 => POKEY_ENABLE_179,
		 ANTIC_ENABLE_179 => ANTIC_ENABLE_179,
		 oldcpu_enable => ENABLE_179_MEMWAIT,
		 CPU_ENABLE_OUT => CPU_SHARED_ENABLE,
		 SCANDOUBLER_ENABLE_LOW => SCANDOUBLER_SHARED_ENABLE_LOW,
		 SCANDOUBLER_ENABLE_HIGH => SCANDOUBLER_SHARED_ENABLE_HIGH);

-- no cart!
CART_RD4 <= '0';
CART_RD5 <= '0';
CART_REQUEST_COMPLETE <= '0';
CART_ROM_DO <= (others=>'0');

mmu1 : address_decoder
PORT MAP(CLK => CLK,
		 CPU_FETCH => CPU_FETCH,
		 CPU_WRITE_N => R_W_N,
		 ANTIC_FETCH => ANTIC_FETCH,
		 antic_refresh => ANTIC_REFRESH,
		 ZPU_FETCH => ZPU_FETCH,
		 ZPU_READ_ENABLE => ZPU_READ_ENABLE,
		 ZPU_32BIT_WRITE_ENABLE => ZPU_32BIT_WRITE_ENABLE,
		 ZPU_16BIT_WRITE_ENABLE => ZPU_16BIT_WRITE_ENABLE,
		 ZPU_8BIT_WRITE_ENABLE => ZPU_8BIT_WRITE_ENABLE,
		 RAM_REQUEST_COMPLETE => RAM_REQUEST_COMPLETE,
		 ROM_REQUEST_COMPLETE => ROM_REQUEST_COMPLETE,
		 CART_REQUEST_COMPLETE => CART_REQUEST_COMPLETE,
		 reset_n => RESET_N,
		 CART_RD4 => CART_RD4,
		 CART_RD5 => CART_RD5,
		 use_sdram => USE_SDRAM,
		 SDRAM_REQUEST_COMPLETE => SDRAM_REQUEST_COMPLETE,
		 ANTIC_ADDR => ANTIC_ADDR,
		 ANTIC_DATA => ANTIC_DO,
		 CACHE_ANTIC_DATA => CACHE_ANTIC_DO,
		 CART_ROM_DATA => CART_ROM_DO,
		 CPU_ADDR => CPU_ADDR,
		 CPU_WRITE_DATA => CPU_DO,
		 GTIA_DATA => GTIA_DO,
		 CACHE_GTIA_DATA => CACHE_GTIA_DO,
		 PIA_DATA => PIA_DO,
		 POKEY2_DATA => POKEY2_DO,
		 CACHE_POKEY2_DATA => CACHE_POKEY2_DO,
		 POKEY_DATA => POKEY_DO,
		 CACHE_POKEY_DATA => CACHE_POKEY_DO,
		 PORTB => PORTB_OUT,
		 RAM_DATA => RAM_DO,
		 ram_select => RAM_SELECT(2 downto 0),
		 ROM_DATA => ROM_DO,
		 rom_select => ROM_SELECT, 
		 SDRAM_DATA => SDRAM_DO,
		 ZPU_ADDR => ZPU_ADDR_FETCH,
		 ZPU_WRITE_DATA => ZPU_DO,
		 MEMORY_READY_ANTIC => MEMORY_READY_ANTIC,
		 MEMORY_READY_ZPU => MEMORY_READY_ZPU,
		 MEMORY_READY_CPU => MEMORY_READY_CPU,
		 GTIA_WR_ENABLE => GTIA_WRITE_ENABLE,
		 POKEY_WR_ENABLE => POKEY_WRITE_ENABLE,
		 POKEY2_WR_ENABLE => POKEY2_WRITE_ENABLE,
		 ANTIC_WR_ENABLE => ANTIC_WRITE_ENABLE,
		 PIA_WR_ENABLE => PIA_WRITE_ENABLE,
		 PIA_RD_ENABLE => PIA_READ_ENABLE,
		 RAM_WR_ENABLE => RAM_WRITE_ENABLE,
		 PBI_WR_ENABLE => PBI_WRITE_ENABLE,
		 RAM_REQUEST => RAM_REQUEST,
		 ROM_REQUEST => ROM_REQUEST,
		 CART_REQUEST => CART_REQUEST,
		 CART_S4_n => CART_S4_n,
		 CART_S5_n => CART_S5_N,
		 CART_CCTL_n => CART_CCTL_N,
		 WIDTH_8bit_ACCESS => WIDTH_8BIT_ACCESS,
		 WIDTH_16bit_ACCESS => WIDTH_16BIT_ACCESS,
		 WIDTH_32bit_ACCESS => WIDTH_32BIT_ACCESS,
		 SDRAM_READ_EN => SDRAM_READ_ENABLE,
		 SDRAM_WRITE_EN => SDRAM_WRITE_ENABLE,
		 SDRAM_REQUEST => SDRAM_REQUEST,
		 SDRAM_REFRESH => SDRAM_REFRESH,
		 MEMORY_DATA => MEMORY_DATA,
		 PBI_ADDR => PBI_ADDR,
		 RAM_ADDR => RAM_ADDR,
		 ROM_ADDR => ROM_ADDR,
		 SDRAM_ADDR => SDRAM_ADDR,
		 WRITE_DATA => WRITE_DATA,
		 d6_wr_enable => covox_write_enable,
		 cart_select => "0000000",
		 cart_activate => '0');

zpu_rom1 : zpu_rom
PORT MAP(clock => CLK,
		 address => ZPU_ADDR_ROM_RAM(13 DOWNTO 2),
		 q => ZPU_ROM_DATA);
--
--b2v_inst23 : zpu_ram
--PORT MAP(wren => ZPU_STACK_WRITE(2),
--		 clock => CLK,
--		 address => ZPU_ADDR_ROM_RAM(11 DOWNTO 2),
--		 data => ZPU_DO(23 DOWNTO 16),
--		 q => ZPU_RAM_DATA(23 DOWNTO 16));

zpu_ram1 : generic_ram_infer
generic map
(
	ADDRESS_WIDTH => 10,
	SPACE => 1024,
	DATA_WIDTH =>8
)
PORT MAP(clock => clk,
		 address => ZPU_ADDR_ROM_RAM(11 downto 2),
		 data => ZPU_DO(23 downto 16),
		 we => ZPU_STACK_WRITE(2),
		 q => ZPU_RAM_DATA(23 downto 16)
		 );	

SYNC_KEYS <= (others=> '0');
SYNC_SWITCHES <= (others=> '1');
zpu_config1 : zpu_config_regs
PORT MAP(CLK => CLK,
		 ENABLE_179 => POKEY_ENABLE_179,
		 WR_EN => ZPU_CONFIG_WRITE_ENABLE,
		 SDCARD_DAT => SD_DAT0,
		 SIO_COMMAND_OUT => SIO_COMMAND_OUT,
		 SIO_DATA_OUT => SIO_DATA_OUT,
		 PLL_LOCKED => PLL_LOCKED,
		 REQUEST_RESET_ZPU => SYSTEM_RESET_REQUEST,
		 ADDR => ZPU_ADDR_ROM_RAM(6 DOWNTO 2),
		 CPU_DATA_IN => ZPU_DO,
		 KEY => VIRTUAL_KEYS, --SYNC_KEYS,
		 SWITCH => SYNC_SWITCHES,
		 SDCARD_CLK => SD_CLK,
		 SDCARD_CMD => SD_CMD,
		 SDCARD_DAT3 => SD_DAT3,
		 SIO_DATA_IN => SIO_DATA_IN,
		 PAUSE_ZPU => ZPU_PAUSE,
		 PAL => PAL,
		 USE_SDRAM => USE_SDRAM,
		 VGA => VGA,
		 COMPOSITE_ON_HSYNC => COMPOSITE_ON_HSYNC,
		 GPIO_ENABLE => GPIO_ENABLE,
		 RESET_6502 => CPU_6502_RESET,
		 RESET_ZPU => ZPU_RESET,
		 RESET_N => RESET_N,
		 PAUSE_6502 => PAUSE_6502,
		 DATA_OUT => ZPU_CONFIG_DO,
		 LEDG => LEDG_dummy,
		 LEDR => LEDR_dummy,
		 RAM_SELECT => RAM_SELECT_dummy,
		 ROM_SELECT => ROM_SELECT_dummy(1 downto 0),
		 THROTTLE_COUNT_6502 => THROTTLE_COUNT_6502,
		 ZPU_HEX => ZPU_HEX,
		 sector_request => dummy_sector_request,
		 sector => dummy_sector,
		 sector_ready => '0'
		 );
ROM_SELECT_dummy(5 downto 2) <= "0000";

--
--b2v_inst25 : zpu_ram
--PORT MAP(wren => ZPU_STACK_WRITE(3),
--		 clock => CLK,
--		 address => ZPU_ADDR_ROM_RAM(11 DOWNTO 2),
--		 data => ZPU_DO(31 DOWNTO 24),
--		 q => ZPU_RAM_DATA(31 DOWNTO 24));

zpu_ram2 : generic_ram_infer
generic map
(
	ADDRESS_WIDTH => 10,
	SPACE => 1024,
	DATA_WIDTH =>8
)
PORT MAP(clock => clk,
		 address => ZPU_ADDR_ROM_RAM(11 downto 2),
		 data => ZPU_DO(31 downto 24),
		 we => ZPU_STACK_WRITE(3),
		 q => ZPU_RAM_DATA(31 downto 24)
		 );	


--b2v_inst26 : zpu_ram
--PORT MAP(wren => ZPU_STACK_WRITE(0),
--		 clock => CLK,
--		 address => ZPU_ADDR_ROM_RAM(11 DOWNTO 2),
--		 data => ZPU_DO(7 DOWNTO 0),
--		 q => ZPU_RAM_DATA(7 DOWNTO 0));

zpu_ram3 : generic_ram_infer
generic map
(
	ADDRESS_WIDTH => 10,
	SPACE => 1024,
	DATA_WIDTH =>8
)
PORT MAP(clock => clk,
		 address => ZPU_ADDR_ROM_RAM(11 downto 2),
		 data => ZPU_DO(7 downto 0),
		 we => ZPU_STACK_WRITE(0),
		 q => ZPU_RAM_DATA(7 downto 0)
		 );	


--b2v_inst27 : zpu_ram
--PORT MAP(wren => ZPU_STACK_WRITE(1),
--		 clock => CLK,
--		 address => ZPU_ADDR_ROM_RAM(11 DOWNTO 2),
--		 data => ZPU_DO(15 DOWNTO 8),
--		 q => ZPU_RAM_DATA(15 DOWNTO 8));

zpu_ram4 : generic_ram_infer
generic map
(
	ADDRESS_WIDTH => 10,
	SPACE => 1024,
	DATA_WIDTH =>8
)
PORT MAP(clock => clk,
		 address => ZPU_ADDR_ROM_RAM(11 downto 2),
		 data => ZPU_DO(15 downto 8),
		 we => ZPU_STACK_WRITE(1),
		 q => ZPU_RAM_DATA(15 downto 8)
		 );	

pokey1 : pokey
PORT MAP(CLK => CLK,
		 CPU_MEMORY_READY => MEMORY_READY_CPU,
		 ANTIC_MEMORY_READY => MEMORY_READY_ANTIC,
		 WR_EN => POKEY_WRITE_ENABLE,
		 RESET_N => RESET_N,
		 SIO_IN1 => SIO_RXD,
		 SIO_IN2 => '1',
		 SIO_IN3 => SIO_DATA_IN,
		 ADDR => PBI_ADDR(3 DOWNTO 0),
		 DATA_IN => WRITE_DATA(7 DOWNTO 0),
		 keyboard_response => KEYBOARD_RESPONSE,
		 POT_IN => POT_IN,
		 IRQ_N_OUT => POKEY_IRQ,
		 SIO_OUT1 => SIO_TXD,
		 SIO_OUT2 => GPIO_SIO_OUT,
		 SIO_OUT3 => SIO_DATA_OUT,
		 POT_RESET => POT_RESET,
		 CHANNEL_0_OUT => POKEY1_CHANNEL0,
		 CHANNEL_1_OUT => POKEY1_CHANNEL1,
		 CHANNEL_2_OUT => POKEY1_CHANNEL2,
		 CHANNEL_3_OUT => POKEY1_CHANNEL3,
		 DATA_OUT => POKEY_DO,
		 keyboard_scan => KEYBOARD_SCAN);

	keyboard_scan_inv <= not(keyboard_scan);

a4051: complete_address_decoder
	generic map (width => 3)
	PORT map ( addr_in => keyboard_scan_inv(5 downto 3), addr_decoded => matrix_in ); 

b4051: complete_address_decoder
	generic map (width => 3)
	PORT map ( addr_in => keyboard_scan_inv(2 downto 0), addr_decoded => matrix_out_match ); 

	process(matrix_out, matrix_out_match)
	begin
		keyboard_response(0) <= '1';

		if (or_reduce(matrix_out(7 downto 0) and matrix_out_match(7 downto 0)) = '1') then
			keyboard_response(0) <= '0';
		end if;
	end process;

	process(static_keys, pause_key)
	begin
		keyboard_response(1) <= '1';

		if (keyboard_scan(5 downto 4)="00" and pause_key = '1') then
			keyboard_response(1) <= '0';
		end if;
		
		if (keyboard_scan(5 downto 4)="10" and static_keys(0) = '1') then
			keyboard_response(1) <= '0';
		end if;

		if (keyboard_scan(5 downto 4)="11" and static_keys(1) = '1') then
			keyboard_response(1) <= '0';
		end if;
	end process;

	CONSOL_START <= static_keys(6);
	CONSOL_SELECT <= static_keys(5);
	CONSOL_OPTION <= static_keys(4);
	system_reset_request <= static_keys(3);

	virtual_keys <= "000"&static_keys(2); -- todo need more static keys!! though on second thoughts using replay menu for options/loading...
	virtual_triggers <= "00"&joy1_n(4)&joy2_n(4); -- todo joystick...
		 	 
gtia1 : gtia
PORT MAP(CLK => CLK,
		 WR_EN => GTIA_WRITE_ENABLE,
		 CPU_MEMORY_READY => MEMORY_READY_CPU,
		 ANTIC_MEMORY_READY => MEMORY_READY_ANTIC,
		 ANTIC_FETCH => ANTIC_FETCH,
		 CPU_ENABLE_ORIGINAL => ENABLE_179_MEMWAIT,
		 RESET_N => RESET_N,
		 PAL => PAL,
		 COLOUR_CLOCK_ORIGINAL => ANTIC_ORIGINAL_COLOUR_CLOCK_OUT,
		 COLOUR_CLOCK => ANTIC_COLOUR_CLOCK_OUT,
		 COLOUR_CLOCK_HIGHRES => ANTIC_HIGHRES_COLOUR_CLOCK_OUT,
		 CONSOL_START => CONSOL_START,
		 CONSOL_SELECT => CONSOL_SELECT,
		 CONSOL_OPTION => CONSOL_OPTION,
		 TRIG0 => joy2_n(4), -- TODO - joystick trigger too
		 TRIG1 => joy1_n(4),
		 --TRIG0 => VIRTUAL_TRIGGERS(0) and joy2_n(4), -- TODO - joystick trigger too
		 --TRIG1 => VIRTUAL_TRIGGERS(1) and joy1_n(4),
		 --TRIG0 => VIRTUAL_TRIGGERS(0),
		 --TRIG1 => VIRTUAL_TRIGGERS(1),
		 TRIG2 => VIRTUAL_TRIGGERS(2),
		 TRIG3 => VIRTUAL_TRIGGERS(3),
		 ADDR => PBI_ADDR(4 DOWNTO 0),
		 AN => ANTIC_AN,
		 CPU_DATA_IN => WRITE_DATA(7 DOWNTO 0),
		 MEMORY_DATA_IN => MEMORY_DATA(7 DOWNTO 0),
		 VSYNC => VGA_VS,
		 HSYNC => VGA_HS,
		 BLANK => GTIA_BLANK,
		 sound => GTIA_SOUND,
		 COLOUR_out => COLOUR,
		 DATA_OUT => GTIA_DO);

	-- colour palette
--	Color             Value         Color             Value
--Black           0,      0	Medium blue     8,    128
--Rust            1,     16       Dark blue       9,    144
--Red-orange      2,     32       Blue-grey      10,    160
--Dark orange     3,     48       Olive green    11,    176
--Red             4,     64       Medium green   12,    192
--Dk lavender     5,     80       Dark green     13,    208
--Cobalt blue     6,     96       Orange-green   14,    224
--Ultramarine     7,    112       Orange         15,    240

-- from altirra	
	palette1 : entity work.gtia_palette(altirra)
		port map (ATARI_COLOUR=>COLOUR, R_next=>VGA_R, G_next=>VGA_G, B_next=>VGA_B);
	--VGA_B <= hcount_temp;
	--VGA_G <= vcount_temp(7 downto 0);
		
-- from lao
--	palette2 : entity work.gtia_palette(laoo)
--		port map (ATARI_COLOUR=>COLOUR, R_next=>R_next, G_next=>G_next, B_next=>B_next);		


irq_glue1 : irq_glue
PORT MAP(pokey_irq => POKEY_IRQ,
		 pia_irqa => PIA_IRQA,
		 pia_irqb => PIA_IRQB,
		 combined_irq => IRQ_n);
		 
pokey1_mirror : reg_file
generic map(BYTES=>16,WIDTH=>4)
port map(
	CLK => CLK,
	ADDR => PBI_ADDR(3 downto 0),
	DATA_IN => WRITE_DATA(7 downto 0),
	WR_EN => POKEY_WRITE_ENABLE,
	DATA_OUT => CACHE_POKEY_DO
);	 

pokey2_mirror : reg_file
generic map(BYTES=>16,WIDTH=>4)
port map(
	CLK => CLK,
	ADDR => PBI_ADDR(3 downto 0),
	DATA_IN => WRITE_DATA(7 downto 0),
	WR_EN => POKEY2_WRITE_ENABLE,
	DATA_OUT => CACHE_POKEY2_DO
);	 		 

gtia_mirror : reg_file
generic map(BYTES=>32,WIDTH=>5)
port map(
	CLK => CLK,
	ADDR => PBI_ADDR(4 downto 0),
	DATA_IN => WRITE_DATA(7 downto 0),
	WR_EN => GTIA_WRITE_ENABLE,
	DATA_OUT => CACHE_GTIA_DO
);	

antic_mirror : reg_file
generic map(BYTES=>16,WIDTH=>4)
port map(
	CLK => CLK,
	ADDR => PBI_ADDR(3 downto 0),
	DATA_IN => WRITE_DATA(7 downto 0),
	WR_EN => ANTIC_WRITE_ENABLE,
	DATA_OUT => CACHE_ANTIC_DO
);	

internalromram1 : internalromram
  PORT map(
    clock => clk,
    reset_n => reset_n,

	ROM_ADDR =>rom_addr,
	ROM_REQUEST_COMPLETE => rom_REQUEST_COMPLETE,
	ROM_REQUEST => rom_REQUEST,
	ROM_DATA => rom_DO,
	
	RAM_ADDR => ram_addr,
	RAM_WR_ENABLE => ram_WRITE_ENABLE,
	RAM_DATA_IN => wriTE_DATA(7 downto 0),
	RAM_REQUEST_COMPLETE => ram_REQUEST_COMPLETE,
	RAM_REQUEST => ram_REQUEST,
	RAM_DATA => ram_do(7 downto 0)
	);

SDRAM_WIDTH_8bit_ACCESS <= WIDTH_8bit_access;
SDRAM_WIDTH_16bit_ACCESS <= WIDTH_16bit_access;
SDRAM_WIDTH_32bit_ACCESS <= WIDTH_32bit_access;
SDRAM_DI <= WRITE_DATA;

covox1 : covox
	PORT map
	( 
		clk => clk,
		addr => pbi_addr(1 downto 0),
		data_in => WRITE_DATA(7 DOWNTO 0),
		wr_en => covox_write_enable,
		covox_channel0 => covox_channel0,
		covox_channel1 => covox_channel1,
		covox_channel2 => covox_channel2,
		covox_channel3 => covox_channel3
	);

END bdf_type;
