
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f6",
X"80738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80fa",
X"a00c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f3",
X"ad2d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580f2ec",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80dcfb04",
X"fd3d0d75",
X"705254ae",
X"aa3f83e0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83e0",
X"8008732e",
X"a13883e0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183e0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83e2c008",
X"248a38b4",
X"fb3fff0b",
X"83e2c00c",
X"800b83e0",
X"800c04ff",
X"3d0d7352",
X"83e09c08",
X"722e8d38",
X"d93f7151",
X"96a03f71",
X"83e09c0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"55805681",
X"54bc1508",
X"762e0981",
X"06819138",
X"7451c83f",
X"7958757a",
X"2580f738",
X"83e2f008",
X"70892a57",
X"83ff0678",
X"84807231",
X"56565773",
X"78258338",
X"73557583",
X"e2c0082e",
X"8438ff82",
X"3f83e2c0",
X"088025a6",
X"3875892b",
X"5198dc3f",
X"83e2f008",
X"8f3dfc11",
X"555c5481",
X"52f81b51",
X"96c63f76",
X"1483e2f0",
X"0c7583e2",
X"c00c7453",
X"76527851",
X"b3a53f83",
X"e0800883",
X"e2f00816",
X"83e2f00c",
X"78763176",
X"1b5b5956",
X"778024ff",
X"8b38617a",
X"710c5475",
X"5475802e",
X"83388154",
X"7383e080",
X"0c8e3d0d",
X"04fc3d0d",
X"fe943f76",
X"51fea83f",
X"863dfc05",
X"53785277",
X"5195e93f",
X"7975710c",
X"5483e080",
X"085483e0",
X"8008802e",
X"83388154",
X"7383e080",
X"0c863d0d",
X"04fe3d0d",
X"7583e2c0",
X"08535380",
X"72248938",
X"71732e84",
X"38fdcf3f",
X"7451fde3",
X"3f725197",
X"ae3f83e0",
X"80085283",
X"e0800880",
X"2e833881",
X"527183e0",
X"800c843d",
X"0d04803d",
X"0d7280c0",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d72bc",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"c40b83e0",
X"800c04fd",
X"3d0d7577",
X"71547053",
X"5553a9fb",
X"3f82c813",
X"08bc150c",
X"82c01308",
X"80c0150c",
X"fce43f73",
X"5193ab3f",
X"7383e09c",
X"0c83e080",
X"085383e0",
X"8008802e",
X"83388153",
X"7283e080",
X"0c853d0d",
X"04fd3d0d",
X"75775553",
X"fcb83f72",
X"802ea538",
X"bc130852",
X"7351a985",
X"3f83e080",
X"088f3877",
X"527251ff",
X"9a3f83e0",
X"8008538a",
X"3982cc13",
X"0853d839",
X"81537283",
X"e0800c85",
X"3d0d04fe",
X"3d0dff0b",
X"83e2c00c",
X"7483e0a0",
X"0c7583e2",
X"bc0cafd9",
X"3f83e080",
X"0881ff06",
X"52815371",
X"993883e2",
X"d8518e94",
X"3f83e080",
X"085283e0",
X"8008802e",
X"83387252",
X"71537283",
X"e0800c84",
X"3d0d04fa",
X"3d0d787a",
X"82c41208",
X"82c41208",
X"70722459",
X"56565757",
X"73732e09",
X"81069138",
X"80c01652",
X"80c01751",
X"a6f63f83",
X"e0800855",
X"7483e080",
X"0c883d0d",
X"04f63d0d",
X"7c5b807b",
X"715c5457",
X"7a772e8c",
X"38811a82",
X"cc140854",
X"5a72f638",
X"805980d9",
X"397a5481",
X"5780707b",
X"7b315a57",
X"55ff1853",
X"74732580",
X"c13882cc",
X"14085273",
X"51ff8c3f",
X"800b83e0",
X"800825a1",
X"3882cc14",
X"0882cc11",
X"0882cc16",
X"0c7482cc",
X"120c5375",
X"802e8638",
X"7282cc17",
X"0c725480",
X"577382cc",
X"15088117",
X"575556ff",
X"b8398119",
X"59800bff",
X"1b545478",
X"73258338",
X"81547681",
X"32707506",
X"515372ff",
X"90388c3d",
X"0d04f73d",
X"0d7b7d5a",
X"5a82d052",
X"83e2bc08",
X"5180e1e8",
X"3f83e080",
X"0857f9da",
X"3f795283",
X"e2c45195",
X"b73f83e0",
X"80085480",
X"5383e080",
X"08732e09",
X"81068283",
X"3883e0a0",
X"080b0b80",
X"f7b85370",
X"5256a6b3",
X"3f0b0b80",
X"f7b85280",
X"c01651a6",
X"a63f75bc",
X"170c7382",
X"c0170c81",
X"0b82c417",
X"0c810b82",
X"c8170c73",
X"82cc170c",
X"ff1782d0",
X"17555781",
X"913983e0",
X"ac337082",
X"2a708106",
X"51545572",
X"81803874",
X"812a8106",
X"587780f6",
X"3874842a",
X"810682c4",
X"150c83e0",
X"ac338106",
X"82c8150c",
X"79527351",
X"a5cd3f73",
X"51a5e43f",
X"83e08008",
X"1453af73",
X"70810555",
X"3472bc15",
X"0c83e0ad",
X"527251a5",
X"ae3f83e0",
X"a40882c0",
X"150c83e0",
X"ba5280c0",
X"1451a59b",
X"3f78802e",
X"8d387351",
X"782d83e0",
X"8008802e",
X"99387782",
X"cc150c75",
X"802e8638",
X"7382cc17",
X"0c7382d0",
X"15ff1959",
X"55567680",
X"2e9b3883",
X"e0a45283",
X"e2c45194",
X"ad3f83e0",
X"80088a38",
X"83e0ad33",
X"5372fed2",
X"3878802e",
X"893883e0",
X"a00851fc",
X"b83f83e0",
X"a0085372",
X"83e0800c",
X"8b3d0d04",
X"ff3d0d80",
X"527351fd",
X"b53f833d",
X"0d04f03d",
X"0d627052",
X"54f6893f",
X"83e08008",
X"7453873d",
X"70535555",
X"f6a93ff7",
X"893f7351",
X"d33f6353",
X"745283e0",
X"800851fa",
X"b83f923d",
X"0d047183",
X"e0800c04",
X"80c01283",
X"e0800c04",
X"803d0d72",
X"82c01108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"7282cc11",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282c4",
X"110883e0",
X"800c5182",
X"3d0d04f9",
X"3d0d7983",
X"e0900857",
X"57817727",
X"81963876",
X"88170827",
X"818e3875",
X"33557482",
X"2e893874",
X"832eb338",
X"80fe3974",
X"54761083",
X"fe065376",
X"882a8c17",
X"08055289",
X"3dfc0551",
X"aa873f83",
X"e0800880",
X"df38029d",
X"0533893d",
X"3371882b",
X"07565680",
X"d1398454",
X"76822b83",
X"fc065376",
X"872a8c17",
X"08055289",
X"3dfc0551",
X"a9d73f83",
X"e08008b0",
X"38029f05",
X"33028405",
X"9e053371",
X"982b7190",
X"2b07028c",
X"059d0533",
X"70882b72",
X"078d3d33",
X"7180ffff",
X"fe800607",
X"51525357",
X"58568339",
X"81557483",
X"e0800c89",
X"3d0d04fb",
X"3d0d83e0",
X"9008fe19",
X"881208fe",
X"05555654",
X"80567473",
X"278d3882",
X"14337571",
X"29941608",
X"05575375",
X"83e0800c",
X"873d0d04",
X"fc3d0d76",
X"52800b83",
X"e0900870",
X"33515253",
X"70832e09",
X"81069138",
X"95123394",
X"13337198",
X"2b71902b",
X"07555551",
X"9b12339a",
X"13337188",
X"2b077407",
X"83e0800c",
X"55863d0d",
X"04fc3d0d",
X"7683e090",
X"08555580",
X"75238815",
X"08537281",
X"2e883888",
X"14087326",
X"85388152",
X"b2397290",
X"38733352",
X"71832e09",
X"81068538",
X"90140853",
X"728c160c",
X"72802e8d",
X"387251fe",
X"d63f83e0",
X"80085285",
X"39901408",
X"52719016",
X"0c805271",
X"83e0800c",
X"863d0d04",
X"fa3d0d78",
X"83e09008",
X"71228105",
X"7083ffff",
X"06575457",
X"5573802e",
X"88389015",
X"08537286",
X"38835280",
X"e739738f",
X"06527180",
X"da388113",
X"90160c8c",
X"15085372",
X"9038830b",
X"84172257",
X"52737627",
X"80c638bf",
X"39821633",
X"ff057484",
X"2a065271",
X"b2387251",
X"fcb13f81",
X"527183e0",
X"800827a8",
X"38835283",
X"e0800888",
X"1708279c",
X"3883e080",
X"088c160c",
X"83e08008",
X"51fdbc3f",
X"83e08008",
X"90160c73",
X"75238052",
X"7183e080",
X"0c883d0d",
X"04f23d0d",
X"60626458",
X"5e5b7533",
X"5574a02e",
X"09810688",
X"38811670",
X"4456ef39",
X"62703356",
X"5674af2e",
X"09810684",
X"38811643",
X"800b881c",
X"0c627033",
X"5155749f",
X"2691387a",
X"51fdd23f",
X"83e08008",
X"56807d34",
X"83813993",
X"3d841c08",
X"7058595f",
X"8a55a076",
X"70810558",
X"34ff1555",
X"74ff2e09",
X"8106ef38",
X"80705a5c",
X"887f085f",
X"5a7b811d",
X"7081ff06",
X"60137033",
X"70af3270",
X"30a07327",
X"71802507",
X"5151525b",
X"535e5755",
X"7480e738",
X"76ae2e09",
X"81068338",
X"8155787a",
X"27750755",
X"74802e9f",
X"38798832",
X"703078ae",
X"32703070",
X"73079f2a",
X"53515751",
X"5675bb38",
X"88598b5a",
X"ffab3976",
X"982b5574",
X"80258738",
X"80f59017",
X"3357ff9f",
X"17557499",
X"268938e0",
X"177081ff",
X"06585578",
X"811a7081",
X"ff06721b",
X"535b5755",
X"767534fe",
X"f8397b1e",
X"7f0c8055",
X"76a02683",
X"38815574",
X"8b19347a",
X"51fc823f",
X"83e08008",
X"80f538a0",
X"547a2270",
X"852b83e0",
X"06545590",
X"1b08527c",
X"51a4923f",
X"83e08008",
X"5783e080",
X"08818138",
X"7c335574",
X"802e80f4",
X"388b1d33",
X"70832a70",
X"81065156",
X"5674b438",
X"8b7d841d",
X"0883e080",
X"08595b5b",
X"58ff1858",
X"77ff2e9a",
X"38797081",
X"055b3379",
X"7081055b",
X"33717131",
X"52565675",
X"802ee238",
X"86397580",
X"2e96387a",
X"51fbe53f",
X"ff863983",
X"e0800856",
X"83e08008",
X"b6388339",
X"7656841b",
X"088b1133",
X"515574a7",
X"388b1d33",
X"70842a70",
X"81065156",
X"56748938",
X"83569439",
X"81569039",
X"7c51fa94",
X"3f83e080",
X"08881c0c",
X"fd813975",
X"83e0800c",
X"903d0d04",
X"f83d0d7a",
X"7c595782",
X"5483fe53",
X"77527651",
X"a2d73f83",
X"5683e080",
X"0880ec38",
X"81173377",
X"3371882b",
X"07565682",
X"567482d4",
X"d52e0981",
X"0680d438",
X"7554b653",
X"77527651",
X"a2ab3f83",
X"e0800898",
X"38811733",
X"77337188",
X"2b0783e0",
X"80085256",
X"56748182",
X"c62eac38",
X"825480d2",
X"53775276",
X"51a2823f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62e83",
X"38815675",
X"83e0800c",
X"8a3d0d04",
X"eb3d0d67",
X"5a800b83",
X"e0900ca1",
X"a43f83e0",
X"80088106",
X"55825674",
X"83ef3874",
X"75538f3d",
X"70535759",
X"feca3f83",
X"e0800881",
X"ff065776",
X"812e0981",
X"0680d438",
X"905483be",
X"53745275",
X"51a1963f",
X"83e08008",
X"80c9388f",
X"3d335574",
X"802e80c9",
X"3802bf05",
X"33028405",
X"be053371",
X"982b7190",
X"2b07028c",
X"05bd0533",
X"70882b72",
X"07953d33",
X"71077058",
X"7b575e52",
X"5e575957",
X"fdee3f83",
X"e0800881",
X"ff065776",
X"832e0981",
X"06863881",
X"5682f239",
X"76802e86",
X"38865682",
X"e839a454",
X"8d537852",
X"7551a0ad",
X"3f815683",
X"e0800882",
X"d43802be",
X"05330284",
X"05bd0533",
X"71882b07",
X"595d77ab",
X"380280ce",
X"05330284",
X"0580cd05",
X"3371982b",
X"71902b07",
X"973d3370",
X"882b7207",
X"02940580",
X"cb053371",
X"0754525e",
X"57595602",
X"b7053378",
X"71290288",
X"05b60533",
X"028c05b5",
X"05337188",
X"2b07701d",
X"707f8c05",
X"0c5f5957",
X"595d8e3d",
X"33821b34",
X"02b90533",
X"903d3371",
X"882b075a",
X"5c78841b",
X"2302bb05",
X"33028405",
X"ba053371",
X"882b0756",
X"5c74ab38",
X"0280ca05",
X"33028405",
X"80c90533",
X"71982b71",
X"902b0796",
X"3d337088",
X"2b720702",
X"940580c7",
X"05337107",
X"51525357",
X"5e5c7476",
X"31783179",
X"842a903d",
X"33547171",
X"31535656",
X"80d2cd3f",
X"83e08008",
X"82057088",
X"1c0c83e0",
X"8008e08a",
X"05565674",
X"83dffe26",
X"83388257",
X"83fff676",
X"27853883",
X"57893986",
X"5676802e",
X"80db3876",
X"7a347683",
X"2e098106",
X"b0380280",
X"d6053302",
X"840580d5",
X"05337198",
X"2b71902b",
X"07993d33",
X"70882b72",
X"07029405",
X"80d30533",
X"71077f90",
X"050c525e",
X"57585686",
X"39771b90",
X"1b0c841a",
X"228c1b08",
X"1971842a",
X"05941c0c",
X"5d800b81",
X"1b347983",
X"e0900c80",
X"567583e0",
X"800c973d",
X"0d04e93d",
X"0d83e090",
X"08568554",
X"75802e81",
X"8238800b",
X"81173499",
X"3de01146",
X"6a548a3d",
X"705458ec",
X"0551f6e5",
X"3f83e080",
X"085483e0",
X"800880df",
X"38893d33",
X"5473802e",
X"913802ab",
X"05337084",
X"2a810651",
X"5574802e",
X"86388354",
X"80c13976",
X"51f4893f",
X"83e08008",
X"a0170c02",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"9c1c0c52",
X"78981b0c",
X"53565957",
X"810b8117",
X"34745473",
X"83e0800c",
X"993d0d04",
X"f53d0d7d",
X"7f617283",
X"e090085a",
X"5d5d595c",
X"807b0c85",
X"5775802e",
X"81e03881",
X"16338106",
X"55845774",
X"802e81d2",
X"38913974",
X"81173486",
X"39800b81",
X"17348157",
X"81c0399c",
X"16089817",
X"08315574",
X"78278338",
X"74587780",
X"2e81a938",
X"98160870",
X"83ff0656",
X"577480cf",
X"38821633",
X"ff057789",
X"2a067081",
X"ff065a55",
X"78a03876",
X"8738a016",
X"08558d39",
X"a4160851",
X"f0e93f83",
X"e0800855",
X"817527ff",
X"a83874a4",
X"170ca416",
X"0851f283",
X"3f83e080",
X"085583e0",
X"8008802e",
X"ff893883",
X"e0800819",
X"a8170c98",
X"160883ff",
X"06848071",
X"31515577",
X"75278338",
X"77557483",
X"ffff0654",
X"98160883",
X"ff0653a8",
X"16085279",
X"577b8338",
X"7b577651",
X"9ad33f83",
X"e08008fe",
X"d0389816",
X"08159817",
X"0c741a78",
X"76317c08",
X"177d0c59",
X"5afed339",
X"80577683",
X"e0800c8d",
X"3d0d04fa",
X"3d0d7883",
X"e0900855",
X"56855573",
X"802e81e3",
X"38811433",
X"81065384",
X"5572802e",
X"81d5389c",
X"14085372",
X"76278338",
X"72569814",
X"0857800b",
X"98150c75",
X"802e81b9",
X"38821433",
X"70892b56",
X"5376802e",
X"b7387452",
X"ff165180",
X"cdce3f83",
X"e08008ff",
X"18765470",
X"53585380",
X"cdbe3f83",
X"e0800873",
X"26963874",
X"30707806",
X"7098170c",
X"777131a4",
X"17085258",
X"51538939",
X"a0140870",
X"a4160c53",
X"747627b9",
X"387251ee",
X"d63f83e0",
X"80085381",
X"0b83e080",
X"08278b38",
X"88140883",
X"e0800826",
X"8838800b",
X"811534b0",
X"3983e080",
X"08a4150c",
X"98140815",
X"98150c75",
X"753156c4",
X"39981408",
X"16709816",
X"0c735256",
X"efc53f83",
X"e080088c",
X"3883e080",
X"08811534",
X"81559439",
X"821433ff",
X"0576892a",
X"0683e080",
X"0805a815",
X"0c805574",
X"83e0800c",
X"883d0d04",
X"ef3d0d63",
X"56855583",
X"e0900880",
X"2e80d238",
X"933df405",
X"84170c64",
X"53883d70",
X"53765257",
X"f1cf3f83",
X"e0800855",
X"83e08008",
X"b438883d",
X"33547380",
X"2ea13802",
X"a7053370",
X"842a7081",
X"06515555",
X"83557380",
X"2e973876",
X"51eef53f",
X"83e08008",
X"88170c75",
X"51efa63f",
X"83e08008",
X"557483e0",
X"800c933d",
X"0d04e43d",
X"0d6ea13d",
X"08405e85",
X"5683e090",
X"08802e84",
X"85389e3d",
X"f405841f",
X"0c7e9838",
X"7d51eef5",
X"3f83e080",
X"085683ee",
X"39814181",
X"f6398341",
X"81f13993",
X"3d7f9605",
X"4159807f",
X"8295055e",
X"56756081",
X"ff053483",
X"41901e08",
X"762e81d3",
X"38a0547d",
X"2270852b",
X"83e00654",
X"58901e08",
X"52785196",
X"dc3f83e0",
X"80084183",
X"e08008ff",
X"b8387833",
X"5c7b802e",
X"ffb4388b",
X"193370bf",
X"06718106",
X"52435574",
X"802e80de",
X"387b81bf",
X"0655748f",
X"2480d338",
X"9a193355",
X"7480cb38",
X"f31d7058",
X"5d815675",
X"8b2e0981",
X"0685388e",
X"568b3975",
X"9a2e0981",
X"0683389c",
X"56751970",
X"70810552",
X"33713381",
X"1a821a5f",
X"5b525b55",
X"74863879",
X"77348539",
X"80df7734",
X"777b5757",
X"7aa02e09",
X"8106c038",
X"81567b81",
X"e5327030",
X"709f2a51",
X"51557bae",
X"2e933874",
X"802e8e38",
X"61832a70",
X"81065155",
X"74802e97",
X"387d51ed",
X"df3f83e0",
X"80084183",
X"e0800887",
X"38901e08",
X"feaf3880",
X"60347580",
X"2e88387c",
X"527f518e",
X"823f6080",
X"2e863880",
X"0b901f0c",
X"60566083",
X"2e853860",
X"81d03889",
X"1f57901e",
X"08802e81",
X"a8388056",
X"75197033",
X"515574a0",
X"2ea03874",
X"852e0981",
X"06843881",
X"e5557477",
X"70810559",
X"34811670",
X"81ff0657",
X"55877627",
X"d7388819",
X"335574a0",
X"2ea938ae",
X"77708105",
X"59348856",
X"75197033",
X"515574a0",
X"2e953874",
X"77708105",
X"59348116",
X"7081ff06",
X"57558a76",
X"27e2388b",
X"19337f88",
X"05349f19",
X"339e1a33",
X"71982b71",
X"902b079d",
X"1c337088",
X"2b72079c",
X"1e337107",
X"640c5299",
X"1d33981e",
X"3371882b",
X"07535153",
X"57595674",
X"7f840523",
X"97193396",
X"1a337188",
X"2b075656",
X"747f8605",
X"23807734",
X"7d51ebf0",
X"3f83e080",
X"08833270",
X"30707207",
X"9f2c83e0",
X"80080652",
X"5656961f",
X"3355748a",
X"38891f52",
X"961f518c",
X"8e3f7583",
X"e0800c9e",
X"3d0d04f4",
X"3d0d7e8f",
X"3dec1156",
X"56589053",
X"f0155277",
X"51e0d23f",
X"83e08008",
X"80d63878",
X"902e0981",
X"0680cd38",
X"02ab0533",
X"80faa80b",
X"80faa833",
X"5758568c",
X"3974762e",
X"8a388417",
X"70335657",
X"74f33876",
X"33705755",
X"74802eac",
X"38821722",
X"708a2b90",
X"3dec0556",
X"70555656",
X"96800a52",
X"7751e081",
X"3f83e080",
X"08863878",
X"752e8538",
X"80568539",
X"81173356",
X"7583e080",
X"0c8e3d0d",
X"04fc3d0d",
X"76705255",
X"8b953f83",
X"e0800815",
X"ff055473",
X"752e8e38",
X"73335372",
X"ae2e8638",
X"ff1454ef",
X"39775281",
X"14518aad",
X"3f83e080",
X"08307083",
X"e0800807",
X"802583e0",
X"800c5386",
X"3d0d04fc",
X"3d0d7670",
X"5255e6ee",
X"3f83e080",
X"08548153",
X"83e08008",
X"80c13874",
X"51e6b13f",
X"83e08008",
X"80f7c853",
X"83e08008",
X"5253ff91",
X"3f83e080",
X"08a13880",
X"f7cc5272",
X"51ff823f",
X"83e08008",
X"923880f7",
X"d0527251",
X"fef33f83",
X"e0800880",
X"2e833881",
X"54735372",
X"83e0800c",
X"863d0d04",
X"fd3d0d75",
X"705254e6",
X"8d3f8153",
X"83e08008",
X"98387351",
X"e5d63f83",
X"e3880852",
X"83e08008",
X"51feba3f",
X"83e08008",
X"537283e0",
X"800c853d",
X"0d04df3d",
X"0da43d08",
X"70525edb",
X"f43f83e0",
X"80083395",
X"3d565473",
X"963880fd",
X"e4527451",
X"898d3f9a",
X"397d5278",
X"51defc3f",
X"84d0397d",
X"51dbda3f",
X"83e08008",
X"527451db",
X"8a3f8043",
X"80428041",
X"804083e3",
X"90085294",
X"3d70525d",
X"e1e43f83",
X"e0800859",
X"800b83e0",
X"8008555b",
X"83e08008",
X"7b2e9438",
X"811b7452",
X"5be4e63f",
X"83e08008",
X"5483e080",
X"08ee3880",
X"5aff5f79",
X"09709f2c",
X"7b065b54",
X"7a7a2484",
X"38ff1b5a",
X"f61a7009",
X"709f2c72",
X"067bff12",
X"5a5a5255",
X"55807525",
X"95387651",
X"e4ab3f83",
X"e0800876",
X"ff185855",
X"57738024",
X"ed38747f",
X"2e8638a1",
X"b53f745f",
X"78ff1b70",
X"585d5880",
X"7a259538",
X"7751e481",
X"3f83e080",
X"0876ff18",
X"58555873",
X"8024ed38",
X"800b83e7",
X"c00c800b",
X"83e7e80c",
X"80f7d451",
X"8d8c3f81",
X"800b83e7",
X"e80c80f7",
X"dc518cfe",
X"3fa80b83",
X"e7c00c76",
X"802e80e4",
X"3883e7c0",
X"08777932",
X"70307072",
X"07802570",
X"872b83e7",
X"e80c5156",
X"78535656",
X"e3b83f83",
X"e0800880",
X"2e883880",
X"f7e4518c",
X"c53f7651",
X"e2fa3f83",
X"e0800852",
X"80f98451",
X"8cb43f76",
X"51e3823f",
X"83e08008",
X"83e7c008",
X"55577574",
X"258638a8",
X"1656f739",
X"7583e7c0",
X"0c86f076",
X"24ff9838",
X"87980b83",
X"e7c00c77",
X"802eb138",
X"7751e2b8",
X"3f83e080",
X"08785255",
X"e2d83f80",
X"f7ec5483",
X"e080088d",
X"38873980",
X"763481d0",
X"3980f7e8",
X"54745373",
X"5280f7bc",
X"518bd33f",
X"805480f7",
X"c4518bca",
X"3f811454",
X"73a82e09",
X"8106ef38",
X"868da051",
X"9da83f80",
X"52903d70",
X"525780c3",
X"b33f8352",
X"765180c3",
X"ab3f6281",
X"8f386180",
X"2e80fb38",
X"7b5473ff",
X"2e963878",
X"802e818a",
X"387851e1",
X"dc3f83e0",
X"8008ff15",
X"5559e739",
X"78802e80",
X"f5387851",
X"e1d83f83",
X"e0800880",
X"2efc8e38",
X"7851e1a0",
X"3f83e080",
X"085280f7",
X"b85183e0",
X"3f83e080",
X"08a3387c",
X"5185983f",
X"83e08008",
X"5574ff16",
X"56548074",
X"25ae3874",
X"1d703355",
X"5673af2e",
X"fecd38e9",
X"397851e0",
X"e13f83e0",
X"8008527c",
X"5184d03f",
X"8f397f88",
X"29601005",
X"7a056105",
X"5afc9039",
X"62802efb",
X"d1388052",
X"765180c2",
X"8b3fa33d",
X"0d04803d",
X"0d9088b8",
X"337081ff",
X"0670842a",
X"81327081",
X"06515151",
X"5170802e",
X"8d38a80b",
X"9088b834",
X"b80b9088",
X"b8347083",
X"e0800c82",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067085",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d3898",
X"0b9088b8",
X"34b80b90",
X"88b83470",
X"83e0800c",
X"823d0d04",
X"930b9088",
X"bc34ff0b",
X"9088a834",
X"04ff3d0d",
X"028f0533",
X"52800b90",
X"88bc348a",
X"519aef3f",
X"df3f80f8",
X"0b9088a0",
X"34800b90",
X"888834fa",
X"12527190",
X"88803480",
X"0b908898",
X"34719088",
X"90349088",
X"b8528072",
X"34b87234",
X"833d0d04",
X"803d0d02",
X"8b053351",
X"709088b4",
X"34febf3f",
X"83e08008",
X"802ef638",
X"823d0d04",
X"803d0d84",
X"39a5a63f",
X"fed93f83",
X"e0800880",
X"2ef33890",
X"88b43370",
X"81ff0683",
X"e0800c51",
X"823d0d04",
X"803d0da3",
X"0b9088bc",
X"34ff0b90",
X"88a83490",
X"88b851a8",
X"7134b871",
X"34823d0d",
X"04803d0d",
X"9088bc33",
X"70982b70",
X"802583e0",
X"800c5151",
X"823d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"832a8132",
X"70810651",
X"51515170",
X"802ee838",
X"b00b9088",
X"b834b80b",
X"9088b834",
X"823d0d04",
X"803d0d90",
X"80ac0881",
X"0683e080",
X"0c823d0d",
X"04fd3d0d",
X"75775454",
X"80732594",
X"38737081",
X"05553352",
X"80f7f051",
X"87843fff",
X"1353e939",
X"853d0d04",
X"fd3d0d75",
X"77535473",
X"33517089",
X"38713351",
X"70802ea1",
X"38733372",
X"33525372",
X"71278538",
X"ff519439",
X"70732785",
X"3881518b",
X"39811481",
X"135354d3",
X"39805170",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"77545472",
X"337081ff",
X"06525270",
X"802ea338",
X"7181ff06",
X"8114ffbf",
X"12535452",
X"70992689",
X"38a01270",
X"81ff0653",
X"51717470",
X"81055634",
X"d2398074",
X"34853d0d",
X"04ffbd3d",
X"0d80c63d",
X"0852a53d",
X"705254ff",
X"b33f80c7",
X"3d085285",
X"3d705253",
X"ffa63f72",
X"527351fe",
X"df3f80c5",
X"3d0d04fe",
X"3d0d7476",
X"53537170",
X"81055333",
X"51707370",
X"81055534",
X"70f03884",
X"3d0d04fe",
X"3d0d7452",
X"80723352",
X"5370732e",
X"8d388112",
X"81147133",
X"53545270",
X"f5387283",
X"e0800c84",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"baa63f83",
X"e080087a",
X"27ee3874",
X"802e80dd",
X"38745275",
X"51ba913f",
X"83e08008",
X"75537652",
X"54ba953f",
X"83e08008",
X"7a537552",
X"56b9f93f",
X"83e08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"e08008c5",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9f",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fc813f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd53f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbb13f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83e0940c",
X"7183e098",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383e094",
X"085283e0",
X"980851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"bdbe5351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fc3d",
X"0d765574",
X"83e39c08",
X"2eaf3880",
X"53745187",
X"c13f83e0",
X"800881ff",
X"06ff1470",
X"81ff0672",
X"30709f2a",
X"51525553",
X"5472802e",
X"843871dd",
X"3873fe38",
X"7483e39c",
X"0c863d0d",
X"04ff3d0d",
X"ff0b83e3",
X"9c0c84a5",
X"3f815187",
X"853f83e0",
X"800881ff",
X"065271ee",
X"3881d33f",
X"7183e080",
X"0c833d0d",
X"04fc3d0d",
X"76028405",
X"a2052202",
X"8805a605",
X"227a5455",
X"5555ff82",
X"3f72802e",
X"a03883e3",
X"b0143375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552dd",
X"39800b83",
X"e0800c86",
X"3d0d04fc",
X"3d0d7678",
X"7a115653",
X"55805371",
X"742e9338",
X"72155170",
X"3383e3b0",
X"13348112",
X"81145452",
X"ea39800b",
X"83e0800c",
X"863d0d04",
X"fd3d0d90",
X"5483e39c",
X"085186f4",
X"3f83e080",
X"0881ff06",
X"ff157130",
X"71307073",
X"079f2a72",
X"9f2a0652",
X"55525553",
X"72db3885",
X"3d0d0480",
X"3d0d83e3",
X"a8081083",
X"e3a00807",
X"9080a80c",
X"823d0d04",
X"800b83e3",
X"a80ce43f",
X"04810b83",
X"e3a80cdb",
X"3f04ed3f",
X"047183e3",
X"a40c0480",
X"3d0d8051",
X"f43f810b",
X"83e3a80c",
X"810b83e3",
X"a00cffbb",
X"3f823d0d",
X"04803d0d",
X"72307074",
X"07802583",
X"e3a00c51",
X"ffa53f82",
X"3d0d0480",
X"3d0d028b",
X"05339080",
X"a40c9080",
X"a8087081",
X"06515170",
X"f5389080",
X"a4087081",
X"ff0683e0",
X"800c5182",
X"3d0d0480",
X"3d0d81ff",
X"51d13f83",
X"e0800881",
X"ff0683e0",
X"800c823d",
X"0d04803d",
X"0d73902b",
X"73079080",
X"b40c823d",
X"0d0404fb",
X"3d0d7802",
X"84059f05",
X"3370982b",
X"55575572",
X"80259b38",
X"7580ff06",
X"56805280",
X"f751e03f",
X"83e08008",
X"81ff0654",
X"73812680",
X"ff388051",
X"fee73fff",
X"a23f8151",
X"fedf3fff",
X"9a3f7551",
X"feed3f74",
X"982a51fe",
X"e63f7490",
X"2a7081ff",
X"065253fe",
X"da3f7488",
X"2a7081ff",
X"065253fe",
X"ce3f7481",
X"ff0651fe",
X"c63f8155",
X"7580c02e",
X"09810686",
X"38819555",
X"8d397580",
X"c82e0981",
X"06843881",
X"87557451",
X"fea53f8a",
X"55fec83f",
X"83e08008",
X"81ff0670",
X"982b5454",
X"7280258c",
X"38ff1570",
X"81ff0656",
X"5374e238",
X"7383e080",
X"0c873d0d",
X"04fa3d0d",
X"fdc53f80",
X"51fdda3f",
X"8a54fe93",
X"3fff1470",
X"81ff0655",
X"5373f338",
X"73745355",
X"80c051fe",
X"a63f83e0",
X"800881ff",
X"06547381",
X"2e098106",
X"829f3883",
X"aa5280c8",
X"51fe8c3f",
X"83e08008",
X"81ff0653",
X"72812e09",
X"810681a8",
X"38745487",
X"3d741154",
X"56fdc83f",
X"83e08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e53802",
X"9a053353",
X"72812e09",
X"810681d9",
X"38029b05",
X"335380ce",
X"90547281",
X"aa2e8d38",
X"81c73980",
X"e4518b9a",
X"3fff1454",
X"73802e81",
X"b838820a",
X"5281e951",
X"fda53f83",
X"e0800881",
X"ff065372",
X"de387252",
X"80fa51fd",
X"923f83e0",
X"800881ff",
X"06537281",
X"90387254",
X"731653fc",
X"d63f83e0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e8",
X"38873d33",
X"70862a70",
X"81065154",
X"548c5572",
X"80e33884",
X"5580de39",
X"745281e9",
X"51fccc3f",
X"83e08008",
X"81ff0653",
X"825581e9",
X"56817327",
X"86387355",
X"80c15680",
X"ce90548a",
X"3980e451",
X"8a8c3fff",
X"14547380",
X"2ea93880",
X"527551fc",
X"9a3f83e0",
X"800881ff",
X"065372e1",
X"38848052",
X"80d051fc",
X"863f83e0",
X"800881ff",
X"06537280",
X"2e833880",
X"557483e3",
X"ac348051",
X"fb873ffb",
X"c23f883d",
X"0d04fb3d",
X"0d775480",
X"0b83e3ac",
X"3370832a",
X"70810651",
X"55575572",
X"752e0981",
X"06853873",
X"892b5473",
X"5280d151",
X"fbbd3f83",
X"e0800881",
X"ff065372",
X"bd3882b8",
X"c054fb83",
X"3f83e080",
X"0881ff06",
X"537281ff",
X"2e098106",
X"8938ff14",
X"5473e738",
X"9f397281",
X"fe2e0981",
X"06963883",
X"e7b05283",
X"e3b051fa",
X"ed3ffad3",
X"3ffad03f",
X"83398155",
X"8051fa89",
X"3ffac43f",
X"7481ff06",
X"83e0800c",
X"873d0d04",
X"fb3d0d77",
X"83e3b056",
X"548151f9",
X"ec3f83e3",
X"ac337083",
X"2a708106",
X"51545672",
X"85387389",
X"2b547352",
X"80d851fa",
X"b63f83e0",
X"800881ff",
X"06537280",
X"e43881ff",
X"51f9d43f",
X"81fe51f9",
X"ce3f8480",
X"53747081",
X"05563351",
X"f9c13fff",
X"137083ff",
X"ff065153",
X"72eb3872",
X"51f9b03f",
X"7251f9ab",
X"3ff9d03f",
X"83e08008",
X"9f0653a7",
X"88547285",
X"2e8c3899",
X"3980e451",
X"87c43fff",
X"1454f9b3",
X"3f83e080",
X"0881ff2e",
X"843873e9",
X"388051f8",
X"e43ff99f",
X"3f800b83",
X"e0800c87",
X"3d0d0471",
X"83e7b40c",
X"8880800b",
X"83e7b00c",
X"8480800b",
X"83e7b80c",
X"04fd3d0d",
X"77701755",
X"7705ff1a",
X"535371ff",
X"2e943873",
X"70810555",
X"33517073",
X"70810555",
X"34ff1252",
X"e939853d",
X"0d04fb3d",
X"0d87a681",
X"0b83e7b4",
X"08565675",
X"3383a680",
X"1634a054",
X"83a08053",
X"83e7b408",
X"5283e7b0",
X"0851ffb1",
X"3fa05483",
X"a4805383",
X"e7b40852",
X"83e7b008",
X"51ff9e3f",
X"905483a8",
X"805383e7",
X"b4085283",
X"e7b00851",
X"ff8b3fa0",
X"53805283",
X"e7b80883",
X"a0800551",
X"86953fa0",
X"53805283",
X"e7b80883",
X"a4800551",
X"86853f90",
X"53805283",
X"e7b80883",
X"a8800551",
X"85f53fff",
X"763483a0",
X"80548053",
X"83e7b408",
X"5283e7b8",
X"0851fec5",
X"3f80d080",
X"5483b080",
X"5383e7b4",
X"085283e7",
X"b80851fe",
X"b03f87ba",
X"3fa25480",
X"5383e7b8",
X"088c8005",
X"5280fb9c",
X"51fe9a3f",
X"860b87a8",
X"8334800b",
X"87a88234",
X"800b87a0",
X"9a34af0b",
X"87a09634",
X"bf0b87a0",
X"9734800b",
X"87a09834",
X"9f0b87a0",
X"9934800b",
X"87a09b34",
X"e00b87a8",
X"8934a20b",
X"87a88034",
X"830b87a4",
X"8f34820b",
X"87a88134",
X"873d0d04",
X"fc3d0d83",
X"a0805480",
X"5383e7b8",
X"085283e7",
X"b40851fd",
X"b83f80d0",
X"805483b0",
X"805383e7",
X"b8085283",
X"e7b40851",
X"fda33fa0",
X"5483a080",
X"5383e7b8",
X"085283e7",
X"b40851fd",
X"903fa054",
X"83a48053",
X"83e7b808",
X"5283e7b4",
X"0851fcfd",
X"3f905483",
X"a8805383",
X"e7b80852",
X"83e7b408",
X"51fcea3f",
X"83e7b408",
X"5583a680",
X"153387a6",
X"8134863d",
X"0d04fa3d",
X"0d787052",
X"55c1e33f",
X"83ffff0b",
X"83e08008",
X"25a93874",
X"51c1e43f",
X"83e08008",
X"9e3883e0",
X"80085788",
X"3dfc0554",
X"84808053",
X"83e7b408",
X"527451ff",
X"bf963fff",
X"bedc3f88",
X"3d0d04fa",
X"3d0d7870",
X"5255c1a2",
X"3f83ffff",
X"0b83e080",
X"08259638",
X"8057883d",
X"fc055484",
X"80805383",
X"e7b40852",
X"7451c095",
X"3f883d0d",
X"04803d0d",
X"90809008",
X"810683e0",
X"800c823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087081",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fd0676",
X"1007720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870822c",
X"bf0683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe830676",
X"822b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087088",
X"2c870683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f1ff06",
X"76882b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"912cbf06",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fc87",
X"ffff0676",
X"912b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087099",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70ffbf0a",
X"0676992b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90808008",
X"70882c81",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"0870892c",
X"810683e0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708a",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8b2c8106",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708c2cbf",
X"0683e080",
X"0c51823d",
X"0d04fe3d",
X"0d7481e6",
X"29872a90",
X"80a00c84",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70810554",
X"34ff1151",
X"f039843d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"8405540c",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"84808053",
X"80528880",
X"0a51ffb3",
X"3f818080",
X"53805282",
X"800a51c6",
X"3f843d0d",
X"04803d0d",
X"8151fcaa",
X"3f72802e",
X"90388051",
X"fdfe3fcd",
X"3f83e7bc",
X"3351fdf4",
X"3f8151fc",
X"bb3f8051",
X"fcb63f80",
X"51fc873f",
X"823d0d04",
X"fd3d0d75",
X"52805480",
X"ff722588",
X"38810bff",
X"80135354",
X"ffbf1251",
X"70992686",
X"38e01252",
X"b039ff9f",
X"12519971",
X"27a738d0",
X"12e01354",
X"51708926",
X"85387252",
X"9839728f",
X"26853872",
X"528f3971",
X"ba2e0981",
X"0685389a",
X"52833980",
X"5273802e",
X"85388180",
X"12527181",
X"ff0683e0",
X"800c853d",
X"0d04803d",
X"0d84d8c0",
X"51807170",
X"81055334",
X"7084e0c0",
X"2e098106",
X"f038823d",
X"0d04fe3d",
X"0d029705",
X"3351fef4",
X"3f83e080",
X"0881ff06",
X"83e7c008",
X"54528073",
X"249b3883",
X"e7e40813",
X"7283e7e8",
X"08075353",
X"71733483",
X"e7c00881",
X"0583e7c0",
X"0c843d0d",
X"04fa3d0d",
X"82800a1b",
X"55805788",
X"3dfc0554",
X"79537452",
X"7851ffba",
X"ac3f883d",
X"0d04fe3d",
X"0d83e7d8",
X"08527451",
X"c1903f83",
X"e080088c",
X"38765375",
X"5283e7d8",
X"0851c63f",
X"843d0d04",
X"fe3d0d83",
X"e7d80853",
X"75527451",
X"ffbbce3f",
X"83e08008",
X"8d387753",
X"765283e7",
X"d80851ff",
X"a03f843d",
X"0d04fe3d",
X"0d83e7d8",
X"0851ffba",
X"c13f83e0",
X"80088180",
X"802e0981",
X"06883883",
X"c1808053",
X"9c3983e7",
X"d80851ff",
X"baa43f83",
X"e0800880",
X"d0802e09",
X"81069338",
X"83c1b080",
X"5383e080",
X"085283e7",
X"d80851fe",
X"d43f843d",
X"0d04803d",
X"0df9fc3f",
X"83e08008",
X"842980fb",
X"c0057008",
X"83e0800c",
X"51823d0d",
X"04ed3d0d",
X"80448043",
X"80428041",
X"80705a5b",
X"fdcc3f80",
X"0b83e7c0",
X"0c800b83",
X"e7e80c80",
X"f8bc51e9",
X"c53f8180",
X"0b83e7e8",
X"0c80f8c0",
X"51e9b73f",
X"80d00b83",
X"e7c00c78",
X"30707a07",
X"80257087",
X"2b83e7e8",
X"0c5155f8",
X"ed3f83e0",
X"80085280",
X"f8c851e9",
X"913f80f8",
X"0b83e7c0",
X"0c788132",
X"70307072",
X"07802570",
X"872b83e7",
X"e80c5156",
X"569db73f",
X"83e08008",
X"5280f8d8",
X"51e8e73f",
X"81a00b83",
X"e7c00c78",
X"82327030",
X"70720780",
X"2570872b",
X"83e7e80c",
X"515656fe",
X"c53f83e0",
X"80085280",
X"f8e851e8",
X"bd3f81c8",
X"0b83e7c0",
X"0c788332",
X"70307072",
X"07802570",
X"872b83e7",
X"e80c5156",
X"83e7d808",
X"5256ffb5",
X"983f83e0",
X"80085280",
X"f8f051e8",
X"8d3f8298",
X"0b83e7c0",
X"0c810b83",
X"e7c45b58",
X"83e7c008",
X"83197a32",
X"70307072",
X"07802570",
X"872b83e7",
X"e80c5157",
X"8e3d7055",
X"ff1b5457",
X"57579af9",
X"3f797084",
X"055b0851",
X"ffb4ce3f",
X"745483e0",
X"80085377",
X"5280f8f8",
X"51e7bf3f",
X"a81783e7",
X"c00c8118",
X"5877852e",
X"098106ff",
X"af3883b8",
X"0b83e7c0",
X"0c788832",
X"70307072",
X"07802570",
X"872b83e7",
X"e80c5156",
X"56f7b93f",
X"80f98855",
X"83e08008",
X"802e8f38",
X"83e7d408",
X"51ffb3f9",
X"3f83e080",
X"08557452",
X"80f99051",
X"e6ec3f84",
X"880b83e7",
X"c00c7889",
X"32703070",
X"72078025",
X"70872b83",
X"e7e80c51",
X"5780f99c",
X"5255e6ca",
X"3f868da0",
X"51f8b33f",
X"8052913d",
X"7052559e",
X"bf3f8352",
X"74519eb8",
X"3f635574",
X"839c3861",
X"19597880",
X"25853874",
X"59903989",
X"79258538",
X"89598739",
X"78892682",
X"fb387882",
X"2b5580f7",
X"90150804",
X"f5d43f83",
X"e0800861",
X"57557581",
X"2e098106",
X"893883e0",
X"80081055",
X"903975ff",
X"2e098106",
X"883883e0",
X"8008812c",
X"55907525",
X"85389055",
X"88397480",
X"24833881",
X"557451f5",
X"ae3f82b0",
X"3999fe3f",
X"83e08008",
X"61055574",
X"80258538",
X"80558839",
X"87752583",
X"38875574",
X"518de13f",
X"828e39f5",
X"9e3f83e0",
X"80086105",
X"55748025",
X"85388055",
X"88398675",
X"25833886",
X"557451f5",
X"973f81ec",
X"39608738",
X"62802e81",
X"e33883e3",
X"8c0883e3",
X"880cadec",
X"0b83e390",
X"0c83e7d8",
X"0851d5e2",
X"3ffa8f3f",
X"81c63960",
X"56807625",
X"9838ad8b",
X"0b83e390",
X"0c83e7b4",
X"15700852",
X"55d5c33f",
X"74085292",
X"39758025",
X"923883e7",
X"b4150851",
X"ffb1c03f",
X"8052fc19",
X"51b83962",
X"802e818c",
X"3883e7b4",
X"15700883",
X"e7c40872",
X"0c83e7c4",
X"0cfc1a70",
X"5351558c",
X"ae3f83e0",
X"80085680",
X"518ca43f",
X"83e08008",
X"52745188",
X"bd3f7552",
X"805188b6",
X"3f80d539",
X"60558075",
X"25b63883",
X"e3980883",
X"e3880cad",
X"ec0b83e3",
X"900c83e7",
X"d40851d4",
X"cd3f83e7",
X"d40851d1",
X"ee3f83e0",
X"800881ff",
X"06705255",
X"f3f73f74",
X"802e9d38",
X"8155a139",
X"74802594",
X"3883e7d4",
X"0851ffb0",
X"b23f8051",
X"f3db3f84",
X"39628738",
X"7a802ef9",
X"b7388055",
X"7483e080",
X"0c953d0d",
X"04fe3d0d",
X"f4873f83",
X"e0800880",
X"2e863880",
X"51818a39",
X"f48c3f83",
X"e0800880",
X"fe38f4ac",
X"3f83e080",
X"08802eb9",
X"388151f1",
X"e93f8051",
X"f3c23fed",
X"e13f800b",
X"83e7c00c",
X"f8df3f83",
X"e0800853",
X"ff0b83e7",
X"c00cefd4",
X"3f7280cb",
X"3883e7bc",
X"3351f39c",
X"3f7251f1",
X"b93f80c0",
X"39f3d43f",
X"83e08008",
X"802eb538",
X"8151f1a6",
X"3f8051f2",
X"ff3fed9e",
X"3fad8b0b",
X"83e3900c",
X"83e7c408",
X"51d2ff3f",
X"ff0b83e7",
X"c00cef90",
X"3f83e7c4",
X"08528051",
X"86b43f81",
X"51f4c63f",
X"843d0d04",
X"fb3d0d80",
X"0b83e7bc",
X"34908080",
X"52868480",
X"8051ffb2",
X"f23f83e0",
X"80088197",
X"388a993f",
X"80fdd451",
X"ffb7b13f",
X"83e08008",
X"559c800a",
X"5480c080",
X"5380f9a4",
X"5283e080",
X"0851f6ac",
X"3f83e7d8",
X"085380f9",
X"b4527451",
X"ffb1fa3f",
X"83e08008",
X"8438f6ba",
X"3f83e7dc",
X"085380f9",
X"c0527451",
X"ffb1e23f",
X"83e08008",
X"b638873d",
X"fc055484",
X"80805386",
X"a8808052",
X"83e7dc08",
X"51ffafed",
X"3f83e080",
X"08933875",
X"8480802e",
X"09810689",
X"38810b83",
X"e7bc3487",
X"39800b83",
X"e7bc3483",
X"e7bc3351",
X"f1a63f81",
X"51f3923f",
X"93ca3f81",
X"51f38a3f",
X"8151fda1",
X"3ffa3983",
X"e08c0802",
X"83e08c0c",
X"fb3d0d02",
X"80f9cc0b",
X"83e38c0c",
X"80f9d00b",
X"83e3840c",
X"80f9d40b",
X"83e3980c",
X"80f9d80b",
X"83e3940c",
X"83e08c08",
X"fc050c80",
X"0b83e7c4",
X"0b83e08c",
X"08f8050c",
X"83e08c08",
X"f4050cff",
X"aff53f83",
X"e0800886",
X"05fc0683",
X"e08c08f0",
X"050c0283",
X"e08c08f0",
X"0508310d",
X"833d7083",
X"e08c08f8",
X"05087084",
X"0583e08c",
X"08f8050c",
X"0c51ffac",
X"b63f83e0",
X"8c08f405",
X"08810583",
X"e08c08f4",
X"050c83e0",
X"8c08f405",
X"08882e09",
X"8106ffab",
X"38869480",
X"8051e9cf",
X"3fff0b83",
X"e7c00c80",
X"0b83e7e8",
X"0c84d8c0",
X"0b83e7e4",
X"0c8151ed",
X"f53f8151",
X"ee9a3f80",
X"51ee953f",
X"8151eebb",
X"3f8251ee",
X"e33f8051",
X"ef8b3f80",
X"51efb53f",
X"80d1ae52",
X"8051deb3",
X"3ffcd93f",
X"83e08c08",
X"fc05080d",
X"800b83e0",
X"800c873d",
X"0d83e08c",
X"0c04803d",
X"0d81ff51",
X"800b83e7",
X"f81234ff",
X"115170f4",
X"38823d0d",
X"04ff3d0d",
X"73703353",
X"51811133",
X"71347181",
X"1234833d",
X"0d04ff3d",
X"0d83ea94",
X"08a82e09",
X"81068b38",
X"83eaac08",
X"83ea940c",
X"8739a80b",
X"83ea940c",
X"83ea9408",
X"86057081",
X"ff065252",
X"d4bb3f83",
X"3d0d04fb",
X"3d0d7779",
X"56568070",
X"71555552",
X"717525ac",
X"38721670",
X"33701470",
X"81ff0655",
X"51515171",
X"74278938",
X"81127081",
X"ff065351",
X"71811470",
X"83ffff06",
X"55525474",
X"7324d638",
X"7183e080",
X"0c873d0d",
X"04fb3d0d",
X"77568939",
X"f9f33f83",
X"51eee33f",
X"d5c23f83",
X"e0800880",
X"2eee3883",
X"ea940886",
X"057081ff",
X"065253d3",
X"c83f810b",
X"9088d434",
X"f9cb3f83",
X"51eebb3f",
X"9088d433",
X"7081ff06",
X"55537380",
X"2eea3873",
X"862a7081",
X"06515372",
X"ffbe3873",
X"982b5380",
X"732480de",
X"38d4b23f",
X"83e08008",
X"5583e080",
X"0880cf38",
X"74167582",
X"2b545490",
X"88c01333",
X"74348115",
X"5574852e",
X"098106e8",
X"38753383",
X"e7f83481",
X"163383e7",
X"f9348216",
X"3383e7fa",
X"34831633",
X"83e7fb34",
X"845283e7",
X"f851fe93",
X"3f83e080",
X"0881ff06",
X"84173355",
X"5372742e",
X"8738fdce",
X"3ffed139",
X"80e451ed",
X"ad3f873d",
X"0d04f43d",
X"0d7e6059",
X"55805d80",
X"75822b71",
X"83ea9812",
X"0c83eab0",
X"175b5b57",
X"76793477",
X"772e83b7",
X"38765277",
X"51ffaad1",
X"3f8e3dfc",
X"05549053",
X"83ea8052",
X"7751ffaa",
X"8c3f7c56",
X"75902e09",
X"81068393",
X"3883ea80",
X"51fcde3f",
X"83ea8251",
X"fcd73f83",
X"ea8451fc",
X"d03f7683",
X"ea900c77",
X"51ffa7d1",
X"3f80f7cc",
X"5283e080",
X"0851c9f1",
X"3f83e080",
X"08812e09",
X"810680d4",
X"387683ea",
X"a80c820b",
X"83ea8034",
X"ff960b83",
X"ea813477",
X"51ffaa9e",
X"3f83e080",
X"085583e0",
X"80087725",
X"883883e0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83ea8234",
X"7483ea83",
X"347683ea",
X"8434ff80",
X"0b83ea85",
X"34819039",
X"83ea8033",
X"83ea8133",
X"71882b07",
X"565b7483",
X"ffff2e09",
X"810680e8",
X"38fe800b",
X"83eaa80c",
X"810b83ea",
X"900cff0b",
X"83ea8034",
X"ff0b83ea",
X"81347751",
X"ffa9ab3f",
X"83e08008",
X"83eab40c",
X"83e08008",
X"5583e080",
X"08802588",
X"3883e080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"ea823474",
X"83ea8334",
X"7683ea84",
X"34ff800b",
X"83ea8534",
X"810b83ea",
X"8f34a539",
X"7485962e",
X"09810680",
X"fe387583",
X"eaa80c77",
X"51ffa8df",
X"3f83ea8f",
X"3383e080",
X"08075574",
X"83ea8f34",
X"83ea8f33",
X"81065574",
X"802e8338",
X"845783ea",
X"843383ea",
X"85337188",
X"2b07565c",
X"7481802e",
X"098106a1",
X"3883ea82",
X"3383ea83",
X"3371882b",
X"07565bad",
X"80752787",
X"38768207",
X"579c3976",
X"81075796",
X"39748280",
X"2e098106",
X"87387683",
X"07578739",
X"7481ff26",
X"8a387783",
X"ea981b0c",
X"7679348e",
X"3d0d0480",
X"3d0d7284",
X"2983ea98",
X"05700883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"7083e7f0",
X"0c708429",
X"80fd9405",
X"700883ea",
X"ac0c5151",
X"823d0d04",
X"fe3d0d81",
X"51de3f80",
X"0b83e9fc",
X"0c800b83",
X"e9f80cff",
X"0b83e7f4",
X"0ca80b83",
X"ea940cae",
X"51cdf63f",
X"800b83ea",
X"98545280",
X"73708405",
X"550c8112",
X"5271842e",
X"098106ef",
X"38843d0d",
X"04fe3d0d",
X"74028405",
X"96052253",
X"5371802e",
X"96387270",
X"81055433",
X"51ce813f",
X"ff127083",
X"ffff0651",
X"52e73984",
X"3d0d04fe",
X"3d0d0292",
X"05225382",
X"ac51e8a2",
X"3f80c351",
X"cdde3f81",
X"9651e896",
X"3f725283",
X"e7f851ff",
X"b43f7252",
X"83e7f851",
X"f8cd3f83",
X"e0800881",
X"ff0651cd",
X"bb3f843d",
X"0d04ffb1",
X"3d0d80d1",
X"3df80551",
X"f8f73f83",
X"e9fc0881",
X"0583e9fc",
X"0c80cf3d",
X"33cf1170",
X"81ff0651",
X"56567483",
X"2688e638",
X"758f06ff",
X"05567583",
X"e7f4082e",
X"9b387583",
X"26963875",
X"83e7f40c",
X"75842983",
X"ea980570",
X"08535575",
X"51f9fb3f",
X"80762488",
X"c2387584",
X"2983ea98",
X"05557408",
X"802e88b3",
X"3883e7f4",
X"08842983",
X"ea980570",
X"08028805",
X"82b90533",
X"525b5574",
X"80d22e84",
X"b0387480",
X"d2249038",
X"74bf2e9c",
X"387480d0",
X"2e81d538",
X"87f23974",
X"80d32e80",
X"d3387480",
X"d72e81c4",
X"3887e139",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"055656cc",
X"b73f80c1",
X"51cbf13f",
X"f6983f83",
X"eaaf3383",
X"e7f83481",
X"5283e7f8",
X"51cd8e3f",
X"8151fde7",
X"3f748b38",
X"83eaac08",
X"83ea940c",
X"8739a80b",
X"83ea940c",
X"cc823f80",
X"c151cbbc",
X"3ff5e33f",
X"900b83ea",
X"8f338106",
X"56567480",
X"2e833898",
X"5683ea84",
X"3383ea85",
X"3371882b",
X"07565974",
X"81802e09",
X"81069c38",
X"83ea8233",
X"83ea8333",
X"71882b07",
X"5657ad80",
X"75278c38",
X"75818007",
X"56853975",
X"a0075675",
X"83e7f834",
X"ff0b83e7",
X"f934e00b",
X"83e7fa34",
X"800b83e7",
X"fb348452",
X"83e7f851",
X"cc833f84",
X"51869b39",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"055659ca",
X"f73f7951",
X"ffa38c3f",
X"83e08008",
X"802e8a38",
X"80ce51ca",
X"a33f85f1",
X"3980c151",
X"ca9a3fcb",
X"8b3fc9c4",
X"3f83eaa8",
X"08588375",
X"259b3883",
X"ea843383",
X"ea853371",
X"882b07fc",
X"1771297a",
X"05838005",
X"5a51578d",
X"39748180",
X"2918ff80",
X"05588180",
X"57805676",
X"762e9238",
X"c9f63f83",
X"e0800883",
X"e7f81734",
X"811656eb",
X"39c9e53f",
X"83e08008",
X"81ff0677",
X"5383e7f8",
X"5256f4bf",
X"3f83e080",
X"0881ff06",
X"5575752e",
X"09810681",
X"95389451",
X"e3e03fc9",
X"df3f80c1",
X"51c9993f",
X"ca8a3f77",
X"527951ff",
X"a19f3f80",
X"5e80d13d",
X"fdf40554",
X"765383e7",
X"f8527951",
X"ff9fa53f",
X"0282b905",
X"33558159",
X"7480d72e",
X"09810680",
X"c5387752",
X"7951ffa0",
X"f03f80d1",
X"3dfdf005",
X"5476538f",
X"3d70537a",
X"5258ffa0",
X"a83f8056",
X"76762ea2",
X"38751883",
X"e7f81733",
X"71337072",
X"32703070",
X"80257030",
X"7f06811d",
X"5d5f5151",
X"51525b55",
X"db3982ac",
X"51e2db3f",
X"78802e86",
X"3880c351",
X"843980ce",
X"51c88d3f",
X"c8fe3fc7",
X"b73f83d8",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055955",
X"80705d59",
X"80e451e2",
X"a53fc8a4",
X"3f80c151",
X"c7de3f83",
X"ea900879",
X"2e82d638",
X"83eab408",
X"80fc0555",
X"80fd5274",
X"5185c13f",
X"83e08008",
X"5b778224",
X"b238ff18",
X"70872b83",
X"ffff8006",
X"80fbe005",
X"83e7f859",
X"57558180",
X"55757081",
X"05573377",
X"70810559",
X"34ff1570",
X"81ff0651",
X"5574ea38",
X"82853977",
X"82e82e81",
X"a3387782",
X"e92e0981",
X"0681aa38",
X"78587787",
X"32703070",
X"72078025",
X"7a8a3270",
X"30707207",
X"80257307",
X"53545a51",
X"57557580",
X"2e973878",
X"78269238",
X"a00b83e7",
X"f81a3481",
X"197081ff",
X"065a55eb",
X"39811870",
X"81ff0659",
X"558a7827",
X"ffbc388f",
X"5883e7f3",
X"183383e7",
X"f81934ff",
X"187081ff",
X"06595577",
X"8426ea38",
X"9058800b",
X"83e7f819",
X"34811870",
X"81ff0670",
X"982b5259",
X"55748025",
X"e93880c6",
X"557a858f",
X"24843880",
X"c2557483",
X"e7f83480",
X"f10b83e7",
X"fb34810b",
X"83e7fc34",
X"7a83e7f9",
X"347a882c",
X"557483e7",
X"fa3480cb",
X"3982f078",
X"2580c438",
X"7780fd29",
X"fd97d305",
X"527951ff",
X"9dcb3f80",
X"d13dfdec",
X"055480fd",
X"5383e7f8",
X"527951ff",
X"9d833f7b",
X"81195956",
X"7580fc24",
X"83387858",
X"77882c55",
X"7483e8f5",
X"347783e8",
X"f6347583",
X"e8f73481",
X"805980cc",
X"3983eaa8",
X"08578378",
X"259b3883",
X"ea843383",
X"ea853371",
X"882b07fc",
X"1a712979",
X"05838005",
X"5951598d",
X"39778180",
X"2917ff80",
X"05578180",
X"59765279",
X"51ff9cd9",
X"3f80d13d",
X"fdec0554",
X"785383e7",
X"f8527951",
X"ff9c923f",
X"7851f6bf",
X"3fc5a13f",
X"c3da3f8b",
X"3983e9f8",
X"08810583",
X"e9f80c80",
X"d13d0d04",
X"f6e03ffc",
X"39fc3d0d",
X"76787184",
X"2983ea98",
X"05700851",
X"53535370",
X"9e3880ce",
X"723480cf",
X"0b811334",
X"80ce0b82",
X"133480c5",
X"0b831334",
X"70841334",
X"80e73983",
X"eab01333",
X"5480d272",
X"3473822a",
X"70810651",
X"5180cf53",
X"70843880",
X"d7537281",
X"1334a00b",
X"82133473",
X"83065170",
X"812e9e38",
X"70812488",
X"3870802e",
X"8f389f39",
X"70822e92",
X"3870832e",
X"92389339",
X"80d8558e",
X"3980d355",
X"893980cd",
X"55843980",
X"c4557483",
X"133480c4",
X"0b841334",
X"800b8513",
X"34863d0d",
X"0483e7f0",
X"0883e080",
X"0c04803d",
X"0d83e7f0",
X"08842980",
X"fdb40570",
X"0883e080",
X"0c51823d",
X"0d04fc3d",
X"0d767853",
X"54815380",
X"55873971",
X"10731054",
X"52737226",
X"5172802e",
X"a7387080",
X"2e863871",
X"8025e838",
X"72802e98",
X"38717426",
X"89387372",
X"31757407",
X"56547281",
X"2a72812a",
X"5353e539",
X"73517883",
X"38745170",
X"83e0800c",
X"863d0d04",
X"fe3d0d80",
X"53755274",
X"51ffa33f",
X"843d0d04",
X"fe3d0d81",
X"53755274",
X"51ff933f",
X"843d0d04",
X"fb3d0d77",
X"79555580",
X"56747625",
X"86387430",
X"55815673",
X"80258838",
X"73307681",
X"32575480",
X"53735274",
X"51fee73f",
X"83e08008",
X"5475802e",
X"873883e0",
X"80083054",
X"7383e080",
X"0c873d0d",
X"04fa3d0d",
X"787a5755",
X"80577477",
X"25863874",
X"30558157",
X"759f2c54",
X"81537574",
X"32743152",
X"7451feaa",
X"3f83e080",
X"08547680",
X"2e873883",
X"e0800830",
X"547383e0",
X"800c883d",
X"0d04fd3d",
X"0d755480",
X"740c800b",
X"84150c80",
X"0b88150c",
X"800b8c15",
X"0c87a680",
X"337081ff",
X"06707184",
X"2a065151",
X"51dae63f",
X"70812a81",
X"32718132",
X"71810671",
X"81063184",
X"170c5353",
X"70832a81",
X"3271822a",
X"81327081",
X"06727131",
X"770c5152",
X"5287a090",
X"3387a091",
X"337081ff",
X"06707306",
X"81328106",
X"88180c51",
X"525283e0",
X"8008802e",
X"80c23883",
X"e0800881",
X"2a708106",
X"83e08008",
X"81063184",
X"160c5183",
X"e0800883",
X"2a83e080",
X"08822a71",
X"81067181",
X"0631760c",
X"525283e0",
X"8008842a",
X"81068815",
X"0c83e080",
X"08852a81",
X"068c150c",
X"853d0d04",
X"fe3d0d74",
X"76545271",
X"51febb3f",
X"72812ea2",
X"38817326",
X"8d387282",
X"2ea83872",
X"832e9c38",
X"e6397108",
X"e2388412",
X"08dd3888",
X"1208d838",
X"a5398812",
X"08812e9e",
X"38913988",
X"1208812e",
X"95387108",
X"91388412",
X"088c388c",
X"1208812e",
X"098106ff",
X"b238843d",
X"0d040000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002b98",
X"00002bd9",
X"00002bfb",
X"00002c1d",
X"00002c43",
X"00002c43",
X"00002c43",
X"00002c43",
X"00002cb4",
X"00002d05",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"43505520",
X"54757262",
X"6f3a2564",
X"78000000",
X"44726976",
X"65205475",
X"72626f3a",
X"25730000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"66726565",
X"7a65722e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"4d454d00",
X"5374616e",
X"64617264",
X"00000000",
X"46617374",
X"28362900",
X"46617374",
X"28352900",
X"46617374",
X"28342900",
X"46617374",
X"28332900",
X"46617374",
X"28322900",
X"46617374",
X"28312900",
X"46617374",
X"28302900",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00003bf8",
X"00003bfc",
X"00003c04",
X"00003c10",
X"00003c1c",
X"00003c28",
X"00003c34",
X"00003c38",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00000028",
X"00000006",
X"00000005",
X"00000004",
X"00000003",
X"00000002",
X"00000001",
X"00000000",
X"00003cdc",
X"00003ce8",
X"00003cf0",
X"00003cf8",
X"00003d00",
X"00003d08",
X"00003d10",
X"00003d18",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
