
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81ca",
X"a0738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81d1",
X"b40c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757581c4",
X"cd2d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7581c2e1",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80ddf304",
X"fd3d0d75",
X"705254ae",
X"a43f83c0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"c0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83c0",
X"8008732e",
X"a13883c0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183c0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83c2d008",
X"248a38b4",
X"f93fff0b",
X"83c2d00c",
X"800b83c0",
X"800c04ff",
X"3d0d7352",
X"83c0ac08",
X"722e8d38",
X"d93f7151",
X"96993f71",
X"83c0ac0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"558154bc",
X"15088191",
X"387451cf",
X"3f795880",
X"7a2580f7",
X"3883c380",
X"0870892a",
X"5783ff06",
X"78848072",
X"31565657",
X"73782583",
X"38735575",
X"83c2d008",
X"2e8438ff",
X"893f83c2",
X"d0088025",
X"a6387589",
X"2b5198dc",
X"3f83c380",
X"088f3dfc",
X"11555c54",
X"8152f81b",
X"5196c63f",
X"761483c3",
X"800c7583",
X"c2d00c74",
X"53765278",
X"51b3aa3f",
X"83c08008",
X"83c38008",
X"1683c380",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8b3861",
X"7a710c54",
X"75547580",
X"2e833881",
X"547383c0",
X"800c8e3d",
X"0d04fc3d",
X"0dfe9b3f",
X"7651feaf",
X"3f863dfc",
X"05537852",
X"775195e9",
X"3f797571",
X"0c5483c0",
X"80085483",
X"c0800880",
X"2e833881",
X"547383c0",
X"800c863d",
X"0d04fe3d",
X"0d7583c2",
X"d0085353",
X"80722489",
X"3871732e",
X"8438fdd6",
X"3f7451fd",
X"ea3f7251",
X"97ae3f83",
X"c0800852",
X"83c08008",
X"802e8338",
X"81527183",
X"c0800c84",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"c0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"c0800c51",
X"823d0d04",
X"80c40b83",
X"c0800c04",
X"fd3d0d75",
X"77715470",
X"535553a9",
X"fc3f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfceb3f",
X"735193ab",
X"3f7383c0",
X"ac0c83c0",
X"80085383",
X"c0800880",
X"2e833881",
X"537283c0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcbf3f",
X"72802ea5",
X"38bc1308",
X"527351a9",
X"863f83c0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"c0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83c0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83c2d0",
X"0c7483c0",
X"b00c7583",
X"c2cc0caf",
X"de3f83c0",
X"800881ff",
X"06528153",
X"71993883",
X"c2e8518e",
X"943f83c0",
X"80085283",
X"c0800880",
X"2e833872",
X"52715372",
X"83c0800c",
X"843d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"51a6f73f",
X"83c08008",
X"557483c0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"c0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283c2cc",
X"085181b1",
X"9e3f83c0",
X"800857f9",
X"e13f7952",
X"83c2d451",
X"95b73f83",
X"c0800854",
X"805383c0",
X"8008732e",
X"09810682",
X"833883c0",
X"b0080b0b",
X"81cfbc53",
X"705256a6",
X"b43f0b0b",
X"81cfbc52",
X"80c01651",
X"a6a73f75",
X"bc170c73",
X"82c0170c",
X"810b82c4",
X"170c810b",
X"82c8170c",
X"7382cc17",
X"0cff1782",
X"d0175557",
X"81913983",
X"c0bc3370",
X"822a7081",
X"06515455",
X"72818038",
X"74812a81",
X"06587780",
X"f6387484",
X"2a810682",
X"c4150c83",
X"c0bc3381",
X"0682c815",
X"0c795273",
X"51a5ce3f",
X"7351a5e5",
X"3f83c080",
X"081453af",
X"73708105",
X"553472bc",
X"150c83c0",
X"bd527251",
X"a5af3f83",
X"c0b40882",
X"c0150c83",
X"c0ca5280",
X"c01451a5",
X"9c3f7880",
X"2e8d3873",
X"51782d83",
X"c0800880",
X"2e993877",
X"82cc150c",
X"75802e86",
X"387382cc",
X"170c7382",
X"d015ff19",
X"59555676",
X"802e9b38",
X"83c0b452",
X"83c2d451",
X"94ad3f83",
X"c080088a",
X"3883c0bd",
X"335372fe",
X"d2387880",
X"2e893883",
X"c0b00851",
X"fcb83f83",
X"c0b00853",
X"7283c080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb53f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f690",
X"3f83c080",
X"08745387",
X"3d705355",
X"55f6b03f",
X"f7903f73",
X"51d33f63",
X"53745283",
X"c0800851",
X"fab83f92",
X"3d0d0471",
X"83c0800c",
X"0480c012",
X"83c0800c",
X"04803d0d",
X"7282c011",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"c0800c51",
X"823d0d04",
X"f93d0d79",
X"83c09008",
X"57578177",
X"27819638",
X"76881708",
X"27818e38",
X"75335574",
X"822e8938",
X"74832eb3",
X"3880fe39",
X"74547610",
X"83fe0653",
X"76882a8c",
X"17080552",
X"893dfc05",
X"51aa8c3f",
X"83c08008",
X"80df3802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d13984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"51a9dc3f",
X"83c08008",
X"b038029f",
X"05330284",
X"059e0533",
X"71982b71",
X"902b0702",
X"8c059d05",
X"3370882b",
X"72078d3d",
X"337180ff",
X"fffe8006",
X"07515253",
X"57585683",
X"39815574",
X"83c0800c",
X"893d0d04",
X"fb3d0d83",
X"c09008fe",
X"19881208",
X"fe055556",
X"54805674",
X"73278d38",
X"82143375",
X"71299416",
X"08055753",
X"7583c080",
X"0c873d0d",
X"04fc3d0d",
X"7652800b",
X"83c09008",
X"70335152",
X"5370832e",
X"09810691",
X"38951233",
X"94133371",
X"982b7190",
X"2b075555",
X"519b1233",
X"9a133371",
X"882b0774",
X"0783c080",
X"0c55863d",
X"0d04fc3d",
X"0d7683c0",
X"90085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"fed63f83",
X"c0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183c080",
X"0c863d0d",
X"04fa3d0d",
X"7883c090",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fcb13f",
X"81527183",
X"c0800827",
X"a8388352",
X"83c08008",
X"88170827",
X"9c3883c0",
X"80088c16",
X"0c83c080",
X"0851fdbc",
X"3f83c080",
X"0890160c",
X"73752380",
X"527183c0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585e5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"9f269138",
X"7a51fdd2",
X"3f83c080",
X"0856807d",
X"34838139",
X"933d841c",
X"08705859",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"3880705a",
X"5c887f08",
X"5f5a7b81",
X"1d7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535e57",
X"557480e7",
X"3876ae2e",
X"09810683",
X"38815578",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675bb",
X"3888598b",
X"5affab39",
X"76982b55",
X"74802587",
X"3881c9b0",
X"173357ff",
X"9f175574",
X"99268938",
X"e0177081",
X"ff065855",
X"78811a70",
X"81ff0672",
X"1b535b57",
X"55767534",
X"fef8397b",
X"1e7f0c80",
X"5576a026",
X"83388155",
X"748b1934",
X"7a51fc82",
X"3f83c080",
X"0880f538",
X"a0547a22",
X"70852b83",
X"e0065455",
X"901b0852",
X"7c51a497",
X"3f83c080",
X"085783c0",
X"80088181",
X"387c3355",
X"74802e80",
X"f4388b1d",
X"3370832a",
X"70810651",
X"565674b4",
X"388b7d84",
X"1d0883c0",
X"8008595b",
X"5b58ff18",
X"5877ff2e",
X"9a387970",
X"81055b33",
X"79708105",
X"5b337171",
X"31525656",
X"75802ee2",
X"38863975",
X"802e9638",
X"7a51fbe5",
X"3fff8639",
X"83c08008",
X"5683c080",
X"08b63883",
X"39765684",
X"1b088b11",
X"33515574",
X"a7388b1d",
X"3370842a",
X"70810651",
X"56567489",
X"38835694",
X"39815690",
X"397c51fa",
X"943f83c0",
X"8008881c",
X"0cfd8139",
X"7583c080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"51a2dc3f",
X"835683c0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"51a2b03f",
X"83c08008",
X"98388117",
X"33773371",
X"882b0783",
X"c0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"7651a287",
X"3f83c080",
X"08983881",
X"17337733",
X"71882b07",
X"83c08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583c080",
X"0c8a3d0d",
X"04eb3d0d",
X"675a800b",
X"83c0900c",
X"a1a93f83",
X"c0800881",
X"06558256",
X"7483ef38",
X"7475538f",
X"3d705357",
X"59feca3f",
X"83c08008",
X"81ff0657",
X"76812e09",
X"810680d4",
X"38905483",
X"be537452",
X"7551a19b",
X"3f83c080",
X"0880c938",
X"8f3d3355",
X"74802e80",
X"c93802bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"33710770",
X"587b575e",
X"525e5759",
X"57fdee3f",
X"83c08008",
X"81ff0657",
X"76832e09",
X"81068638",
X"815682f2",
X"3976802e",
X"86388656",
X"82e839a4",
X"548d5378",
X"527551a0",
X"b23f8156",
X"83c08008",
X"82d43802",
X"be053302",
X"8405bd05",
X"3371882b",
X"07595d77",
X"ab380280",
X"ce053302",
X"840580cd",
X"05337198",
X"2b71902b",
X"07973d33",
X"70882b72",
X"07029405",
X"80cb0533",
X"71075452",
X"5e575956",
X"02b70533",
X"78712902",
X"8805b605",
X"33028c05",
X"b5053371",
X"882b0770",
X"1d707f8c",
X"050c5f59",
X"57595d8e",
X"3d33821b",
X"3402b905",
X"33903d33",
X"71882b07",
X"5a5c7884",
X"1b2302bb",
X"05330284",
X"05ba0533",
X"71882b07",
X"565c74ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"07515253",
X"575e5c74",
X"76317831",
X"79842a90",
X"3d335471",
X"71315356",
X"5681a283",
X"3f83c080",
X"08820570",
X"881c0c83",
X"c08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83c0900c",
X"80567583",
X"c0800c97",
X"3d0d04e9",
X"3d0d83c0",
X"90085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e53f83c0",
X"80085483",
X"c0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f489",
X"3f83c080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383c080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83c09008",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0e93f",
X"83c08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"833f83c0",
X"80085583",
X"c0800880",
X"2eff8938",
X"83c08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"519ad83f",
X"83c08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83c0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83c09008",
X"55568555",
X"73802e81",
X"e3388114",
X"33810653",
X"84557280",
X"2e81d538",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b9388214",
X"3370892b",
X"56537680",
X"2eb73874",
X"52ff1651",
X"819d843f",
X"83c08008",
X"ff187654",
X"70535853",
X"819cf43f",
X"83c08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed63f83",
X"c0800853",
X"810b83c0",
X"8008278b",
X"38881408",
X"83c08008",
X"26883880",
X"0b811534",
X"b03983c0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc53f",
X"83c08008",
X"8c3883c0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683c0",
X"800805a8",
X"150c8055",
X"7483c080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83c09008",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1cf3f",
X"83c08008",
X"5583c080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef5",
X"3f83c080",
X"0888170c",
X"7551efa6",
X"3f83c080",
X"08557483",
X"c0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683c0",
X"9008802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f53f83c0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"96e13f83",
X"c0800841",
X"83c08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"eddf3f83",
X"c0800841",
X"83c08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"8e833f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f03f83c0",
X"80088332",
X"70307072",
X"079f2c83",
X"c0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"8c8f3f75",
X"83c0800c",
X"9e3d0d04",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"7751e0d2",
X"3f83c080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3381d1bc",
X"0b81d1bc",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"527751e0",
X"813f83c0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583c0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"558b963f",
X"83c08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"8114518a",
X"ae3f83c0",
X"80083070",
X"83c08008",
X"07802583",
X"c0800c53",
X"863d0d04",
X"fc3d0d76",
X"705255e6",
X"ee3f83c0",
X"80085481",
X"5383c080",
X"0880c138",
X"7451e6b1",
X"3f83c080",
X"0881cfcc",
X"5383c080",
X"085253ff",
X"913f83c0",
X"8008a138",
X"81cfd052",
X"7251ff82",
X"3f83c080",
X"08923881",
X"cfd45272",
X"51fef33f",
X"83c08008",
X"802e8338",
X"81547353",
X"7283c080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"e68d3f81",
X"5383c080",
X"08983873",
X"51e5d63f",
X"83c39808",
X"5283c080",
X"0851feba",
X"3f83c080",
X"08537283",
X"c0800c85",
X"3d0d04df",
X"3d0da43d",
X"0870525e",
X"dbfb3f83",
X"c0800833",
X"953d5654",
X"73963881",
X"d2d85274",
X"51898e3f",
X"9a397d52",
X"7851defc",
X"3f84cd39",
X"7d51dbe1",
X"3f83c080",
X"08527451",
X"db913f80",
X"43804280",
X"41804083",
X"c3a00852",
X"943d7052",
X"5de1e43f",
X"83c08008",
X"59800b83",
X"c0800855",
X"5b83c080",
X"087b2e94",
X"38811b74",
X"525be4e6",
X"3f83c080",
X"085483c0",
X"8008ee38",
X"805aff5f",
X"7909709f",
X"2c7b065b",
X"547a7a24",
X"8438ff1b",
X"5af61a70",
X"09709f2c",
X"72067bff",
X"125a5a52",
X"55558075",
X"25953876",
X"51e4ab3f",
X"83c08008",
X"76ff1858",
X"55577380",
X"24ed3874",
X"7f2e8638",
X"a0c73f74",
X"5f78ff1b",
X"70585d58",
X"807a2595",
X"387751e4",
X"813f83c0",
X"800876ff",
X"18585558",
X"738024ed",
X"38800b83",
X"c7d00c80",
X"0b83c894",
X"0c81cfd8",
X"518d913f",
X"81800b83",
X"c8940c81",
X"cfe0518d",
X"833fa80b",
X"83c7d00c",
X"76802e80",
X"e43883c7",
X"d0087779",
X"32703070",
X"72078025",
X"70872b83",
X"c8940c51",
X"56785356",
X"56e3b83f",
X"83c08008",
X"802e8838",
X"81cfe851",
X"8cca3f76",
X"51e2fa3f",
X"83c08008",
X"5281d0fc",
X"518cb93f",
X"7651e382",
X"3f83c080",
X"0883c7d0",
X"08555775",
X"74258638",
X"a81656f7",
X"397583c7",
X"d00c86f0",
X"7624ff98",
X"3887980b",
X"83c7d00c",
X"77802eb1",
X"387751e2",
X"b83f83c0",
X"80087852",
X"55e2d83f",
X"81cff054",
X"83c08008",
X"8d388739",
X"80763481",
X"ce3981cf",
X"ec547453",
X"735281cf",
X"c0518bd8",
X"3f805481",
X"cfc8518b",
X"cf3f8114",
X"5473a82e",
X"098106ef",
X"38868da0",
X"519cbb3f",
X"8052903d",
X"705257af",
X"ee3f8352",
X"7651afe7",
X"3f62818f",
X"3861802e",
X"80fb387b",
X"5473ff2e",
X"96387880",
X"2e818938",
X"7851e1de",
X"3f83c080",
X"08ff1555",
X"59e73978",
X"802e80f4",
X"387851e1",
X"da3f83c0",
X"8008802e",
X"fc903878",
X"51e1a23f",
X"83c08008",
X"5281cfbc",
X"5183e33f",
X"83c08008",
X"a3387c51",
X"859b3f83",
X"c0800855",
X"74ff1656",
X"54807425",
X"ae38741d",
X"70335556",
X"73af2efe",
X"cf38e939",
X"7851e0e3",
X"3f83c080",
X"08527c51",
X"84d33f8f",
X"397f8829",
X"6010057a",
X"0561055a",
X"fc923962",
X"802efbd3",
X"38805276",
X"51aec83f",
X"a33d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"842a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"a80b9088",
X"b834b80b",
X"9088b834",
X"7083c080",
X"0c823d0d",
X"04803d0d",
X"9088b833",
X"7081ff06",
X"70852a81",
X"32708106",
X"51515151",
X"70802e8d",
X"38980b90",
X"88b834b8",
X"0b9088b8",
X"347083c0",
X"800c823d",
X"0d04930b",
X"9088bc34",
X"ff0b9088",
X"a83404ff",
X"3d0d028f",
X"05335280",
X"0b9088bc",
X"348a519a",
X"853fdf3f",
X"80f80b90",
X"88a03480",
X"0b908888",
X"34fa1252",
X"71908880",
X"34800b90",
X"88983471",
X"90889034",
X"9088b852",
X"807234b8",
X"7234833d",
X"0d04803d",
X"0d028b05",
X"33517090",
X"88b434fe",
X"bf3f83c0",
X"8008802e",
X"f638823d",
X"0d04803d",
X"0d8439a7",
X"943ffed9",
X"3f83c080",
X"08802ef3",
X"389088b4",
X"337081ff",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0da30b90",
X"88bc34ff",
X"0b9088a8",
X"349088b8",
X"51a87134",
X"b8713482",
X"3d0d0480",
X"3d0d9088",
X"bc337081",
X"c0067030",
X"70802583",
X"c0800c51",
X"5151823d",
X"0d04803d",
X"0d9088b8",
X"337081ff",
X"0670832a",
X"81327081",
X"06515151",
X"5170802e",
X"e838b00b",
X"9088b834",
X"b80b9088",
X"b834823d",
X"0d04803d",
X"0d9080ac",
X"08810683",
X"c0800c82",
X"3d0d04fd",
X"3d0d7577",
X"54548073",
X"25943873",
X"70810555",
X"335281cf",
X"f4518788",
X"3fff1353",
X"e939853d",
X"0d04fd3d",
X"0d757753",
X"54733351",
X"70893871",
X"33517080",
X"2ea13873",
X"33723352",
X"53727127",
X"8538ff51",
X"94397073",
X"27853881",
X"518b3981",
X"14811353",
X"54d33980",
X"517083c0",
X"800c853d",
X"0d04fd3d",
X"0d757754",
X"54723370",
X"81ff0652",
X"5270802e",
X"a3387181",
X"ff068114",
X"ffbf1253",
X"54527099",
X"268938a0",
X"127081ff",
X"06535171",
X"74708105",
X"5634d239",
X"80743485",
X"3d0d04ff",
X"bd3d0d80",
X"c63d0852",
X"a53d7052",
X"54ffb33f",
X"80c73d08",
X"52853d70",
X"5253ffa6",
X"3f725273",
X"51fedf3f",
X"80c53d0d",
X"04fe3d0d",
X"74765353",
X"71708105",
X"53335170",
X"73708105",
X"553470f0",
X"38843d0d",
X"04fe3d0d",
X"74528072",
X"33525370",
X"732e8d38",
X"81128114",
X"71335354",
X"5270f538",
X"7283c080",
X"0c843d0d",
X"04f63d0d",
X"7c7e6062",
X"5a5d5b56",
X"80598155",
X"8539747a",
X"29557452",
X"75518189",
X"da3f83c0",
X"80087a27",
X"ed387480",
X"2e80e038",
X"74527551",
X"8189c43f",
X"83c08008",
X"75537652",
X"548189ea",
X"3f83c080",
X"087a5375",
X"52568189",
X"aa3f83c0",
X"80087930",
X"707b079f",
X"2a707780",
X"24075151",
X"54557287",
X"3883c080",
X"08c23876",
X"8118b016",
X"55585889",
X"74258b38",
X"b714537a",
X"853880d7",
X"14537278",
X"34811959",
X"ff9c3980",
X"77348c3d",
X"0d04f73d",
X"0d7b7d7f",
X"62029005",
X"bb053357",
X"59565a5a",
X"b0587283",
X"38a05875",
X"70708105",
X"52337159",
X"54559039",
X"8074258e",
X"38ff1477",
X"70810559",
X"33545472",
X"ef3873ff",
X"15555380",
X"73258938",
X"77527951",
X"782def39",
X"75337557",
X"5372802e",
X"90387252",
X"7951782d",
X"75708105",
X"573353ed",
X"398b3d0d",
X"04ee3d0d",
X"64666969",
X"70708105",
X"52335b4a",
X"5c5e5e76",
X"802e82f9",
X"3876a52e",
X"09810682",
X"e0388070",
X"41677070",
X"81055233",
X"714a5957",
X"5f76b02e",
X"0981068c",
X"38757081",
X"05573376",
X"4857815f",
X"d0175675",
X"892680da",
X"3876675c",
X"59805c93",
X"39778a24",
X"80c3387b",
X"8a29187b",
X"7081055d",
X"335a5cd0",
X"197081ff",
X"06585889",
X"7727a438",
X"ff9f1970",
X"81ff06ff",
X"a91b5a51",
X"56857627",
X"9238ffbf",
X"197081ff",
X"06515675",
X"85268a38",
X"c9195877",
X"8025ffb9",
X"387a477b",
X"407881ff",
X"06577680",
X"e42e80e5",
X"387680e4",
X"24a73876",
X"80d82e81",
X"86387680",
X"d8249038",
X"76802e81",
X"cc3876a5",
X"2e81b638",
X"81b93976",
X"80e32e81",
X"8c3881af",
X"397680f5",
X"2e9b3876",
X"80f5248b",
X"387680f3",
X"2e818138",
X"81993976",
X"80f82e80",
X"ca38818f",
X"39913d70",
X"55578053",
X"8a527984",
X"1b710853",
X"5b56fbfd",
X"3f7655ab",
X"3979841b",
X"7108943d",
X"705b5b52",
X"5b567580",
X"258c3875",
X"3056ad78",
X"340280c1",
X"05577654",
X"80538a52",
X"7551fbd1",
X"3f77557e",
X"54b83991",
X"3d705577",
X"80d83270",
X"30708025",
X"56515856",
X"90527984",
X"1b710853",
X"5b57fbad",
X"3f7555db",
X"3979841b",
X"83123354",
X"5b569839",
X"79841b71",
X"08575b56",
X"80547f53",
X"7c527d51",
X"fc9c3f87",
X"3976527d",
X"517c2d66",
X"70335881",
X"0547fd83",
X"39943d0d",
X"047283c0",
X"940c7183",
X"c0980c04",
X"fb3d0d88",
X"3d707084",
X"05520857",
X"54755383",
X"c0940852",
X"83c09808",
X"51fcc63f",
X"873d0d04",
X"ff3d0d73",
X"70085351",
X"02930533",
X"72347008",
X"8105710c",
X"833d0d04",
X"fc3d0d87",
X"3d881155",
X"7854bdbc",
X"5351fc99",
X"3f805287",
X"3d51d13f",
X"863d0d04",
X"fc3d0d76",
X"557483c3",
X"ac082eaf",
X"38805374",
X"5187c13f",
X"83c08008",
X"81ff06ff",
X"147081ff",
X"06723070",
X"9f2a5152",
X"55535472",
X"802e8438",
X"71dd3873",
X"fe387483",
X"c3ac0c86",
X"3d0d04ff",
X"3d0dff0b",
X"83c3ac0c",
X"84a53f81",
X"5187853f",
X"83c08008",
X"81ff0652",
X"71ee3881",
X"d33f7183",
X"c0800c83",
X"3d0d04fc",
X"3d0d7602",
X"8405a205",
X"22028805",
X"a605227a",
X"54555555",
X"ff823f72",
X"802ea038",
X"83c3c014",
X"33757081",
X"05573481",
X"147083ff",
X"ff06ff15",
X"7083ffff",
X"06565255",
X"52dd3980",
X"0b83c080",
X"0c863d0d",
X"04fc3d0d",
X"76787a11",
X"56535580",
X"5371742e",
X"93387215",
X"51703383",
X"c3c01334",
X"81128114",
X"5452ea39",
X"800b83c0",
X"800c863d",
X"0d04fd3d",
X"0d905483",
X"c3ac0851",
X"86f43f83",
X"c0800881",
X"ff06ff15",
X"71307130",
X"7073079f",
X"2a729f2a",
X"06525552",
X"555372db",
X"38853d0d",
X"04803d0d",
X"83c3b808",
X"1083c3b0",
X"08079080",
X"a80c823d",
X"0d04800b",
X"83c3b80c",
X"e43f0481",
X"0b83c3b8",
X"0cdb3f04",
X"ed3f0471",
X"83c3b40c",
X"04803d0d",
X"8051f43f",
X"810b83c3",
X"b80c810b",
X"83c3b00c",
X"ffbb3f82",
X"3d0d0480",
X"3d0d7230",
X"70740780",
X"2583c3b0",
X"0c51ffa5",
X"3f823d0d",
X"04803d0d",
X"028b0533",
X"9080a40c",
X"9080a808",
X"70810651",
X"5170f538",
X"9080a408",
X"7081ff06",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"81ff51d1",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"823d0d04",
X"803d0d73",
X"902b7307",
X"9080b40c",
X"823d0d04",
X"04fb3d0d",
X"78028405",
X"9f053370",
X"982b5557",
X"55728025",
X"9b387580",
X"ff065680",
X"5280f751",
X"e03f83c0",
X"800881ff",
X"06547381",
X"2680ff38",
X"8051fee7",
X"3fffa23f",
X"8151fedf",
X"3fff9a3f",
X"7551feed",
X"3f74982a",
X"51fee63f",
X"74902a70",
X"81ff0652",
X"53feda3f",
X"74882a70",
X"81ff0652",
X"53fece3f",
X"7481ff06",
X"51fec63f",
X"81557580",
X"c02e0981",
X"06863881",
X"95558d39",
X"7580c82e",
X"09810684",
X"38818755",
X"7451fea5",
X"3f8a55fe",
X"c83f83c0",
X"800881ff",
X"0670982b",
X"54547280",
X"258c38ff",
X"157081ff",
X"06565374",
X"e2387383",
X"c0800c87",
X"3d0d04fa",
X"3d0dfdc5",
X"3f8051fd",
X"da3f8a54",
X"fe933fff",
X"147081ff",
X"06555373",
X"f3387374",
X"535580c0",
X"51fea63f",
X"83c08008",
X"81ff0654",
X"73812e09",
X"8106829f",
X"3883aa52",
X"80c851fe",
X"8c3f83c0",
X"800881ff",
X"06537281",
X"2e098106",
X"81a83874",
X"54873d74",
X"115456fd",
X"c83f83c0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e5",
X"38029a05",
X"33537281",
X"2e098106",
X"81d93802",
X"9b053353",
X"80ce9054",
X"7281aa2e",
X"8d3881c7",
X"3980e451",
X"8aa83fff",
X"14547380",
X"2e81b838",
X"820a5281",
X"e951fda5",
X"3f83c080",
X"0881ff06",
X"5372de38",
X"725280fa",
X"51fd923f",
X"83c08008",
X"81ff0653",
X"72819038",
X"72547316",
X"53fcd63f",
X"83c08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e83887",
X"3d337086",
X"2a708106",
X"5154548c",
X"557280e3",
X"38845580",
X"de397452",
X"81e951fc",
X"cc3f83c0",
X"800881ff",
X"06538255",
X"81e95681",
X"73278638",
X"735580c1",
X"5680ce90",
X"548a3980",
X"e451899a",
X"3fff1454",
X"73802ea9",
X"38805275",
X"51fc9a3f",
X"83c08008",
X"81ff0653",
X"72e13884",
X"805280d0",
X"51fc863f",
X"83c08008",
X"81ff0653",
X"72802e83",
X"38805574",
X"83c3bc34",
X"8051fb87",
X"3ffbc23f",
X"883d0d04",
X"fb3d0d77",
X"54800b83",
X"c3bc3370",
X"832a7081",
X"06515557",
X"5572752e",
X"09810685",
X"3873892b",
X"54735280",
X"d151fbbd",
X"3f83c080",
X"0881ff06",
X"5372bd38",
X"82b8c054",
X"fb833f83",
X"c0800881",
X"ff065372",
X"81ff2e09",
X"81068938",
X"ff145473",
X"e7389f39",
X"7281fe2e",
X"09810696",
X"3883c7c0",
X"5283c3c0",
X"51faed3f",
X"fad33ffa",
X"d03f8339",
X"81558051",
X"fa893ffa",
X"c43f7481",
X"ff0683c0",
X"800c873d",
X"0d04fb3d",
X"0d7783c3",
X"c0565481",
X"51f9ec3f",
X"83c3bc33",
X"70832a70",
X"81065154",
X"56728538",
X"73892b54",
X"735280d8",
X"51fab63f",
X"83c08008",
X"81ff0653",
X"7280e438",
X"81ff51f9",
X"d43f81fe",
X"51f9ce3f",
X"84805374",
X"70810556",
X"3351f9c1",
X"3fff1370",
X"83ffff06",
X"515372eb",
X"387251f9",
X"b03f7251",
X"f9ab3ff9",
X"d03f83c0",
X"80089f06",
X"53a78854",
X"72852e8c",
X"38993980",
X"e45186d2",
X"3fff1454",
X"f9b33f83",
X"c0800881",
X"ff2e8438",
X"73e93880",
X"51f8e43f",
X"f99f3f80",
X"0b83c080",
X"0c873d0d",
X"047183c7",
X"c40c8880",
X"800b83c7",
X"c00c8480",
X"800b83c7",
X"c80c04f0",
X"3d0d8380",
X"805683c7",
X"c4081683",
X"c7c00817",
X"56547433",
X"743483c7",
X"c8081654",
X"80743481",
X"16567583",
X"80a02e09",
X"8106db38",
X"83d08056",
X"83c7c408",
X"1683c7c0",
X"08175654",
X"74337434",
X"83c7c808",
X"16548074",
X"34811656",
X"7583d090",
X"2e098106",
X"db3883a8",
X"805683c7",
X"c4081683",
X"c7c00817",
X"56547433",
X"743483c7",
X"c8081654",
X"80743481",
X"16567583",
X"a8902e09",
X"8106db38",
X"805683c7",
X"c4081683",
X"c7c80817",
X"55557333",
X"75348116",
X"56758180",
X"802e0981",
X"06e43886",
X"f83f893d",
X"58a25381",
X"cbb05277",
X"5180ffce",
X"3f80578c",
X"805683c7",
X"c8081677",
X"19555573",
X"33753481",
X"16811858",
X"5676a22e",
X"098106e6",
X"38860b87",
X"a8833480",
X"0b87a882",
X"34800b87",
X"809a34af",
X"0b878096",
X"34bf0b87",
X"80973480",
X"0b878098",
X"349f0b87",
X"80993480",
X"0b87809b",
X"34f80b87",
X"a8893476",
X"87a88034",
X"820b87d0",
X"8f34820b",
X"87a88134",
X"923d0d04",
X"fe3d0d80",
X"5383c7c8",
X"081383c7",
X"c4081452",
X"52703372",
X"34811353",
X"72818080",
X"2e098106",
X"e4388380",
X"805383c7",
X"c8081383",
X"c7c40814",
X"52527033",
X"72348113",
X"53728380",
X"a02e0981",
X"06e43883",
X"d0805383",
X"c7c80813",
X"83c7c408",
X"14525270",
X"33723481",
X"13537283",
X"d0902e09",
X"8106e438",
X"83a88053",
X"83c7c808",
X"1383c7c4",
X"08145252",
X"70337234",
X"81135372",
X"83a8902e",
X"098106e4",
X"38843d0d",
X"04803d0d",
X"90809008",
X"810683c0",
X"800c823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087081",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fd0676",
X"1007720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870822c",
X"bf0683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe830676",
X"822b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087088",
X"2c870683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f1ff06",
X"76882b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"912cbf06",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fc87",
X"ffff0676",
X"912b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087099",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70ffbf0a",
X"0676992b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90808008",
X"70882c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"0870892c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708a",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8b2c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708c2cbf",
X"0683c080",
X"0c51823d",
X"0d04fe3d",
X"0d7481e6",
X"29872a90",
X"80a00c84",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70810554",
X"34ff1151",
X"f039843d",
X"0d04fe3d",
X"0d7575ff",
X"19535353",
X"70ff2e8d",
X"38727270",
X"8405540c",
X"ff1151f0",
X"39843d0d",
X"04fe3d0d",
X"81808053",
X"80528880",
X"0a51ffb3",
X"3fa08053",
X"80528280",
X"0a51c73f",
X"843d0d04",
X"803d0d81",
X"51fcab3f",
X"72802e90",
X"388051fd",
X"ff3fce3f",
X"81d2b033",
X"51fdf53f",
X"8151fcbc",
X"3f8051fc",
X"b73f8051",
X"fc883f82",
X"3d0d04fd",
X"3d0d7552",
X"805480ff",
X"72258838",
X"810bff80",
X"135354ff",
X"bf125170",
X"99268638",
X"e01252b0",
X"39ff9f12",
X"51997127",
X"a738d012",
X"e0135451",
X"70892685",
X"38725298",
X"39728f26",
X"85387252",
X"8f3971ba",
X"2e098106",
X"85389a52",
X"83398052",
X"73802e85",
X"38818012",
X"527181ff",
X"0683c080",
X"0c853d0d",
X"04803d0d",
X"84d8c051",
X"80717081",
X"05533470",
X"84e0c02e",
X"098106f0",
X"38823d0d",
X"04fe3d0d",
X"02970533",
X"51fef43f",
X"83c08008",
X"81ff0683",
X"c7d00854",
X"52807324",
X"9b3883c8",
X"90081372",
X"83c89408",
X"07535371",
X"733483c7",
X"d0088105",
X"83c7d00c",
X"843d0d04",
X"fa3d0d82",
X"800a1b55",
X"8057883d",
X"fc055479",
X"53745278",
X"51ffbb9a",
X"3f883d0d",
X"04fe3d0d",
X"83c7e808",
X"527451c1",
X"fe3f83c0",
X"80088c38",
X"76537552",
X"83c7e808",
X"51c63f84",
X"3d0d04fe",
X"3d0d83c7",
X"e8085375",
X"527451ff",
X"bcbc3f83",
X"c080088d",
X"38775376",
X"5283c7e8",
X"0851ffa0",
X"3f843d0d",
X"04fd3d0d",
X"83c7e808",
X"51ffbbaf",
X"3f83c080",
X"0890802e",
X"098106ad",
X"38805483",
X"c1808053",
X"83c08008",
X"5283c7e8",
X"0851fef0",
X"3f87c180",
X"80143387",
X"c1908015",
X"34811454",
X"7390802e",
X"098106e9",
X"38853d0d",
X"0481cffc",
X"0b83c080",
X"0c04fc3d",
X"0d765473",
X"902e80ff",
X"38739024",
X"8e387384",
X"2e983873",
X"862ea638",
X"82b93973",
X"932e8195",
X"3873942e",
X"81cf3882",
X"aa398180",
X"80538280",
X"805283c7",
X"e40851fe",
X"8f3f82b5",
X"39805481",
X"80805380",
X"c0805283",
X"c7e40851",
X"fdfa3f82",
X"80805380",
X"c0805283",
X"c7e40851",
X"fdea3f84",
X"81808014",
X"338481c0",
X"80153484",
X"82808014",
X"338482c0",
X"80153481",
X"14547380",
X"c0802e09",
X"8106dc38",
X"81eb3982",
X"80805381",
X"80805283",
X"c7e40851",
X"fdb23f80",
X"54848280",
X"80143384",
X"81808015",
X"34811454",
X"73818080",
X"2e098106",
X"e83881bd",
X"39818080",
X"5380c080",
X"5283c7e4",
X"0851fd84",
X"3f805584",
X"81808015",
X"54733384",
X"81c08016",
X"34733384",
X"82808016",
X"34733384",
X"82c08016",
X"34811555",
X"7480c080",
X"2e098106",
X"d63880fd",
X"39818080",
X"53a08052",
X"83c7e408",
X"51fcc53f",
X"80558481",
X"80801554",
X"73338481",
X"a0801634",
X"73338481",
X"c0801634",
X"73338481",
X"e0801634",
X"73338482",
X"80801634",
X"73338482",
X"a0801634",
X"73338482",
X"c0801634",
X"73338482",
X"e0801634",
X"81155574",
X"a0802e09",
X"8106ffb6",
X"389f39fb",
X"9c3f800b",
X"83c7d00c",
X"800b83c8",
X"940c81d0",
X"8051e888",
X"3f81b78d",
X"c051f8fe",
X"3f863d0d",
X"04fc3d0d",
X"76705255",
X"ffbed03f",
X"83c08008",
X"54815383",
X"c0800880",
X"c2387451",
X"ffbe923f",
X"83c08008",
X"81d09c53",
X"83c08008",
X"5253d6f2",
X"3f83c080",
X"08a13881",
X"d0a05272",
X"51d6e33f",
X"83c08008",
X"923881d0",
X"a4527251",
X"d6d43f83",
X"c0800880",
X"2e833881",
X"54735372",
X"83c0800c",
X"863d0d04",
X"f13d0d80",
X"d5a10b83",
X"c3a00c83",
X"c7e40851",
X"d8813f83",
X"c7e40851",
X"ffb3fe3f",
X"ff0b81d0",
X"a05383c0",
X"80085256",
X"d6943f83",
X"c0800880",
X"2e9f3880",
X"58913ddc",
X"11555590",
X"53f01552",
X"83c7e408",
X"51ffb5da",
X"3f02b705",
X"335681a3",
X"3983c7e4",
X"0851ffb6",
X"b63f83c0",
X"80085783",
X"c0800882",
X"80802e09",
X"81068338",
X"845683c0",
X"80088180",
X"802e0981",
X"0680df38",
X"805b805a",
X"8059f995",
X"3f800b83",
X"c7d00c80",
X"0b83c894",
X"0c81d0a8",
X"51e6813f",
X"80d00b83",
X"c7d00c81",
X"d0b851e5",
X"f33f80f8",
X"0b83c7d0",
X"0c81d0cc",
X"51e5e53f",
X"758025a2",
X"38805289",
X"3d705255",
X"8a913f83",
X"5274518a",
X"8a3f7855",
X"74802583",
X"38905680",
X"7525dd38",
X"86567680",
X"c0802e09",
X"81068538",
X"93568c39",
X"76a0802e",
X"09810683",
X"38945675",
X"51faaf3f",
X"913d0d04",
X"f73d0d80",
X"59805880",
X"57807056",
X"56f88e3f",
X"800b83c7",
X"d00c800b",
X"83c8940c",
X"81d0e051",
X"e4fa3f81",
X"800b83c8",
X"940c81d0",
X"e451e4ec",
X"3f80d00b",
X"83c7d00c",
X"74307076",
X"07802570",
X"872b83c8",
X"940c5153",
X"f3b03f83",
X"c0800852",
X"81d0ec51",
X"e4c63f80",
X"f80b83c7",
X"d00c7481",
X"32703070",
X"72078025",
X"70872b83",
X"c8940c51",
X"5454f9ad",
X"3f83c080",
X"085281d0",
X"f851e49c",
X"3f81a00b",
X"83c7d00c",
X"74823270",
X"30707207",
X"80257087",
X"2b83c894",
X"0c515483",
X"c7e80852",
X"54ffb0f9",
X"3f83c080",
X"085281d1",
X"8051e3ec",
X"3f81c80b",
X"83c7d00c",
X"74833270",
X"30707207",
X"80257087",
X"2b83c894",
X"0c515483",
X"c7e40852",
X"54ffb0c9",
X"3f81d188",
X"5383c080",
X"08802e8f",
X"3883c7e4",
X"0851ffb0",
X"b43f83c0",
X"80085372",
X"5281d190",
X"51e3a53f",
X"81f00b83",
X"c7d00c74",
X"84327030",
X"70720780",
X"2570872b",
X"83c8940c",
X"515581d1",
X"985253e3",
X"833f868d",
X"a051f3fa",
X"3f805287",
X"3d705253",
X"87ad3f83",
X"52725187",
X"a63f7715",
X"55748025",
X"85388055",
X"90398475",
X"25853884",
X"55873974",
X"842681a0",
X"38748429",
X"81cbd405",
X"53720804",
X"f1a03f83",
X"c0800877",
X"55537381",
X"2e098106",
X"893883c0",
X"80081053",
X"903973ff",
X"2e098106",
X"883883c0",
X"8008812c",
X"53907325",
X"85389053",
X"88397280",
X"24833881",
X"537251f0",
X"fa3f80d4",
X"39f18c3f",
X"83c08008",
X"17537280",
X"25853880",
X"53883987",
X"73258338",
X"87537251",
X"f1863fb4",
X"39768638",
X"78802eac",
X"3883c39c",
X"0883c398",
X"0cade50b",
X"83c3a00c",
X"83c7e808",
X"51d2c03f",
X"f5ff3f90",
X"3978802e",
X"8b38faa0",
X"3f81538c",
X"39788738",
X"75802efc",
X"9c388053",
X"7283c080",
X"0c8b3d0d",
X"04ff3d0d",
X"83c88051",
X"80df863f",
X"83c7f051",
X"80defe3f",
X"f19f3f83",
X"c0800880",
X"2e863880",
X"5180da39",
X"f1a43f83",
X"c0800880",
X"ce38f1c4",
X"3f83c080",
X"08802eaa",
X"388151ef",
X"813febc7",
X"3f800b83",
X"c7d00cfb",
X"bb3f83c0",
X"800852ff",
X"0b83c7d0",
X"0cedcd3f",
X"71a13871",
X"51eedf3f",
X"9f39f0fb",
X"3f83c080",
X"08802e94",
X"388151ee",
X"cd3feb93",
X"3ff9913f",
X"edaa3f81",
X"51f28d3f",
X"833d0d04",
X"fe3d0d80",
X"5283c880",
X"5180cebd",
X"3f815283",
X"c7f05180",
X"ceb33f82",
X"80805380",
X"52818180",
X"8051f187",
X"3f80c080",
X"53805284",
X"81808051",
X"f1983f90",
X"80805286",
X"84808051",
X"ffb0fd3f",
X"83c08008",
X"a43881d2",
X"c051ffb5",
X"c03f83c7",
X"e8085381",
X"d1a05283",
X"c0800851",
X"ffb09f3f",
X"83c08008",
X"8438f3f1",
X"3f8151f1",
X"9b3ffe8d",
X"3ffc3983",
X"c08c0802",
X"83c08c0c",
X"fb3d0d02",
X"81d1ac0b",
X"83c39c0c",
X"81d0a40b",
X"83c3940c",
X"81d0a00b",
X"83c3a80c",
X"81d1b00b",
X"83c3a40c",
X"83c08c08",
X"fc050c80",
X"0b83c7d4",
X"0b83c08c",
X"08f8050c",
X"83c08c08",
X"f4050cff",
X"aef63f83",
X"c0800886",
X"05fc0683",
X"c08c08f0",
X"050c0283",
X"c08c08f0",
X"0508310d",
X"833d7083",
X"c08c08f8",
X"05087084",
X"0583c08c",
X"08f8050c",
X"0c51ffab",
X"be3f83c0",
X"8c08f405",
X"08810583",
X"c08c08f4",
X"050c83c0",
X"8c08f405",
X"08872e09",
X"8106ffab",
X"38869480",
X"8051e8d5",
X"3fff0b83",
X"c7d00c80",
X"0b83c894",
X"0c84d8c0",
X"0b83c890",
X"0c8151ec",
X"893f8151",
X"ecae3f80",
X"51eca93f",
X"8151eccf",
X"3f8251ec",
X"f73f8051",
X"ed9f3f80",
X"51edc93f",
X"80d0b952",
X"8051ddb9",
X"3ffda53f",
X"83c08c08",
X"fc05080d",
X"800b83c0",
X"800c873d",
X"0d83c08c",
X"0c04fc3d",
X"0d765580",
X"750c800b",
X"84160c80",
X"0b88160c",
X"83c88051",
X"80db823f",
X"83c7f051",
X"80dafa3f",
X"87d08933",
X"87d08f33",
X"70822a70",
X"81067030",
X"70720770",
X"09709f2c",
X"77069e06",
X"54515156",
X"51515454",
X"edcb3f80",
X"73980653",
X"5471882e",
X"09810683",
X"38815471",
X"98327030",
X"70802576",
X"71318419",
X"0c515152",
X"80738606",
X"53547182",
X"2e098106",
X"83388154",
X"71863270",
X"30708025",
X"76713178",
X"0c515152",
X"72943270",
X"30708025",
X"88180c51",
X"5283c080",
X"08802e80",
X"c23883c0",
X"8008812a",
X"70810683",
X"c0800881",
X"06318417",
X"0c5283c0",
X"8008832a",
X"83c08008",
X"822a7181",
X"06718106",
X"31770c53",
X"5383c080",
X"08842a81",
X"0688160c",
X"83c08008",
X"852a8106",
X"8c160c86",
X"3d0d04fe",
X"3d0d7476",
X"54527151",
X"fe903f72",
X"812ea238",
X"8173268d",
X"3872822e",
X"ab387283",
X"2e9f38e6",
X"397108e2",
X"38841208",
X"dd388812",
X"08d838a0",
X"39881208",
X"812e0981",
X"06cc3894",
X"39881208",
X"812e8d38",
X"71088938",
X"84120880",
X"2effb738",
X"843d0d04",
X"fb3d0d78",
X"0284059f",
X"05335556",
X"800b81cd",
X"d4565381",
X"732b7406",
X"5271802e",
X"83388152",
X"74708205",
X"56227073",
X"902b0790",
X"809c0c51",
X"81135372",
X"882e0981",
X"06d93880",
X"5383c89c",
X"13335170",
X"81ff2eb2",
X"38701081",
X"cbf40570",
X"22555180",
X"73177033",
X"701081cb",
X"f4057022",
X"51515152",
X"5273712e",
X"91388112",
X"5271862e",
X"098106f1",
X"38739080",
X"9c0c8113",
X"5372862e",
X"098106ff",
X"b8388053",
X"72167033",
X"51517081",
X"ff2e9438",
X"701081cb",
X"f4057022",
X"70848080",
X"0790809c",
X"0c515181",
X"13537286",
X"2e098106",
X"d7388053",
X"72165170",
X"3383c89c",
X"14348113",
X"5372862e",
X"098106ec",
X"38873d0d",
X"0404ff3d",
X"0d740284",
X"058f0533",
X"52527088",
X"38719080",
X"940c8e39",
X"70812e09",
X"81068638",
X"71908098",
X"0c833d0d",
X"04fb3d0d",
X"029f0533",
X"79982b70",
X"982c7c98",
X"2b70982c",
X"83c8b815",
X"70337098",
X"2b70982c",
X"51585c5a",
X"51555154",
X"5470732e",
X"09810694",
X"3883c898",
X"14337098",
X"2b70982c",
X"51525670",
X"722eb138",
X"72753471",
X"83c89815",
X"3483c899",
X"3383c8b9",
X"3371982b",
X"71902b07",
X"83c89833",
X"70882b72",
X"0783c8b8",
X"33710790",
X"80b80c52",
X"59535452",
X"873d0d04",
X"fe3d0d74",
X"81113371",
X"3371882b",
X"0783c080",
X"0c535184",
X"3d0d0483",
X"c8a43383",
X"c0800c04",
X"f53d0d02",
X"bb053302",
X"8405bf05",
X"33028805",
X"80c30533",
X"028c0580",
X"c6052266",
X"5c5a5e5c",
X"567a557b",
X"548953a1",
X"527d5180",
X"d0c03f83",
X"c0800881",
X"ff0683c0",
X"800c8d3d",
X"0d0483c0",
X"8c080283",
X"c08c0cf5",
X"3d0d83c0",
X"8c088805",
X"0883c08c",
X"088f0533",
X"83c08c08",
X"92052202",
X"8c057390",
X"0583c08c",
X"08e8050c",
X"83c08c08",
X"f8050c83",
X"c08c08f0",
X"050c83c0",
X"8c08ec05",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08f005",
X"0883c08c",
X"08e0050c",
X"83c08c08",
X"fc050c83",
X"c08c08f0",
X"05088927",
X"8a38890b",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"05088605",
X"87fffc06",
X"83c08c08",
X"e0050c02",
X"83c08c08",
X"e0050831",
X"0d853d70",
X"5583c08c",
X"08ec0508",
X"5483c08c",
X"08f00508",
X"5383c08c",
X"08f40508",
X"5283c08c",
X"08e4050c",
X"80d9f23f",
X"83c08008",
X"81ff0683",
X"c08c08e4",
X"050883c0",
X"8c08ec05",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"e0050880",
X"2e8c3883",
X"c08c08f8",
X"05080d89",
X"c83983c0",
X"8c08f005",
X"08802e89",
X"a63883c0",
X"8c08ec05",
X"08810533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508842e",
X"a938840b",
X"83c08c08",
X"e0050825",
X"88c73883",
X"c08c08e0",
X"0508852e",
X"859b3883",
X"c08c08e0",
X"0508a12e",
X"87ad3888",
X"ac39800b",
X"83c08c08",
X"ec050885",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08fc050c",
X"83c08c08",
X"e0050883",
X"2e098106",
X"88833883",
X"c08c08e8",
X"05088105",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e0050881",
X"2687e638",
X"810b83c0",
X"8c08e005",
X"0880d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08fc",
X"050c83c0",
X"8c08ec05",
X"08820533",
X"83c08c08",
X"e0050887",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088b",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"e005088c",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088d",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"e005088e",
X"052383c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"e005088a",
X"053483c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"70940508",
X"fcffff06",
X"7194050c",
X"83c08c08",
X"e0050c83",
X"c08c08ec",
X"05088605",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"f4050c83",
X"c08c08e0",
X"050883c0",
X"8c08fc05",
X"082e0981",
X"06b63883",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c83",
X"c08c08fc",
X"050883c0",
X"8c08e005",
X"088b0534",
X"83c08c08",
X"ec050887",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"812e8f38",
X"83c08c08",
X"e0050882",
X"2eb73884",
X"8c3983c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c820b",
X"83c08c08",
X"e005088a",
X"053483d9",
X"3983c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08fc0508",
X"83c08c08",
X"e005088a",
X"053483a1",
X"3983c08c",
X"08fc0508",
X"802e8395",
X"3883c08c",
X"08ec0508",
X"83053383",
X"0683c08c",
X"08e0050c",
X"83c08c08",
X"e0050883",
X"2e098106",
X"82f33883",
X"c08c08ec",
X"05088205",
X"3370982b",
X"83c08c08",
X"e0050c83",
X"c08c08e4",
X"050c83c0",
X"8c08e005",
X"08802582",
X"cc3883c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c83",
X"c08c08f4",
X"050c83c0",
X"8c08ec05",
X"08860533",
X"83c08c08",
X"e0050880",
X"d6053483",
X"c08c08e0",
X"05088405",
X"83c08c08",
X"ec050882",
X"05338f06",
X"83c08c08",
X"e4050c83",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0883c08c",
X"08e00508",
X"3483c08c",
X"08ec0508",
X"84053383",
X"c08c08e0",
X"05088105",
X"34800b83",
X"c08c08e0",
X"05088205",
X"3483c08c",
X"08e00508",
X"08ff83ff",
X"06828007",
X"83c08c08",
X"e005080c",
X"83c08c08",
X"e8050881",
X"05338105",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"050883c0",
X"8c08e805",
X"08810534",
X"81833983",
X"c08c08fc",
X"0508802e",
X"80f73883",
X"c08c08ec",
X"05088605",
X"3383c08c",
X"08e0050c",
X"83c08c08",
X"e00508a2",
X"2e098106",
X"80d73883",
X"c08c08ec",
X"05088805",
X"3383c08c",
X"08ec0508",
X"87053371",
X"82802905",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c5283c0",
X"8c08e405",
X"0c83c08c",
X"08f4050c",
X"83c08c08",
X"e4050883",
X"c08c08e0",
X"05088805",
X"2383c08c",
X"08ec0508",
X"3383c08c",
X"08f00508",
X"71317083",
X"ffff0683",
X"c08c08f0",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08ec0508",
X"0583c08c",
X"08ec050c",
X"f6d03983",
X"c08c08f8",
X"05080d83",
X"c08c08f0",
X"050883c0",
X"8c08e005",
X"0c83c08c",
X"08f80508",
X"0d83c08c",
X"08e00508",
X"83c0800c",
X"8d3d0d83",
X"c08c0c04",
X"83c08c08",
X"0283c08c",
X"0ce63d0d",
X"83c08c08",
X"88050802",
X"840583c0",
X"8c08e805",
X"0c83c08c",
X"08d4050c",
X"800b83c8",
X"c03483c0",
X"8c08d405",
X"08900583",
X"c08c08c0",
X"050c800b",
X"83c08c08",
X"c0050834",
X"800b83c0",
X"8c08c005",
X"08810534",
X"800b83c0",
X"8c08c405",
X"0c83c08c",
X"08c40508",
X"80d82983",
X"c08c08c0",
X"05080583",
X"c08c08ff",
X"b4050c80",
X"0b83c08c",
X"08ffb405",
X"0880d805",
X"0c83c08c",
X"08ffb405",
X"08840583",
X"c08c08ff",
X"b4050c83",
X"c08c08c4",
X"050883c0",
X"8c08ffb4",
X"05083488",
X"0b83c08c",
X"08ffb405",
X"08810534",
X"800b83c0",
X"8c08ffb4",
X"05088205",
X"3483c08c",
X"08ffb405",
X"0808ffa1",
X"ff06a080",
X"0783c08c",
X"08ffb405",
X"080c83c0",
X"8c08c405",
X"08810570",
X"81ff0683",
X"c08c08c4",
X"050c83c0",
X"8c08ffb4",
X"050c810b",
X"83c08c08",
X"c4050827",
X"fedb3883",
X"c08c08ec",
X"05705483",
X"c08c08c8",
X"050c9252",
X"83c08c08",
X"d4050851",
X"80cd993f",
X"83c08008",
X"81ff0670",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"8dea3883",
X"c08c08f4",
X"0551f18c",
X"3f83c080",
X"0883ffff",
X"0683c08c",
X"08f60552",
X"83c08c08",
X"e4050cf0",
X"f33f83c0",
X"800883ff",
X"ff0683c0",
X"8c08fd05",
X"3383c08c",
X"08ffb805",
X"0883c08c",
X"08c4050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"e0050c83",
X"c08c08c4",
X"050883c0",
X"8c08ffbc",
X"05082780",
X"fe3883c0",
X"8c08c805",
X"085483c0",
X"8c08c405",
X"08538952",
X"83c08c08",
X"d4050851",
X"80cc9e3f",
X"83c08008",
X"81ff0683",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b8050880",
X"f23883c0",
X"8c08ee05",
X"51eff13f",
X"83c08008",
X"83ffff06",
X"5383c08c",
X"08c40508",
X"5283c08c",
X"08d40508",
X"51f0b33f",
X"83c08c08",
X"c4050881",
X"057081ff",
X"0683c08c",
X"08c4050c",
X"83c08c08",
X"ffb4050c",
X"fef13983",
X"c08c08c0",
X"05088105",
X"3383c08c",
X"08ffb405",
X"0c81db0b",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb40508",
X"802e8be0",
X"38943983",
X"c08c08ff",
X"b8050883",
X"c08c08ff",
X"bc050c8b",
X"cb3983c0",
X"8c08f105",
X"335283c0",
X"8c08d405",
X"085180cb",
X"9c3f800b",
X"83c08c08",
X"c0050881",
X"053383c0",
X"8c08ffb4",
X"050c83c0",
X"8c08c405",
X"0c83c08c",
X"08c40508",
X"83c08c08",
X"ffb40508",
X"2789e638",
X"83c08c08",
X"c4050880",
X"d8297083",
X"c08c08c0",
X"05080570",
X"88057083",
X"053383c0",
X"8c08cc05",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"d8050c83",
X"c08c08cc",
X"050887a6",
X"3883c08c",
X"08c80508",
X"22028405",
X"71860587",
X"fffc0683",
X"c08c08ff",
X"b4050c83",
X"c08c08dc",
X"050c83c0",
X"8c08ffb8",
X"050c0283",
X"c08c08ff",
X"b4050831",
X"0d893d70",
X"5983c08c",
X"08ffb805",
X"085883c0",
X"8c08ffbc",
X"05088705",
X"335783c0",
X"8c08ffb4",
X"050ca255",
X"83c08c08",
X"cc050854",
X"86538181",
X"5283c08c",
X"08d40508",
X"51be933f",
X"83c08008",
X"81ff0683",
X"c08c08d0",
X"050c83c0",
X"8c08d005",
X"0881c138",
X"83c08c08",
X"ffbc0508",
X"96055383",
X"c08c08ff",
X"b8050852",
X"83c08c08",
X"ffb40508",
X"51a1c63f",
X"83c08008",
X"81ff0683",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b4050880",
X"2e818538",
X"83c08c08",
X"ffbc0508",
X"940583c0",
X"8c08ffbc",
X"05089605",
X"3370862a",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"cc050c83",
X"c08c08ff",
X"b4050883",
X"2e098106",
X"80c63883",
X"c08c08ff",
X"b4050883",
X"c08c08c8",
X"05088205",
X"3483c8a4",
X"33708105",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb40508",
X"83c8a434",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"cc050834",
X"83c08c08",
X"dc05080d",
X"83c08c08",
X"d0050881",
X"ff0683c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"0508fbff",
X"3883c08c",
X"08d80508",
X"83c08c08",
X"c0050805",
X"88057082",
X"05335183",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b4050883",
X"2e098106",
X"80e33883",
X"c08c08ff",
X"b8050883",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b4050881",
X"057081ff",
X"065183c0",
X"8c08ffb4",
X"050c810b",
X"83c08c08",
X"ffb40508",
X"27dd3880",
X"0b83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb405",
X"08810570",
X"81ff0651",
X"83c08c08",
X"ffb4050c",
X"970b83c0",
X"8c08ffb4",
X"050827dd",
X"3883c08c",
X"08e40508",
X"80f93270",
X"30708025",
X"515183c0",
X"8c08ffb4",
X"050c83c0",
X"8c08e005",
X"08912e09",
X"810680f9",
X"3883c08c",
X"08ffb405",
X"08802e80",
X"ec3883c0",
X"8c08c405",
X"0880e238",
X"850b83c0",
X"8c08c005",
X"08a60534",
X"a00b83c0",
X"8c08c005",
X"08a70534",
X"850b83c0",
X"8c08c005",
X"08a80534",
X"80c00b83",
X"c08c08c0",
X"0508a905",
X"34860b83",
X"c08c08c0",
X"0508aa05",
X"34900b83",
X"c08c08c0",
X"0508ab05",
X"34860b83",
X"c08c08c0",
X"0508ac05",
X"34a00b83",
X"c08c08c0",
X"0508ad05",
X"3483c08c",
X"08e40508",
X"89d83270",
X"30708025",
X"515183c0",
X"8c08ffb4",
X"050c83c0",
X"8c08e005",
X"0883edec",
X"2e098106",
X"80f63881",
X"7083c08c",
X"08ffb405",
X"080683c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb4",
X"0508802e",
X"80ce3883",
X"c08c08c4",
X"050880c4",
X"38840b83",
X"c08c08c0",
X"0508aa05",
X"3480c00b",
X"83c08c08",
X"c00508ab",
X"0534840b",
X"83c08c08",
X"c00508ac",
X"0534900b",
X"83c08c08",
X"c00508ad",
X"053483c0",
X"8c08ffb8",
X"050883c0",
X"8c08c005",
X"088c0534",
X"83c08c08",
X"e4050880",
X"f9327030",
X"70802551",
X"5183c08c",
X"08ffb405",
X"0c83c08c",
X"08e00508",
X"862e0981",
X"0680c338",
X"817083c0",
X"8c08ffb4",
X"05080683",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b4050880",
X"2e9c3883",
X"c08c08c4",
X"05089338",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"c005088d",
X"053483c0",
X"8c08c405",
X"0880d829",
X"83c08c08",
X"c0050805",
X"70840570",
X"83053383",
X"c08c08ff",
X"b4050c83",
X"c08c08c8",
X"050c83c0",
X"8c08ffbc",
X"050c8058",
X"805783c0",
X"8c08ffb4",
X"05085680",
X"5580548a",
X"53a15283",
X"c08c08d4",
X"050851b7",
X"8d3f83c0",
X"800881ff",
X"06703070",
X"9f2a5183",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"b80508a0",
X"2e8c3883",
X"c08c08ff",
X"b40508f6",
X"c23883c0",
X"8c08ffbc",
X"05088b05",
X"3383c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb405",
X"08802eb3",
X"3883c08c",
X"08c80508",
X"83053383",
X"c08c08ff",
X"b4050c80",
X"58805783",
X"c08c08ff",
X"b4050856",
X"80558054",
X"8b53a152",
X"83c08c08",
X"d4050851",
X"b6883f83",
X"c08c08c4",
X"05088105",
X"7081ff06",
X"83c08c08",
X"c0050881",
X"05335283",
X"c08c08c4",
X"050c83c0",
X"8c08ffb4",
X"050cf689",
X"39800b83",
X"c08c08c4",
X"050c83c0",
X"8c08c405",
X"0880d829",
X"83c08c08",
X"d4050805",
X"709a0533",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb40508",
X"822e0981",
X"06a93883",
X"c8c05681",
X"55805483",
X"c08c08ff",
X"b4050853",
X"83c08c08",
X"ffb80508",
X"97053352",
X"83c08c08",
X"d4050851",
X"e48a3f83",
X"c08c08c4",
X"05088105",
X"7081ff06",
X"83c08c08",
X"c4050c83",
X"c08c08ff",
X"b4050c81",
X"0b83c08c",
X"08c40508",
X"27fefb38",
X"810b83c0",
X"8c08c005",
X"0834800b",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"e805080d",
X"83c08c08",
X"ffbc0508",
X"83c0800c",
X"9c3d0d83",
X"c08c0c04",
X"f53d0d90",
X"1e57800b",
X"81183354",
X"59787327",
X"819d3878",
X"80d82917",
X"8a113354",
X"5472832e",
X"09810680",
X"f8389414",
X"335ba98c",
X"3f83c080",
X"085a8056",
X"7581c429",
X"1a871133",
X"54547280",
X"2e80c038",
X"730881cb",
X"e82e0981",
X"06b53880",
X"74595574",
X"80d82918",
X"9a113354",
X"5472832e",
X"09810692",
X"38a41470",
X"3354547a",
X"73278738",
X"ff135372",
X"74348115",
X"7081ff06",
X"56538175",
X"27d13881",
X"167081ff",
X"0657538f",
X"7627ffa4",
X"3883c8a4",
X"33ff0553",
X"7283c8a4",
X"34811970",
X"81ff0681",
X"19335e5a",
X"537b7926",
X"fee53880",
X"0b83c080",
X"0c8d3d0d",
X"0483c08c",
X"080283c0",
X"8c0ce63d",
X"0d83c08c",
X"08880508",
X"02840571",
X"90057033",
X"7083c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"dc050c83",
X"c08c08e0",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"94b53880",
X"0b83c08c",
X"08c80508",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08d4",
X"050c83c0",
X"8c08d405",
X"0883c08c",
X"08ffa405",
X"082593fd",
X"3883c08c",
X"08d40508",
X"80d82983",
X"c08c08c8",
X"05080584",
X"05708605",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffa405",
X"08802e93",
X"8938a6b2",
X"3f83c08c",
X"08ffb805",
X"0880d405",
X"0883c080",
X"082692f2",
X"380283c0",
X"8c08ffb8",
X"05088105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08d8050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"fc052383",
X"c08c08ff",
X"a4050886",
X"0583fc06",
X"83c08c08",
X"ffa4050c",
X"0283c08c",
X"08ffa405",
X"08310d85",
X"3d705583",
X"c08c08fc",
X"055483c0",
X"8c08ffb8",
X"05085383",
X"c08c08e0",
X"05085283",
X"c08c08c0",
X"050cae8a",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"91bb3883",
X"c08c08ff",
X"b8050887",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"80d53883",
X"c08c08ff",
X"b8050886",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508822e",
X"098106b3",
X"3883c08c",
X"08fc0522",
X"83c08c08",
X"ffa4050c",
X"870b83c0",
X"8c08ffa4",
X"05082797",
X"3883c08c",
X"08c00508",
X"82055283",
X"c08c08c0",
X"05083351",
X"dba63f83",
X"c08c08ff",
X"b8050886",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508832e",
X"09810690",
X"a43883c0",
X"8c08ffb8",
X"05089205",
X"70820533",
X"83c08c08",
X"fc052283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08c4",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffa8",
X"0508268f",
X"e438800b",
X"83c08c08",
X"e4050c80",
X"0b83c08c",
X"08ffb005",
X"0c83c08c",
X"08ffb005",
X"081083c0",
X"8c0805f8",
X"0583c08c",
X"08ffb005",
X"08842983",
X"c08c08ff",
X"b0050810",
X"0583c08c",
X"08c40508",
X"05708405",
X"703383c0",
X"8c08c005",
X"08057033",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffbc0508",
X"2383c08c",
X"08ffa805",
X"08810533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"902e0981",
X"06be3883",
X"c08c08ff",
X"a8050833",
X"83c08c08",
X"c0050805",
X"81057033",
X"70828029",
X"83c08c08",
X"ffb40508",
X"05515183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"bc050823",
X"83c08c08",
X"ffac0508",
X"86052283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a80508a2",
X"3883c08c",
X"08ffac05",
X"08880522",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"81ff2e80",
X"e53883c0",
X"8c08ffbc",
X"05082270",
X"83c08c08",
X"ffa80508",
X"31708280",
X"29713183",
X"c08c08ff",
X"ac050888",
X"05227083",
X"c08c08ff",
X"a8050831",
X"70733553",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffac050c",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffbc05",
X"082383c0",
X"8c08ffb0",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa4050c",
X"810b83c0",
X"8c08ffb0",
X"050827fc",
X"e03883c0",
X"8c08f805",
X"2283c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08bf2691",
X"3883c08c",
X"08e40508",
X"820783c0",
X"8c08e405",
X"0c81c00b",
X"83c08c08",
X"ffa40508",
X"27913883",
X"c08c08e4",
X"05088107",
X"83c08c08",
X"e4050c83",
X"c08c08fa",
X"052283c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508bf26",
X"913883c0",
X"8c08e405",
X"08880783",
X"c08c08e4",
X"050c81c0",
X"0b83c08c",
X"08ffa405",
X"08279138",
X"83c08c08",
X"e4050884",
X"0783c08c",
X"08e4050c",
X"800b83c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffb0",
X"05081083",
X"c08c08c4",
X"05080570",
X"90057033",
X"83c08c08",
X"c0050805",
X"70337281",
X"05337072",
X"06515351",
X"83c08c08",
X"ffa8050c",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e9b",
X"38900b83",
X"c08c08ff",
X"b005082b",
X"83c08c08",
X"e4050807",
X"83c08c08",
X"e4050c83",
X"c08c08ff",
X"b0050881",
X"057081ff",
X"0683c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa405",
X"0c970b83",
X"c08c08ff",
X"b0050827",
X"fef43883",
X"c08c08ff",
X"b8050890",
X"053383c0",
X"8c08e405",
X"0883c08c",
X"08ffb405",
X"0c83c08c",
X"08c4050c",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffb80508",
X"8c05082e",
X"83ff3883",
X"c08c08ff",
X"b4050883",
X"c08c08ff",
X"b805088c",
X"050c83c0",
X"8c08ffb8",
X"05088905",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e83",
X"b93883c0",
X"8c08e405",
X"83c08c08",
X"ffb40508",
X"8f0683c0",
X"8c08e405",
X"0c83c08c",
X"08cc050c",
X"800b83c0",
X"8c08f005",
X"0c800b83",
X"c08c08f4",
X"0523800b",
X"81cde433",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffbc0508",
X"2e82d338",
X"83c08c08",
X"f00581cd",
X"e40b83c0",
X"8c08ffac",
X"050c83c0",
X"8c08d005",
X"0c83c08c",
X"08ffac05",
X"083383c0",
X"8c08ffac",
X"05088105",
X"3381722b",
X"81722b07",
X"7083c08c",
X"08ffb405",
X"08065283",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"a805082e",
X"09810681",
X"be3883c0",
X"8c08ffbc",
X"05088526",
X"80f63883",
X"c08c08ff",
X"ac050882",
X"05337081",
X"ff0683c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"80ca3883",
X"c08c08ff",
X"bc050883",
X"c08c08ff",
X"bc050881",
X"057081ff",
X"0683c08c",
X"08d00508",
X"73055383",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b0050883",
X"c08c08ff",
X"a4050834",
X"83c08c08",
X"ffac0508",
X"83053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e9d3881",
X"0b83c08c",
X"08ffa405",
X"082b83c0",
X"8c08cc05",
X"08080783",
X"c08c08cc",
X"05080c83",
X"c08c08ff",
X"ac050884",
X"05703383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a40508fd",
X"c83883c0",
X"8c08f005",
X"528051d0",
X"c33f83c0",
X"8c08e405",
X"085283c0",
X"8c08c405",
X"0851d1fe",
X"3f83c08c",
X"08fb0533",
X"7081800a",
X"29810a05",
X"70982c55",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"f9053370",
X"81800a29",
X"810a0570",
X"982c5583",
X"c08c08ff",
X"a4050c83",
X"c08c08c4",
X"05085383",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a8050cd1",
X"d43f83c0",
X"8c08ffb8",
X"05088805",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e84",
X"e03883c0",
X"8c08ffb8",
X"05089005",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08812684",
X"c0388070",
X"81ce980b",
X"81ce980b",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"b405082e",
X"81ae3883",
X"c08c08ff",
X"ac050884",
X"2983c08c",
X"08ffa805",
X"08057033",
X"83c08c08",
X"c0050805",
X"70337281",
X"05337072",
X"06515351",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802eaa38",
X"810b83c0",
X"8c08ffac",
X"05082b83",
X"c08c08ff",
X"b4050807",
X"7083ffff",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffac05",
X"08810570",
X"81ff0681",
X"ce987184",
X"29710570",
X"81053351",
X"5383c08c",
X"08ffa805",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08fed438",
X"83c08c08",
X"ffb80508",
X"8a052283",
X"c08c08c0",
X"050c83c0",
X"8c08ffb4",
X"050883c0",
X"8c08c005",
X"082e82ad",
X"38800b83",
X"c08c08e8",
X"050c800b",
X"83c08c08",
X"ec052380",
X"7083c08c",
X"08e80583",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"b0050c81",
X"af3983c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffac",
X"05082c70",
X"81065183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e80e738",
X"83c08c08",
X"ffb00508",
X"83c08c08",
X"ffb00508",
X"81057081",
X"ff0683c0",
X"8c08ffbc",
X"05087305",
X"83c08c08",
X"ffb80508",
X"90053383",
X"c08c08ff",
X"ac050884",
X"29055353",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa8050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa80508",
X"81ce9a05",
X"3383c08c",
X"08ffa405",
X"083483c0",
X"8c08ffac",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"ffa4050c",
X"8f0b83c0",
X"8c08ffac",
X"05082783",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b0050885",
X"268c3883",
X"c08c08ff",
X"a40508fe",
X"a93883c0",
X"8c08e805",
X"528051ca",
X"f33f83c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffb8",
X"05088a05",
X"2383c08c",
X"08ffb805",
X"0880d205",
X"3383c08c",
X"08ffb805",
X"0880d405",
X"080583c0",
X"8c08ffb8",
X"050880d4",
X"050c83c0",
X"8c08d805",
X"080d83c0",
X"8c08d405",
X"0881800a",
X"2981800a",
X"0570982c",
X"83c08c08",
X"c8050881",
X"053383c0",
X"8c08ffa8",
X"050c5183",
X"c08c08d4",
X"050c83c0",
X"8c08ffa8",
X"050883c0",
X"8c08d405",
X"0824ec85",
X"38800b83",
X"c08c08ff",
X"a8050c83",
X"c08c08dc",
X"05080d83",
X"c08c08ff",
X"a8050883",
X"c0800c9c",
X"3d0d83c0",
X"8c0c04f3",
X"3d0d02bf",
X"05330284",
X"0580c305",
X"3383c8c0",
X"335a5b59",
X"79802e8d",
X"38787806",
X"5776802e",
X"8e388189",
X"39787806",
X"5776802e",
X"80ff3883",
X"c8c03370",
X"7a075858",
X"79883878",
X"09707906",
X"51577683",
X"c8c03492",
X"973f83c0",
X"80085e80",
X"5c8f5d7d",
X"1c871133",
X"58587680",
X"2e80c138",
X"770881cb",
X"e82e0981",
X"06b63880",
X"5b815a7d",
X"1c701c9a",
X"11335959",
X"5976822e",
X"09810694",
X"3883c8c0",
X"56815580",
X"54765397",
X"18335278",
X"51cbc53f",
X"ff1a80d8",
X"1c5c5a79",
X"8025d038",
X"ff1d81c4",
X"1d5d5d7c",
X"8025ffa7",
X"388f3d0d",
X"04e93d0d",
X"696c0288",
X"0580ea05",
X"225c5a5b",
X"80707141",
X"5e58ff78",
X"797a7b7c",
X"7d464c4a",
X"45405d43",
X"62993d34",
X"62028405",
X"80dd0534",
X"77792280",
X"ffff0654",
X"45727923",
X"79782e88",
X"87387a70",
X"81055c33",
X"70842a71",
X"8c067082",
X"2a5a5656",
X"8306ff1b",
X"7083ffff",
X"065c5456",
X"80547574",
X"2e91387a",
X"7081055c",
X"33ff1b70",
X"83ffff06",
X"5c545481",
X"76279b38",
X"7381ff06",
X"7b708105",
X"5d335574",
X"82802905",
X"ff1b7083",
X"ffff065c",
X"54548276",
X"27aa3873",
X"83ffff06",
X"7b708105",
X"5d337090",
X"2b72077d",
X"7081055f",
X"3370982b",
X"7207fe1f",
X"7083ffff",
X"06405252",
X"52525454",
X"7e802e80",
X"c4387686",
X"f738748a",
X"2e098106",
X"9438811f",
X"7081ff06",
X"811e7081",
X"ff065f52",
X"405386dc",
X"39748c2e",
X"09810686",
X"d338ff1f",
X"7081ff06",
X"ff1e7081",
X"ff065f52",
X"40537b63",
X"2586bd38",
X"ff4386b8",
X"3976812e",
X"83bb3876",
X"81248938",
X"76802e8d",
X"3886a539",
X"76822e84",
X"a638869c",
X"39f81553",
X"72842684",
X"95387284",
X"2981ced8",
X"05537208",
X"0464802e",
X"80cd3878",
X"22838080",
X"06537283",
X"80802e09",
X"8106bc38",
X"80567564",
X"27a43875",
X"1e7083ff",
X"ff067710",
X"1b901172",
X"832a5851",
X"57515373",
X"75347287",
X"0681712b",
X"51537281",
X"16348116",
X"7081ff06",
X"57539776",
X"27cc387f",
X"84074080",
X"0b993d43",
X"56611670",
X"3370982b",
X"70982c51",
X"51515380",
X"732480fb",
X"38607329",
X"1e7083ff",
X"ff067a22",
X"83808006",
X"52585372",
X"8380802e",
X"09810680",
X"de386088",
X"32703070",
X"72078025",
X"63903270",
X"30707207",
X"80257307",
X"53545851",
X"55537380",
X"2ebd3876",
X"87065372",
X"b6387584",
X"29761005",
X"79118411",
X"79832a57",
X"57515373",
X"75346081",
X"16346586",
X"14236688",
X"14237587",
X"387f8107",
X"408d3975",
X"812e0981",
X"0685387f",
X"82074081",
X"167081ff",
X"06575381",
X"7627fee5",
X"38636129",
X"1e7083ff",
X"ff065f53",
X"80704642",
X"ff028405",
X"80dd0534",
X"ff0b993d",
X"3483f539",
X"811c7081",
X"ff065d53",
X"80427381",
X"2e098106",
X"8e387781",
X"800a2981",
X"800a0558",
X"80d33973",
X"802e8938",
X"73822e09",
X"81068d38",
X"7c81800a",
X"2981800a",
X"055da439",
X"815f83b8",
X"39ff1c70",
X"81ff065d",
X"537b6325",
X"8338ff43",
X"7c802e92",
X"387c8180",
X"0a2981ff",
X"0a055d7c",
X"982c5d83",
X"93397780",
X"2e923877",
X"81800a29",
X"81ff0a05",
X"5877982c",
X"5882fd39",
X"7753839e",
X"39748926",
X"80f43874",
X"842981ce",
X"ec055372",
X"08047387",
X"2e82e138",
X"73852e82",
X"db387388",
X"2e82d538",
X"738c2e82",
X"cf387389",
X"2e098106",
X"86388145",
X"82c23973",
X"812e0981",
X"0682b938",
X"62802582",
X"b3387b98",
X"2b70982c",
X"514382a8",
X"397383ff",
X"ff064682",
X"9f397383",
X"ffff0647",
X"82963973",
X"81ff0641",
X"828e3973",
X"811a3482",
X"87397381",
X"ff064481",
X"ff397e53",
X"82a03974",
X"812e81e3",
X"38748124",
X"89387480",
X"2e8d3881",
X"e7397482",
X"2e81d838",
X"81de3974",
X"567b8338",
X"81567453",
X"73862e09",
X"81069738",
X"75810653",
X"72802e8e",
X"38782282",
X"ffff06fe",
X"80800753",
X"b6397b83",
X"38815373",
X"822e0981",
X"06973872",
X"81065372",
X"802e8e38",
X"782281ff",
X"ff068180",
X"80075393",
X"397b9638",
X"fc145372",
X"81268e38",
X"7822ff80",
X"80075372",
X"792380e5",
X"39805573",
X"812e0981",
X"06833873",
X"55775377",
X"802e8938",
X"74810653",
X"7280ca38",
X"72d01554",
X"55728126",
X"83388155",
X"77802eb9",
X"38748106",
X"5372802e",
X"b0387822",
X"83808006",
X"53728380",
X"802e0981",
X"069f3873",
X"b02e0981",
X"06873861",
X"993d3491",
X"3973b12e",
X"09810689",
X"38610284",
X"0580dd05",
X"34618105",
X"538c3961",
X"74318105",
X"53843961",
X"14537283",
X"ffff0642",
X"79f7fb38",
X"7d832a53",
X"72821a34",
X"78228380",
X"80065372",
X"8380802e",
X"09810688",
X"3881537f",
X"872e8338",
X"80537283",
X"c0800c99",
X"3d0d04fd",
X"3d0d7583",
X"11338212",
X"3371982b",
X"71902b07",
X"81143370",
X"882b7207",
X"75337107",
X"83c0800c",
X"52535456",
X"5452853d",
X"0d04f63d",
X"0d02b705",
X"33028405",
X"bb053302",
X"8805bf05",
X"335b5b5b",
X"80588057",
X"78882b7a",
X"07568055",
X"7a548153",
X"a3527c51",
X"92cc3f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f63d",
X"0d02b705",
X"33028405",
X"bb053302",
X"8805bf05",
X"335b5b5b",
X"80588057",
X"78882b7a",
X"07568055",
X"7a548353",
X"a3527c51",
X"92903f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f73d",
X"0d02b305",
X"33028405",
X"b6052260",
X"5a585680",
X"55805480",
X"5381a352",
X"7b5191e2",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8b3d0d04",
X"ee3d0d64",
X"90115c5c",
X"807b3480",
X"0b841c0c",
X"800b881c",
X"34810b89",
X"1c34880b",
X"8a1c3480",
X"0b8b1c34",
X"881b08c1",
X"06810788",
X"1c0c8f3d",
X"70545d88",
X"527b519b",
X"eb3f83c0",
X"800881ff",
X"06705b59",
X"7881a938",
X"903d335e",
X"81db5a7d",
X"892e0981",
X"06819938",
X"7c539252",
X"7b519bc4",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"8182387c",
X"58885778",
X"56a95578",
X"54865381",
X"a0527b51",
X"90d03f83",
X"c0800881",
X"ff06705b",
X"597880e0",
X"3802ba05",
X"337b347c",
X"5478537d",
X"527b519b",
X"ac3f83c0",
X"800881ff",
X"06705b59",
X"7880c138",
X"02bd0533",
X"527b519b",
X"c43f83c0",
X"800881ff",
X"06705b59",
X"78aa3881",
X"7b335a5a",
X"79792699",
X"38805479",
X"5388527b",
X"51fdbb3f",
X"811a7081",
X"ff067c33",
X"525b59e4",
X"39810b88",
X"1c34805a",
X"7983c080",
X"0c943d0d",
X"04800b83",
X"c0800c04",
X"f93d0d79",
X"028405ab",
X"05338e3d",
X"70545858",
X"58ffbeb0",
X"3f8a3d8a",
X"0551ffbe",
X"a73f7551",
X"fc8d3f83",
X"c0800884",
X"86812ebe",
X"3883c080",
X"08848681",
X"26993883",
X"c0800884",
X"82802e80",
X"e63883c0",
X"80088482",
X"812e9f38",
X"81b43983",
X"c0800880",
X"c082832e",
X"80f43883",
X"c0800880",
X"c086832e",
X"80e83881",
X"993983c0",
X"9c335580",
X"5674762e",
X"09810681",
X"8b387454",
X"76539152",
X"7751fbd6",
X"3f745476",
X"53905277",
X"51fbcb3f",
X"74547653",
X"84527751",
X"fbfc3f81",
X"0b83c09c",
X"3481b156",
X"80de3980",
X"54765391",
X"527751fb",
X"a93f8054",
X"76539052",
X"7751fb9e",
X"3f800b83",
X"c09c3476",
X"52871833",
X"5197963f",
X"b5398054",
X"76539452",
X"7751fb82",
X"3f805476",
X"53905277",
X"51faf73f",
X"7551ffbc",
X"db3f83c0",
X"8008892a",
X"81065376",
X"52871833",
X"5190cd3f",
X"800b83c0",
X"9c348056",
X"7583c080",
X"0c893d0d",
X"04f23d0d",
X"6090115a",
X"58800b88",
X"1a337159",
X"56567476",
X"2e82a538",
X"82ac3f84",
X"190883c0",
X"80082682",
X"95387833",
X"5a810b8e",
X"3d23903d",
X"f81155f4",
X"05539918",
X"5277518a",
X"e53f83c0",
X"800881ff",
X"06705755",
X"74772e09",
X"810681d9",
X"38863974",
X"5681d239",
X"81568257",
X"8e3d3377",
X"06557480",
X"2ebb3880",
X"0b8d3d34",
X"903df005",
X"54845375",
X"527751fa",
X"cd3f83c0",
X"800881ff",
X"0655749d",
X"387b5375",
X"527751fc",
X"e73f83c0",
X"800881ff",
X"06557481",
X"b12e818b",
X"3874ffb3",
X"38761081",
X"fc068117",
X"7081ff06",
X"58565787",
X"7627ffa8",
X"38815675",
X"7a2680eb",
X"38800b8d",
X"3d348c3d",
X"70555784",
X"53755277",
X"51f9f73f",
X"83c08008",
X"81ff0655",
X"7480c138",
X"7651ffba",
X"d73f83c0",
X"80088287",
X"06557482",
X"812e0981",
X"06aa3802",
X"ae053381",
X"07557402",
X"8405ae05",
X"347b5375",
X"527751fb",
X"eb3f83c0",
X"800881ff",
X"06557481",
X"b12e9038",
X"74feb838",
X"81167081",
X"ff065755",
X"ff913980",
X"567581ff",
X"0656973f",
X"83c08008",
X"8fd00584",
X"1a0c7557",
X"7683c080",
X"0c903d0d",
X"04049080",
X"a00883c0",
X"800c04ff",
X"3d0d7387",
X"e82951ff",
X"a2e03f83",
X"3d0d0404",
X"83c8c40b",
X"83c0800c",
X"04fd3d0d",
X"75775454",
X"800b83c8",
X"a434728a",
X"38909080",
X"0b84150c",
X"90397281",
X"2e098106",
X"88389098",
X"800b8415",
X"0c841408",
X"83c8bc0c",
X"800b8815",
X"0c800b8c",
X"150c83c8",
X"bc085382",
X"0b878014",
X"348151ff",
X"9e3f83c8",
X"bc085380",
X"0b881434",
X"83c8bc08",
X"53810b87",
X"80143483",
X"c8bc0853",
X"800b8c14",
X"3483c8bc",
X"0853800b",
X"a4143491",
X"7434800b",
X"83c0a034",
X"800b83c0",
X"a434800b",
X"83c0a834",
X"80547381",
X"c42983c8",
X"c8055380",
X"0b831434",
X"81147081",
X"ff065553",
X"8f7427e6",
X"38853d0d",
X"04fe3d0d",
X"74768211",
X"3370bf06",
X"81712bff",
X"05565151",
X"52539071",
X"278338ff",
X"52765171",
X"712383c8",
X"bc085187",
X"13339012",
X"34800b83",
X"c0a43480",
X"0b83c0a8",
X"34881333",
X"8a143352",
X"5271802e",
X"aa387081",
X"ff065184",
X"52708338",
X"70527183",
X"c0a4348a",
X"13337030",
X"70802584",
X"2b708807",
X"51515253",
X"7083c0a8",
X"34903970",
X"81ff0651",
X"70833898",
X"527183c0",
X"a834800b",
X"83c0800c",
X"843d0d04",
X"f13d0d61",
X"6568028c",
X"0580cb05",
X"33029005",
X"80ce0522",
X"02940580",
X"d6052242",
X"40415a40",
X"40fd8b3f",
X"83c08008",
X"a788055b",
X"8070715b",
X"5b528394",
X"3983c8bc",
X"08517d94",
X"123483c0",
X"a4338107",
X"55807054",
X"567f8626",
X"80ea387f",
X"842981cf",
X"a00583c8",
X"bc085351",
X"70080480",
X"0b841334",
X"a1397733",
X"70307080",
X"25837131",
X"51515253",
X"70841334",
X"8d39810b",
X"841334b8",
X"39830b84",
X"13348170",
X"5456ad39",
X"810b8413",
X"34a23977",
X"33703070",
X"80258371",
X"31515152",
X"53708413",
X"34807833",
X"52527083",
X"38815271",
X"78348153",
X"74880755",
X"83c0a833",
X"83c8bc08",
X"5257810b",
X"81d01234",
X"83c8bc08",
X"51810b81",
X"9012347e",
X"802eae38",
X"72802ea9",
X"387eff1e",
X"52547083",
X"ffff0653",
X"7283ffff",
X"2e973873",
X"70810555",
X"3383c8bc",
X"08535170",
X"81c01334",
X"ff1351de",
X"3983c8bc",
X"08a81133",
X"53517688",
X"123483c8",
X"bc085174",
X"713481ff",
X"52913983",
X"c8bc08a0",
X"11337081",
X"06515253",
X"708f38fa",
X"fd3f7a83",
X"c0800826",
X"e6388188",
X"39810ba0",
X"143483c8",
X"bc08a811",
X"3380ff06",
X"70780752",
X"53517080",
X"2e80ed38",
X"71862a70",
X"81065151",
X"70802e91",
X"38807833",
X"52537083",
X"38815372",
X"783480e0",
X"3971842a",
X"70810651",
X"5170802e",
X"9b388119",
X"7083ffff",
X"067d3070",
X"9f2a5152",
X"5a51787c",
X"2e098106",
X"af38a439",
X"71832a70",
X"81065151",
X"70802e93",
X"38811a70",
X"81ff065b",
X"5179832e",
X"09810690",
X"388a3971",
X"a3065170",
X"802e8538",
X"71519239",
X"f9e43f7a",
X"83c08008",
X"26fce238",
X"7181bf06",
X"517083c0",
X"800c913d",
X"0d04f63d",
X"0d02b305",
X"33028405",
X"b7053302",
X"8805ba05",
X"22595959",
X"800b8c3d",
X"348c3dfc",
X"05568055",
X"80547653",
X"77527851",
X"fbf23f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f33d",
X"0d7f6264",
X"028c0580",
X"c2052272",
X"22811533",
X"425f415e",
X"59598078",
X"237d5378",
X"33528151",
X"ffa03f83",
X"c0800881",
X"ff065675",
X"802e8638",
X"755481ad",
X"3983c8bc",
X"08a81133",
X"821b3370",
X"862a7081",
X"0673982b",
X"5351575c",
X"56577980",
X"25833881",
X"5673762e",
X"873881f0",
X"54818239",
X"818c1733",
X"7081ff06",
X"79227d71",
X"31902b70",
X"902c7009",
X"709f2c72",
X"06705252",
X"53515357",
X"57547574",
X"24833875",
X"55748480",
X"8029fc80",
X"80057090",
X"2c515574",
X"ff2e9438",
X"83c8bc08",
X"81801133",
X"5154737c",
X"7081055e",
X"34db3977",
X"22760554",
X"73782379",
X"09709f2a",
X"70810682",
X"1c3381bf",
X"0671862b",
X"07515151",
X"5473821a",
X"347c7626",
X"8a387722",
X"547a7426",
X"febb3880",
X"547383c0",
X"800c8f3d",
X"0d04f93d",
X"0d7a5780",
X"0b893d23",
X"893dfc05",
X"53765279",
X"51f8da3f",
X"83c08008",
X"81ff0670",
X"57557496",
X"387c547b",
X"53883d22",
X"527651fd",
X"e53f83c0",
X"800881ff",
X"06567583",
X"c0800c89",
X"3d0d04f0",
X"3d0d6266",
X"02880580",
X"ce052241",
X"5d5e8002",
X"840580d2",
X"05227f81",
X"0533ff11",
X"5a5d5a5d",
X"81da5876",
X"bf2680e9",
X"3878802e",
X"80e1387a",
X"58787b27",
X"83387858",
X"821e3370",
X"872a585a",
X"76923d34",
X"923dfc05",
X"5677557b",
X"547e537d",
X"33528251",
X"f8de3f83",
X"c0800881",
X"ff065d80",
X"0b923d33",
X"585a7680",
X"2e833881",
X"5a821e33",
X"80ff067a",
X"872b0757",
X"76821f34",
X"7c913878",
X"78317083",
X"ffff0679",
X"1e5e5a57",
X"ff9b397c",
X"587783c0",
X"800c923d",
X"0d04f83d",
X"0d7b0284",
X"05b20522",
X"5858800b",
X"8a3d238a",
X"3dfc0553",
X"77527a51",
X"f6f73f83",
X"c0800881",
X"ff067057",
X"55749638",
X"7d547653",
X"893d2252",
X"7751feaf",
X"3f83c080",
X"0881ff06",
X"567583c0",
X"800c8a3d",
X"0d04ec3d",
X"0d666e02",
X"880580df",
X"0533028c",
X"0580e305",
X"33029005",
X"80e70533",
X"02940580",
X"eb053302",
X"980580ee",
X"05224143",
X"415f5c40",
X"570280f2",
X"0522963d",
X"23963df0",
X"05538417",
X"70537752",
X"59f6863f",
X"83c08008",
X"81ff0658",
X"7781e538",
X"777a8180",
X"06584080",
X"77258338",
X"81407994",
X"3d347b02",
X"840580c9",
X"05347c02",
X"840580ca",
X"05347d02",
X"840580cb",
X"05347a95",
X"3d347a88",
X"2a577602",
X"840580cd",
X"0534953d",
X"22577602",
X"840580ce",
X"05347688",
X"2a577602",
X"840580cf",
X"05347792",
X"3d34963d",
X"ec115757",
X"8855f417",
X"54923d22",
X"53775277",
X"51f6953f",
X"83c08008",
X"81ff0658",
X"7780ed38",
X"7e802e80",
X"cb38923d",
X"22790858",
X"587f802e",
X"9c387681",
X"80800779",
X"0c7e5496",
X"3dfc0553",
X"7783ffff",
X"06527851",
X"f9fc3f99",
X"39768280",
X"8007790c",
X"7e54953d",
X"22537783",
X"ffff0652",
X"7851fc8f",
X"3f83c080",
X"0881ff06",
X"58779d38",
X"923d2253",
X"80527f30",
X"70802584",
X"71315351",
X"57f9873f",
X"83c08008",
X"81ff0658",
X"7783c080",
X"0c963d0d",
X"04f63d0d",
X"7c028405",
X"b705335b",
X"5b805880",
X"57805680",
X"55795485",
X"5380527a",
X"51fda33f",
X"83c08008",
X"81ff0659",
X"78853879",
X"871c3478",
X"83c0800c",
X"8c3d0d04",
X"f93d0d02",
X"a7053302",
X"8405ab05",
X"33028805",
X"af053358",
X"5957800b",
X"83c8cb33",
X"54547274",
X"2e9f3881",
X"147081ff",
X"06555373",
X"8f2681b6",
X"387381c4",
X"2983c8c8",
X"05831133",
X"515372e3",
X"387381c4",
X"2983c8c4",
X"0555800b",
X"87163476",
X"88163475",
X"8a163477",
X"89163480",
X"750c83c8",
X"bc088c16",
X"0c800b84",
X"1634880b",
X"85163480",
X"0b861634",
X"841508ff",
X"a1ff06a0",
X"80078416",
X"0c811470",
X"81ff0653",
X"537451fe",
X"bc3f83c0",
X"800881ff",
X"06705553",
X"7280cd38",
X"8a397308",
X"750c7254",
X"80c23972",
X"81d2b455",
X"5681d2b4",
X"08802eb2",
X"38758429",
X"14700876",
X"53700851",
X"5454722d",
X"83c08008",
X"81ff0653",
X"72802ece",
X"38811670",
X"81ff0681",
X"d2b47184",
X"29115356",
X"57537208",
X"d0388054",
X"7383c080",
X"0c893d0d",
X"04f93d0d",
X"7957800b",
X"84180883",
X"c8bc0c58",
X"f0883f88",
X"170883c0",
X"80082783",
X"ed38effa",
X"3f83c080",
X"08810588",
X"180c83c8",
X"bc08b811",
X"337081ff",
X"06515154",
X"73812ea4",
X"38738124",
X"88387378",
X"2e8a38b8",
X"3973822e",
X"9538b139",
X"763381f0",
X"06547390",
X"2ea63891",
X"7734a139",
X"73587633",
X"81f00654",
X"73902e09",
X"81069138",
X"efa83f83",
X"c0800881",
X"c8058c18",
X"0ca07734",
X"80567581",
X"c42983c8",
X"cb113355",
X"5573802e",
X"aa3883c8",
X"c4157008",
X"56547480",
X"2e9d3888",
X"1508802e",
X"96388c14",
X"0883c8bc",
X"082e0981",
X"06893873",
X"51881508",
X"54732d81",
X"167081ff",
X"0657548f",
X"7627ffba",
X"38763354",
X"73b02e81",
X"993873b0",
X"248f3873",
X"912eab38",
X"73a02e80",
X"f53882a6",
X"397380d0",
X"2e81e438",
X"7380d024",
X"8b387380",
X"c02e8199",
X"38828f39",
X"7381802e",
X"81fb3882",
X"85398056",
X"7581c429",
X"83c8c811",
X"83113356",
X"59557380",
X"2ea83883",
X"c8c41570",
X"08565474",
X"802e9b38",
X"8c140883",
X"c8bc082e",
X"0981068e",
X"38735184",
X"15085473",
X"2d800b83",
X"19348116",
X"7081ff06",
X"57548f76",
X"27ffb938",
X"92773481",
X"b539edc2",
X"3f8c1708",
X"83c08008",
X"2781a738",
X"b0773481",
X"a13983c8",
X"bc085480",
X"0b8c1534",
X"83c8bc08",
X"54840b88",
X"153480c0",
X"7734ed96",
X"3f83c080",
X"08b2058c",
X"180c80fa",
X"39ed873f",
X"8c170883",
X"c0800827",
X"80ec3883",
X"c8bc0854",
X"810b8c15",
X"3483c8bc",
X"0854800b",
X"88153483",
X"c8bc0854",
X"880ba015",
X"34ecdb3f",
X"83c08008",
X"94058c18",
X"0c80d077",
X"34bc3983",
X"c8bc08a0",
X"11337083",
X"2a708106",
X"51515555",
X"73802ea6",
X"38880ba0",
X"1634ecae",
X"3f8c1708",
X"83c08008",
X"279438ff",
X"8077348e",
X"39775380",
X"528051fa",
X"8b3fff90",
X"773483c8",
X"bc08a011",
X"3370832a",
X"70810651",
X"51555573",
X"802e8638",
X"880ba016",
X"34893d0d",
X"04f63d0d",
X"02b30533",
X"028405b7",
X"05335b5b",
X"800b83c8",
X"c8708412",
X"72745d59",
X"575b5856",
X"83153353",
X"72802e80",
X"f3387333",
X"537a732e",
X"09810680",
X"e7388114",
X"33537973",
X"2e098106",
X"80da3880",
X"557481c4",
X"2983c8cc",
X"05703383",
X"1b335855",
X"5373762e",
X"0981068a",
X"38811333",
X"527351ff",
X"9c3f8115",
X"7081ff06",
X"56538f75",
X"27d33880",
X"0b83c8c4",
X"19700856",
X"54557375",
X"2e913872",
X"51841408",
X"53722d83",
X"c0800881",
X"ff065580",
X"0b831834",
X"7453a039",
X"811681c4",
X"1981c417",
X"81c41781",
X"c41d81c4",
X"1c5c5d57",
X"5759568f",
X"7625fee8",
X"38805372",
X"83c0800c",
X"8c3d0d04",
X"f83d0d02",
X"ae05227d",
X"59578056",
X"81558054",
X"86538180",
X"527a51f5",
X"953f83c0",
X"800881ff",
X"0683c080",
X"0c8a3d0d",
X"04f73d0d",
X"02b20522",
X"028405b7",
X"0533605a",
X"5b578056",
X"82557954",
X"86538180",
X"527b51f4",
X"e53f83c0",
X"800881ff",
X"0683c080",
X"0c8b3d0d",
X"04f83d0d",
X"02af0533",
X"59805880",
X"57805680",
X"55785489",
X"5380527a",
X"51f4bb3f",
X"83c08008",
X"81ff0683",
X"c0800c8a",
X"3d0d0483",
X"c08c0802",
X"83c08c0c",
X"fd3d0d80",
X"5383c08c",
X"088c0508",
X"5283c08c",
X"08880508",
X"5183d43f",
X"83c08008",
X"7083c080",
X"0c54853d",
X"0d83c08c",
X"0c0483c0",
X"8c080283",
X"c08c0cfd",
X"3d0d8153",
X"83c08c08",
X"8c050852",
X"83c08c08",
X"88050851",
X"83a13f83",
X"c0800870",
X"83c0800c",
X"54853d0d",
X"83c08c0c",
X"0483c08c",
X"080283c0",
X"8c0cf93d",
X"0d800b83",
X"c08c08fc",
X"050c83c0",
X"8c088805",
X"088025b9",
X"3883c08c",
X"08880508",
X"3083c08c",
X"0888050c",
X"800b83c0",
X"8c08f405",
X"0c83c08c",
X"08fc0508",
X"8a38810b",
X"83c08c08",
X"f4050c83",
X"c08c08f4",
X"050883c0",
X"8c08fc05",
X"0c83c08c",
X"088c0508",
X"8025b938",
X"83c08c08",
X"8c050830",
X"83c08c08",
X"8c050c80",
X"0b83c08c",
X"08f0050c",
X"83c08c08",
X"fc05088a",
X"38810b83",
X"c08c08f0",
X"050c83c0",
X"8c08f005",
X"0883c08c",
X"08fc050c",
X"805383c0",
X"8c088c05",
X"085283c0",
X"8c088805",
X"085181df",
X"3f83c080",
X"087083c0",
X"8c08f805",
X"0c5483c0",
X"8c08fc05",
X"08802e90",
X"3883c08c",
X"08f80508",
X"3083c08c",
X"08f8050c",
X"83c08c08",
X"f8050870",
X"83c0800c",
X"54893d0d",
X"83c08c0c",
X"0483c08c",
X"080283c0",
X"8c0cfb3d",
X"0d800b83",
X"c08c08fc",
X"050c83c0",
X"8c088805",
X"08802599",
X"3883c08c",
X"08880508",
X"3083c08c",
X"0888050c",
X"810b83c0",
X"8c08fc05",
X"0c83c08c",
X"088c0508",
X"80259038",
X"83c08c08",
X"8c050830",
X"83c08c08",
X"8c050c81",
X"5383c08c",
X"088c0508",
X"5283c08c",
X"08880508",
X"51bd3f83",
X"c0800870",
X"83c08c08",
X"f8050c54",
X"83c08c08",
X"fc050880",
X"2e903883",
X"c08c08f8",
X"05083083",
X"c08c08f8",
X"050c83c0",
X"8c08f805",
X"087083c0",
X"800c5487",
X"3d0d83c0",
X"8c0c0483",
X"c08c0802",
X"83c08c0c",
X"fd3d0d81",
X"0b83c08c",
X"08fc050c",
X"800b83c0",
X"8c08f805",
X"0c83c08c",
X"088c0508",
X"83c08c08",
X"88050827",
X"b93883c0",
X"8c08fc05",
X"08802eae",
X"38800b83",
X"c08c088c",
X"050824a2",
X"3883c08c",
X"088c0508",
X"1083c08c",
X"088c050c",
X"83c08c08",
X"fc050810",
X"83c08c08",
X"fc050cff",
X"b83983c0",
X"8c08fc05",
X"08802e80",
X"e13883c0",
X"8c088c05",
X"0883c08c",
X"08880508",
X"26ad3883",
X"c08c0888",
X"050883c0",
X"8c088c05",
X"083183c0",
X"8c088805",
X"0c83c08c",
X"08f80508",
X"83c08c08",
X"fc050807",
X"83c08c08",
X"f8050c83",
X"c08c08fc",
X"0508812a",
X"83c08c08",
X"fc050c83",
X"c08c088c",
X"0508812a",
X"83c08c08",
X"8c050cff",
X"953983c0",
X"8c089005",
X"08802e93",
X"3883c08c",
X"08880508",
X"7083c08c",
X"08f4050c",
X"51913983",
X"c08c08f8",
X"05087083",
X"c08c08f4",
X"050c5183",
X"c08c08f4",
X"050883c0",
X"800c853d",
X"0d83c08c",
X"0c0483c0",
X"8c080283",
X"c08c0cff",
X"3d0d800b",
X"83c08c08",
X"fc050c83",
X"c08c0888",
X"05088106",
X"ff117009",
X"7083c08c",
X"088c0508",
X"0683c08c",
X"08fc0508",
X"1183c08c",
X"08fc050c",
X"83c08c08",
X"88050881",
X"2a83c08c",
X"0888050c",
X"83c08c08",
X"8c050810",
X"83c08c08",
X"8c050c51",
X"51515183",
X"c08c0888",
X"0508802e",
X"8438ffab",
X"3983c08c",
X"08fc0508",
X"7083c080",
X"0c51833d",
X"0d83c08c",
X"0c04fc3d",
X"0d767079",
X"7b555555",
X"558f7227",
X"8c387275",
X"07830651",
X"70802ea9",
X"38ff1252",
X"71ff2e98",
X"38727081",
X"05543374",
X"70810556",
X"34ff1252",
X"71ff2e09",
X"8106ea38",
X"7483c080",
X"0c863d0d",
X"04745172",
X"70840554",
X"08717084",
X"05530c72",
X"70840554",
X"08717084",
X"05530c72",
X"70840554",
X"08717084",
X"05530c72",
X"70840554",
X"08717084",
X"05530cf0",
X"1252718f",
X"26c93883",
X"72279538",
X"72708405",
X"54087170",
X"8405530c",
X"fc125271",
X"8326ed38",
X"7054ff81",
X"39000000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00002d58",
X"00002d99",
X"00002db9",
X"00002ddd",
X"00002de9",
X"000038c4",
X"00004108",
X"000041c1",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3a00",
X"0c0c3b00",
X"0a0a0008",
X"0b0b0008",
X"07070008",
X"0a0b4300",
X"080b4200",
X"04044500",
X"05054400",
X"06060004",
X"08080004",
X"09090004",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"00004e4d",
X"00005154",
X"00004f60",
X"00005154",
X"00004f9d",
X"00004fee",
X"0000502d",
X"00005036",
X"00005154",
X"00005154",
X"00005154",
X"00005154",
X"0000503f",
X"00005047",
X"0000504e",
X"00005254",
X"0000534d",
X"00005461",
X"00005757",
X"00005772",
X"0000575e",
X"00005772",
X"00005779",
X"00005784",
X"0000578b",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"31364b00",
X"556e6b6e",
X"6f776e20",
X"74797065",
X"206f6620",
X"63617274",
X"72696467",
X"65210000",
X"41353200",
X"43415200",
X"42494e00",
X"31366b20",
X"63617274",
X"20747970",
X"65000000",
X"4c656674",
X"20666f72",
X"206f6e65",
X"20636869",
X"70000000",
X"52696768",
X"7420666f",
X"72207477",
X"6f206368",
X"69700000",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a257300",
X"45786974",
X"00000000",
X"35323030",
X"2e726f6d",
X"00000000",
X"524f4d00",
X"4d454d00",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"00000000",
X"00006794",
X"000065e8",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"35323030",
X"00000000",
X"2f617461",
X"72353230",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
