
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f2",
X"80738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80f5",
X"b40c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580ef",
X"bf2d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580eefe",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80da8a04",
X"fd3d0d75",
X"705254ad",
X"b13f83e0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83e0",
X"8008732e",
X"a13883e0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183e0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83e2c008",
X"248a38b4",
X"823fff0b",
X"83e2c00c",
X"800b83e0",
X"800c04ff",
X"3d0d7352",
X"83e09c08",
X"722e8d38",
X"d93f7151",
X"96993f71",
X"83e09c0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"558154bc",
X"15088191",
X"387451cf",
X"3f795880",
X"7a2580f7",
X"3883e2f0",
X"0870892a",
X"5783ff06",
X"78848072",
X"31565657",
X"73782583",
X"38735575",
X"83e2c008",
X"2e8438ff",
X"893f83e2",
X"c0088025",
X"a6387589",
X"2b5198dc",
X"3f83e2f0",
X"088f3dfc",
X"11555c54",
X"8152f81b",
X"5196c63f",
X"761483e2",
X"f00c7583",
X"e2c00c74",
X"53765278",
X"51b2b33f",
X"83e08008",
X"83e2f008",
X"1683e2f0",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8b3861",
X"7a710c54",
X"75547580",
X"2e833881",
X"547383e0",
X"800c8e3d",
X"0d04fc3d",
X"0dfe9b3f",
X"7651feaf",
X"3f863dfc",
X"05537852",
X"775195e9",
X"3f797571",
X"0c5483e0",
X"80085483",
X"e0800880",
X"2e833881",
X"547383e0",
X"800c863d",
X"0d04fe3d",
X"0d7583e2",
X"c0085353",
X"80722489",
X"3871732e",
X"8438fdd6",
X"3f7451fd",
X"ea3f7251",
X"97ae3f83",
X"e0800852",
X"83e08008",
X"802e8338",
X"81527183",
X"e0800c84",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"e0800c51",
X"823d0d04",
X"80c40b83",
X"e0800c04",
X"fd3d0d75",
X"77715470",
X"535553a9",
X"893f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfceb3f",
X"735193ab",
X"3f7383e0",
X"9c0c83e0",
X"80085383",
X"e0800880",
X"2e833881",
X"537283e0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcbf3f",
X"72802ea5",
X"38bc1308",
X"527351a8",
X"933f83e0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"e0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83e0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83e2c0",
X"0c7483e0",
X"a00c7583",
X"e2bc0cae",
X"e73f83e0",
X"800881ff",
X"06528153",
X"71993883",
X"e2d8518e",
X"943f83e0",
X"80085283",
X"e0800880",
X"2e833872",
X"52715372",
X"83e0800c",
X"843d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"51a6843f",
X"83e08008",
X"557483e0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"e0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283e2bc",
X"085180de",
X"813f83e0",
X"800857f9",
X"e13f7952",
X"83e2c451",
X"95b73f83",
X"e0800854",
X"805383e0",
X"8008732e",
X"09810682",
X"833883e0",
X"a0080b0b",
X"80f3b453",
X"705256a5",
X"c13f0b0b",
X"80f3b452",
X"80c01651",
X"a5b43f75",
X"bc170c73",
X"82c0170c",
X"810b82c4",
X"170c810b",
X"82c8170c",
X"7382cc17",
X"0cff1782",
X"d0175557",
X"81913983",
X"e0ac3370",
X"822a7081",
X"06515455",
X"72818038",
X"74812a81",
X"06587780",
X"f6387484",
X"2a810682",
X"c4150c83",
X"e0ac3381",
X"0682c815",
X"0c795273",
X"51a4db3f",
X"7351a4f2",
X"3f83e080",
X"081453af",
X"73708105",
X"553472bc",
X"150c83e0",
X"ad527251",
X"a4bc3f83",
X"e0a40882",
X"c0150c83",
X"e0ba5280",
X"c01451a4",
X"a93f7880",
X"2e8d3873",
X"51782d83",
X"e0800880",
X"2e993877",
X"82cc150c",
X"75802e86",
X"387382cc",
X"170c7382",
X"d015ff19",
X"59555676",
X"802e9b38",
X"83e0a452",
X"83e2c451",
X"94ad3f83",
X"e080088a",
X"3883e0ad",
X"335372fe",
X"d2387880",
X"2e893883",
X"e0a00851",
X"fcb83f83",
X"e0a00853",
X"7283e080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb53f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f690",
X"3f83e080",
X"08745387",
X"3d705355",
X"55f6b03f",
X"f7903f73",
X"51d33f63",
X"53745283",
X"e0800851",
X"fab83f92",
X"3d0d0471",
X"83e0800c",
X"0480c012",
X"83e0800c",
X"04803d0d",
X"7282c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"e0800c51",
X"823d0d04",
X"f93d0d79",
X"83e09008",
X"57578177",
X"27819638",
X"76881708",
X"27818e38",
X"75335574",
X"822e8938",
X"74832eb3",
X"3880fe39",
X"74547610",
X"83fe0653",
X"76882a8c",
X"17080552",
X"893dfc05",
X"51a9953f",
X"83e08008",
X"80df3802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d13984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"51a8e53f",
X"83e08008",
X"b038029f",
X"05330284",
X"059e0533",
X"71982b71",
X"902b0702",
X"8c059d05",
X"3370882b",
X"72078d3d",
X"337180ff",
X"fffe8006",
X"07515253",
X"57585683",
X"39815574",
X"83e0800c",
X"893d0d04",
X"fb3d0d83",
X"e09008fe",
X"19881208",
X"fe055556",
X"54805674",
X"73278d38",
X"82143375",
X"71299416",
X"08055753",
X"7583e080",
X"0c873d0d",
X"04fc3d0d",
X"7652800b",
X"83e09008",
X"70335152",
X"5370832e",
X"09810691",
X"38951233",
X"94133371",
X"982b7190",
X"2b075555",
X"519b1233",
X"9a133371",
X"882b0774",
X"0783e080",
X"0c55863d",
X"0d04fc3d",
X"0d7683e0",
X"90085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"fed63f83",
X"e0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183e080",
X"0c863d0d",
X"04fa3d0d",
X"7883e090",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fcb13f",
X"81527183",
X"e0800827",
X"a8388352",
X"83e08008",
X"88170827",
X"9c3883e0",
X"80088c16",
X"0c83e080",
X"0851fdbc",
X"3f83e080",
X"0890160c",
X"73752380",
X"527183e0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585e5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"9f269138",
X"7a51fdd2",
X"3f83e080",
X"0856807d",
X"34838139",
X"933d841c",
X"08705859",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"3880705a",
X"5c887f08",
X"5f5a7b81",
X"1d7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535e57",
X"557480e7",
X"3876ae2e",
X"09810683",
X"38815578",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675bb",
X"3888598b",
X"5affab39",
X"76982b55",
X"74802587",
X"3880f190",
X"173357ff",
X"9f175574",
X"99268938",
X"e0177081",
X"ff065855",
X"78811a70",
X"81ff0672",
X"1b535b57",
X"55767534",
X"fef8397b",
X"1e7f0c80",
X"5576a026",
X"83388155",
X"748b1934",
X"7a51fc82",
X"3f83e080",
X"0880f538",
X"a0547a22",
X"70852b83",
X"e0065455",
X"901b0852",
X"7c51a3a0",
X"3f83e080",
X"085783e0",
X"80088181",
X"387c3355",
X"74802e80",
X"f4388b1d",
X"3370832a",
X"70810651",
X"565674b4",
X"388b7d84",
X"1d0883e0",
X"8008595b",
X"5b58ff18",
X"5877ff2e",
X"9a387970",
X"81055b33",
X"79708105",
X"5b337171",
X"31525656",
X"75802ee2",
X"38863975",
X"802e9638",
X"7a51fbe5",
X"3fff8639",
X"83e08008",
X"5683e080",
X"08b63883",
X"39765684",
X"1b088b11",
X"33515574",
X"a7388b1d",
X"3370842a",
X"70810651",
X"56567489",
X"38835694",
X"39815690",
X"397c51fa",
X"943f83e0",
X"8008881c",
X"0cfd8139",
X"7583e080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"51a1e53f",
X"835683e0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"51a1b93f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"7651a190",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583e080",
X"0c8a3d0d",
X"04eb3d0d",
X"675a800b",
X"83e0900c",
X"a0b23f83",
X"e0800881",
X"06558256",
X"7483ef38",
X"7475538f",
X"3d705357",
X"59feca3f",
X"83e08008",
X"81ff0657",
X"76812e09",
X"810680d4",
X"38905483",
X"be537452",
X"7551a0a4",
X"3f83e080",
X"0880c938",
X"8f3d3355",
X"74802e80",
X"c93802bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"33710770",
X"587b575e",
X"525e5759",
X"57fdee3f",
X"83e08008",
X"81ff0657",
X"76832e09",
X"81068638",
X"815682f2",
X"3976802e",
X"86388656",
X"82e839a4",
X"548d5378",
X"5275519f",
X"bb3f8156",
X"83e08008",
X"82d43802",
X"be053302",
X"8405bd05",
X"3371882b",
X"07595d77",
X"ab380280",
X"ce053302",
X"840580cd",
X"05337198",
X"2b71902b",
X"07973d33",
X"70882b72",
X"07029405",
X"80cb0533",
X"71075452",
X"5e575956",
X"02b70533",
X"78712902",
X"8805b605",
X"33028c05",
X"b5053371",
X"882b0770",
X"1d707f8c",
X"050c5f59",
X"57595d8e",
X"3d33821b",
X"3402b905",
X"33903d33",
X"71882b07",
X"5a5c7884",
X"1b2302bb",
X"05330284",
X"05ba0533",
X"71882b07",
X"565c74ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"07515253",
X"575e5c74",
X"76317831",
X"79842a90",
X"3d335471",
X"71315356",
X"5680cee6",
X"3f83e080",
X"08820570",
X"881c0c83",
X"e08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83e0900c",
X"80567583",
X"e0800c97",
X"3d0d04e9",
X"3d0d83e0",
X"90085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e53f83e0",
X"80085483",
X"e0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f489",
X"3f83e080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383e080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83e09008",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0e93f",
X"83e08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"833f83e0",
X"80085583",
X"e0800880",
X"2eff8938",
X"83e08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"5199e13f",
X"83e08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83e0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83e09008",
X"55568555",
X"73802e81",
X"e3388114",
X"33810653",
X"84557280",
X"2e81d538",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b9388214",
X"3370892b",
X"56537680",
X"2eb73874",
X"52ff1651",
X"80c9e73f",
X"83e08008",
X"ff187654",
X"70535853",
X"80c9d73f",
X"83e08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed63f83",
X"e0800853",
X"810b83e0",
X"8008278b",
X"38881408",
X"83e08008",
X"26883880",
X"0b811534",
X"b03983e0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc53f",
X"83e08008",
X"8c3883e0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683e0",
X"800805a8",
X"150c8055",
X"7483e080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83e09008",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1cf3f",
X"83e08008",
X"5583e080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef5",
X"3f83e080",
X"0888170c",
X"7551efa6",
X"3f83e080",
X"08557483",
X"e0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683e0",
X"9008802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f53f83e0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"95ea3f83",
X"e0800841",
X"83e08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"eddf3f83",
X"e0800841",
X"83e08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"8d903f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f03f83e0",
X"80088332",
X"70307072",
X"079f2c83",
X"e0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"8b9c3f75",
X"83e0800c",
X"9e3d0d04",
X"f93d0d80",
X"0b83e080",
X"0c893d0d",
X"04fc3d0d",
X"76705255",
X"8b983f83",
X"e0800815",
X"ff055473",
X"752e8e38",
X"73335372",
X"ae2e8638",
X"ff1454ef",
X"39775281",
X"14518ab0",
X"3f83e080",
X"08307083",
X"e0800807",
X"802583e0",
X"800c5386",
X"3d0d04fc",
X"3d0d7670",
X"5255e7e3",
X"3f83e080",
X"08548153",
X"83e08008",
X"80c13874",
X"51e7a63f",
X"83e08008",
X"80f3c453",
X"83e08008",
X"5253ff91",
X"3f83e080",
X"08a13880",
X"f3c85272",
X"51ff823f",
X"83e08008",
X"923880f3",
X"cc527251",
X"fef33f83",
X"e0800880",
X"2e833881",
X"54735372",
X"83e0800c",
X"863d0d04",
X"fd3d0d75",
X"705254e7",
X"823f8153",
X"83e08008",
X"98387351",
X"e6cb3f83",
X"e3880852",
X"83e08008",
X"51feba3f",
X"83e08008",
X"537283e0",
X"800c853d",
X"0d04df3d",
X"0da43d08",
X"70525edc",
X"f03f83e0",
X"80083395",
X"3d565473",
X"963880f8",
X"b8527451",
X"89903f9a",
X"397d5278",
X"51dff13f",
X"84cf397d",
X"51dcd63f",
X"83e08008",
X"527451dc",
X"863f8043",
X"80428041",
X"804083e3",
X"90085294",
X"3d70525d",
X"e2d93f83",
X"e0800859",
X"800b83e0",
X"8008555b",
X"83e08008",
X"7b2e9438",
X"811b7452",
X"5be5db3f",
X"83e08008",
X"5483e080",
X"08ee3880",
X"5aff5f79",
X"09709f2c",
X"7b065b54",
X"7a7a2484",
X"38ff1b5a",
X"f61a7009",
X"709f2c72",
X"067bff12",
X"5a5a5255",
X"55807525",
X"95387651",
X"e5a03f83",
X"e0800876",
X"ff185855",
X"57738024",
X"ed38747f",
X"2e8638a0",
X"d83f745f",
X"78ff1b70",
X"585d5880",
X"7a259538",
X"7751e4f6",
X"3f83e080",
X"0876ff18",
X"58555873",
X"8024ed38",
X"800b83e7",
X"c00c800b",
X"83e7e40c",
X"80f3d051",
X"8d8f3f81",
X"800b83e7",
X"e40c80f3",
X"d8518d81",
X"3fa80b83",
X"e7c00c76",
X"802e80e4",
X"3883e7c0",
X"08777932",
X"70307072",
X"07802570",
X"872b83e7",
X"e40c5156",
X"78535656",
X"e4ad3f83",
X"e0800880",
X"2e883880",
X"f3e0518c",
X"c83f7651",
X"e3ef3f83",
X"e0800852",
X"80f4ec51",
X"8cb73f76",
X"51e3f73f",
X"83e08008",
X"83e7c008",
X"55577574",
X"258638a8",
X"1656f739",
X"7583e7c0",
X"0c86f076",
X"24ff9838",
X"87980b83",
X"e7c00c77",
X"802eb138",
X"7751e3ad",
X"3f83e080",
X"08785255",
X"e3cd3f80",
X"f3e85483",
X"e080088d",
X"38873980",
X"763481d0",
X"3980f3e4",
X"54745373",
X"5280f3b8",
X"518bd63f",
X"805480f3",
X"c0518bcd",
X"3f811454",
X"73a82e09",
X"8106ef38",
X"868da051",
X"9cdd3f80",
X"52903d70",
X"525780c0",
X"ae3f8352",
X"765180c0",
X"a63f6281",
X"8f386180",
X"2e80fb38",
X"7b5473ff",
X"2e963878",
X"802e8189",
X"387851e2",
X"d13f83e0",
X"8008ff15",
X"5559e739",
X"78802e80",
X"f4387851",
X"e2cd3f83",
X"e0800880",
X"2efc8e38",
X"7851e295",
X"3f83e080",
X"085280f3",
X"b45183e3",
X"3f83e080",
X"08a3387c",
X"51859b3f",
X"83e08008",
X"5574ff16",
X"56548074",
X"25ae3874",
X"1d703355",
X"5673af2e",
X"fecd38e9",
X"397851e1",
X"d63f83e0",
X"8008527c",
X"5184d33f",
X"8f397f88",
X"29601005",
X"7a056105",
X"5afc9039",
X"62802efb",
X"d1388052",
X"7651bf87",
X"3fa33d0d",
X"04803d0d",
X"9088b833",
X"7081ff06",
X"70842a81",
X"32708106",
X"51515151",
X"70802e8d",
X"38a80b90",
X"88b834b8",
X"0b9088b8",
X"347083e0",
X"800c823d",
X"0d04803d",
X"0d9088b8",
X"337081ff",
X"0670852a",
X"81327081",
X"06515151",
X"5170802e",
X"8d38980b",
X"9088b834",
X"b80b9088",
X"b8347083",
X"e0800c82",
X"3d0d0493",
X"0b9088bc",
X"34ff0b90",
X"88a83404",
X"ff3d0d02",
X"8f053352",
X"800b9088",
X"bc348a51",
X"9aa53fdf",
X"3f80f80b",
X"9088a034",
X"800b9088",
X"8834fa12",
X"52719088",
X"8034800b",
X"90889834",
X"71908890",
X"349088b8",
X"52807234",
X"b8723483",
X"3d0d0480",
X"3d0d028b",
X"05335170",
X"9088b434",
X"febf3f83",
X"e0800880",
X"2ef63882",
X"3d0d0480",
X"3d0d8439",
X"a3fc3ffe",
X"d93f83e0",
X"8008802e",
X"f3389088",
X"b4337081",
X"ff0683e0",
X"800c5182",
X"3d0d0480",
X"3d0da30b",
X"9088bc34",
X"ff0b9088",
X"a8349088",
X"b851a871",
X"34b87134",
X"823d0d04",
X"803d0d90",
X"88bc3370",
X"81c00670",
X"30708025",
X"83e0800c",
X"51515182",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067083",
X"2a813270",
X"81065151",
X"51517080",
X"2ee838b0",
X"0b9088b8",
X"34b80b90",
X"88b83482",
X"3d0d0480",
X"3d0d9080",
X"ac088106",
X"83e0800c",
X"823d0d04",
X"fd3d0d75",
X"77545480",
X"73259438",
X"73708105",
X"55335280",
X"f3ec5187",
X"843fff13",
X"53e93985",
X"3d0d04fd",
X"3d0d7577",
X"53547333",
X"51708938",
X"71335170",
X"802ea138",
X"73337233",
X"52537271",
X"278538ff",
X"51943970",
X"73278538",
X"81518b39",
X"81148113",
X"5354d339",
X"80517083",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"54547233",
X"7081ff06",
X"52527080",
X"2ea33871",
X"81ff0681",
X"14ffbf12",
X"53545270",
X"99268938",
X"a0127081",
X"ff065351",
X"71747081",
X"055634d2",
X"39807434",
X"853d0d04",
X"ffbd3d0d",
X"80c63d08",
X"52a53d70",
X"5254ffb3",
X"3f80c73d",
X"0852853d",
X"705253ff",
X"a63f7252",
X"7351fedf",
X"3f80c53d",
X"0d04fe3d",
X"0d747653",
X"53717081",
X"05533351",
X"70737081",
X"05553470",
X"f038843d",
X"0d04fe3d",
X"0d745280",
X"72335253",
X"70732e8d",
X"38811281",
X"14713353",
X"545270f5",
X"387283e0",
X"800c843d",
X"0d04f63d",
X"0d7c7e60",
X"625a5d5b",
X"56805981",
X"55853974",
X"7a295574",
X"527551b7",
X"b13f83e0",
X"80087a27",
X"ee387480",
X"2e80dd38",
X"74527551",
X"b79c3f83",
X"e0800875",
X"53765254",
X"b7a03f83",
X"e080087a",
X"53755256",
X"b7843f83",
X"e0800879",
X"30707b07",
X"9f2a7077",
X"80240751",
X"51545572",
X"873883e0",
X"8008c538",
X"768118b0",
X"16555858",
X"8974258b",
X"38b71453",
X"7a853880",
X"d7145372",
X"78348119",
X"59ff9f39",
X"8077348c",
X"3d0d04f7",
X"3d0d7b7d",
X"7f620290",
X"05bb0533",
X"5759565a",
X"5ab05872",
X"8338a058",
X"75707081",
X"05523371",
X"59545590",
X"39807425",
X"8e38ff14",
X"77708105",
X"59335454",
X"72ef3873",
X"ff155553",
X"80732589",
X"38775279",
X"51782def",
X"39753375",
X"57537280",
X"2e903872",
X"52795178",
X"2d757081",
X"05573353",
X"ed398b3d",
X"0d04ee3d",
X"0d646669",
X"69707081",
X"0552335b",
X"4a5c5e5e",
X"76802e82",
X"f93876a5",
X"2e098106",
X"82e03880",
X"70416770",
X"70810552",
X"33714a59",
X"575f76b0",
X"2e098106",
X"8c387570",
X"81055733",
X"76485781",
X"5fd01756",
X"75892680",
X"da387667",
X"5c59805c",
X"9339778a",
X"2480c338",
X"7b8a2918",
X"7b708105",
X"5d335a5c",
X"d0197081",
X"ff065858",
X"897727a4",
X"38ff9f19",
X"7081ff06",
X"ffa91b5a",
X"51568576",
X"279238ff",
X"bf197081",
X"ff065156",
X"7585268a",
X"38c91958",
X"778025ff",
X"b9387a47",
X"7b407881",
X"ff065776",
X"80e42e80",
X"e5387680",
X"e424a738",
X"7680d82e",
X"81863876",
X"80d82490",
X"3876802e",
X"81cc3876",
X"a52e81b6",
X"3881b939",
X"7680e32e",
X"818c3881",
X"af397680",
X"f52e9b38",
X"7680f524",
X"8b387680",
X"f32e8181",
X"38819939",
X"7680f82e",
X"80ca3881",
X"8f39913d",
X"70555780",
X"538a5279",
X"841b7108",
X"535b56fc",
X"813f7655",
X"ab397984",
X"1b710894",
X"3d705b5b",
X"525b5675",
X"80258c38",
X"753056ad",
X"78340280",
X"c1055776",
X"5480538a",
X"527551fb",
X"d53f7755",
X"7e54b839",
X"913d7055",
X"7780d832",
X"70307080",
X"25565158",
X"56905279",
X"841b7108",
X"535b57fb",
X"b13f7555",
X"db397984",
X"1b831233",
X"545b5698",
X"3979841b",
X"7108575b",
X"5680547f",
X"537c527d",
X"51fc9c3f",
X"87397652",
X"7d517c2d",
X"66703358",
X"810547fd",
X"8339943d",
X"0d047283",
X"e0940c71",
X"83e0980c",
X"04fb3d0d",
X"883d7070",
X"84055208",
X"57547553",
X"83e09408",
X"5283e098",
X"0851fcc6",
X"3f873d0d",
X"04ff3d0d",
X"73700853",
X"51029305",
X"33723470",
X"08810571",
X"0c833d0d",
X"04fc3d0d",
X"873d8811",
X"557854bc",
X"c55351fc",
X"993f8052",
X"873d51d1",
X"3f863d0d",
X"04fc3d0d",
X"76557483",
X"e398082e",
X"af388053",
X"745187c1",
X"3f83e080",
X"0881ff06",
X"ff147081",
X"ff067230",
X"709f2a51",
X"52555354",
X"72802e84",
X"3871dd38",
X"73fe3874",
X"83e3980c",
X"863d0d04",
X"ff3d0dff",
X"0b83e398",
X"0c84a53f",
X"81518785",
X"3f83e080",
X"0881ff06",
X"5271ee38",
X"81d33f71",
X"83e0800c",
X"833d0d04",
X"fc3d0d76",
X"028405a2",
X"05220288",
X"05a60522",
X"7a545555",
X"55ff823f",
X"72802ea0",
X"3883e3ac",
X"14337570",
X"81055734",
X"81147083",
X"ffff06ff",
X"157083ff",
X"ff065652",
X"5552dd39",
X"800b83e0",
X"800c863d",
X"0d04fc3d",
X"0d76787a",
X"11565355",
X"80537174",
X"2e933872",
X"15517033",
X"83e3ac13",
X"34811281",
X"145452ea",
X"39800b83",
X"e0800c86",
X"3d0d04fd",
X"3d0d9054",
X"83e39808",
X"5186f43f",
X"83e08008",
X"81ff06ff",
X"15713071",
X"30707307",
X"9f2a729f",
X"2a065255",
X"52555372",
X"db38853d",
X"0d04803d",
X"0d83e3a4",
X"081083e3",
X"9c080790",
X"80a80c82",
X"3d0d0480",
X"0b83e3a4",
X"0ce43f04",
X"810b83e3",
X"a40cdb3f",
X"04ed3f04",
X"7183e3a0",
X"0c04803d",
X"0d8051f4",
X"3f810b83",
X"e3a40c81",
X"0b83e39c",
X"0cffbb3f",
X"823d0d04",
X"803d0d72",
X"30707407",
X"802583e3",
X"9c0c51ff",
X"a53f823d",
X"0d04803d",
X"0d028b05",
X"339080a4",
X"0c9080a8",
X"08708106",
X"515170f5",
X"389080a4",
X"087081ff",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d81ff51",
X"d13f83e0",
X"800881ff",
X"0683e080",
X"0c823d0d",
X"04803d0d",
X"73902b73",
X"079080b4",
X"0c823d0d",
X"0404fb3d",
X"0d780284",
X"059f0533",
X"70982b55",
X"57557280",
X"259b3875",
X"80ff0656",
X"805280f7",
X"51e03f83",
X"e0800881",
X"ff065473",
X"812680ff",
X"388051fe",
X"e73fffa2",
X"3f8151fe",
X"df3fff9a",
X"3f7551fe",
X"ed3f7498",
X"2a51fee6",
X"3f74902a",
X"7081ff06",
X"5253feda",
X"3f74882a",
X"7081ff06",
X"5253fece",
X"3f7481ff",
X"0651fec6",
X"3f815575",
X"80c02e09",
X"81068638",
X"8195558d",
X"397580c8",
X"2e098106",
X"84388187",
X"557451fe",
X"a53f8a55",
X"fec83f83",
X"e0800881",
X"ff067098",
X"2b545472",
X"80258c38",
X"ff157081",
X"ff065653",
X"74e23873",
X"83e0800c",
X"873d0d04",
X"fa3d0dfd",
X"c53f8051",
X"fdda3f8a",
X"54fe933f",
X"ff147081",
X"ff065553",
X"73f33873",
X"74535580",
X"c051fea6",
X"3f83e080",
X"0881ff06",
X"5473812e",
X"09810682",
X"9f3883aa",
X"5280c851",
X"fe8c3f83",
X"e0800881",
X"ff065372",
X"812e0981",
X"0681a838",
X"7454873d",
X"74115456",
X"fdc83f83",
X"e0800873",
X"34811470",
X"81ff0655",
X"53837427",
X"e538029a",
X"05335372",
X"812e0981",
X"0681d938",
X"029b0533",
X"5380ce90",
X"547281aa",
X"2e8d3881",
X"c73980e4",
X"518acc3f",
X"ff145473",
X"802e81b8",
X"38820a52",
X"81e951fd",
X"a53f83e0",
X"800881ff",
X"065372de",
X"38725280",
X"fa51fd92",
X"3f83e080",
X"0881ff06",
X"53728190",
X"38725473",
X"1653fcd6",
X"3f83e080",
X"08733481",
X"147081ff",
X"06555383",
X"7427e838",
X"873d3370",
X"862a7081",
X"06515454",
X"8c557280",
X"e3388455",
X"80de3974",
X"5281e951",
X"fccc3f83",
X"e0800881",
X"ff065382",
X"5581e956",
X"81732786",
X"38735580",
X"c15680ce",
X"90548a39",
X"80e45189",
X"be3fff14",
X"5473802e",
X"a9388052",
X"7551fc9a",
X"3f83e080",
X"0881ff06",
X"5372e138",
X"84805280",
X"d051fc86",
X"3f83e080",
X"0881ff06",
X"5372802e",
X"83388055",
X"7483e3a8",
X"348051fb",
X"873ffbc2",
X"3f883d0d",
X"04fb3d0d",
X"7754800b",
X"83e3a833",
X"70832a70",
X"81065155",
X"57557275",
X"2e098106",
X"85387389",
X"2b547352",
X"80d151fb",
X"bd3f83e0",
X"800881ff",
X"065372bd",
X"3882b8c0",
X"54fb833f",
X"83e08008",
X"81ff0653",
X"7281ff2e",
X"09810689",
X"38ff1454",
X"73e7389f",
X"397281fe",
X"2e098106",
X"963883e7",
X"ac5283e3",
X"ac51faed",
X"3ffad33f",
X"fad03f83",
X"39815580",
X"51fa893f",
X"fac43f74",
X"81ff0683",
X"e0800c87",
X"3d0d04fb",
X"3d0d7783",
X"e3ac5654",
X"8151f9ec",
X"3f83e3a8",
X"3370832a",
X"70810651",
X"54567285",
X"3873892b",
X"54735280",
X"d851fab6",
X"3f83e080",
X"0881ff06",
X"537280e4",
X"3881ff51",
X"f9d43f81",
X"fe51f9ce",
X"3f848053",
X"74708105",
X"563351f9",
X"c13fff13",
X"7083ffff",
X"06515372",
X"eb387251",
X"f9b03f72",
X"51f9ab3f",
X"f9d03f83",
X"e080089f",
X"0653a788",
X"5472852e",
X"8c389939",
X"80e45186",
X"f63fff14",
X"54f9b33f",
X"83e08008",
X"81ff2e84",
X"3873e938",
X"8051f8e4",
X"3ff99f3f",
X"800b83e0",
X"800c873d",
X"0d047183",
X"e7b00c88",
X"80800b83",
X"e7ac0c84",
X"80800b83",
X"e7b40c04",
X"fd3d0d77",
X"70175577",
X"05ff1a53",
X"5371ff2e",
X"94387370",
X"81055533",
X"51707370",
X"81055534",
X"ff1252e9",
X"39853d0d",
X"04fc3d0d",
X"87a68155",
X"743383e7",
X"b834a054",
X"83a08053",
X"83e7b008",
X"5283e7ac",
X"0851ffb8",
X"3fa05483",
X"a4805383",
X"e7b00852",
X"83e7ac08",
X"51ffa53f",
X"905483a8",
X"805383e7",
X"b0085283",
X"e7ac0851",
X"ff923fa0",
X"53805283",
X"e7b40883",
X"a0800551",
X"85ce3fa0",
X"53805283",
X"e7b40883",
X"a4800551",
X"85be3f90",
X"53805283",
X"e7b40883",
X"a8800551",
X"85ae3fff",
X"753483a0",
X"80548053",
X"83e7b008",
X"5283e7b4",
X"0851fecc",
X"3f80d080",
X"5483b080",
X"5383e7b0",
X"085283e7",
X"b40851fe",
X"b73f86e1",
X"3fa25480",
X"5383e7b4",
X"088c8005",
X"5280f6b0",
X"51fea13f",
X"860b87a8",
X"8334800b",
X"87a88234",
X"800b87a0",
X"9a34af0b",
X"87a09634",
X"bf0b87a0",
X"9734800b",
X"87a09834",
X"9f0b87a0",
X"9934800b",
X"87a09b34",
X"e00b87a8",
X"8934a20b",
X"87a88034",
X"830b87a4",
X"8f34820b",
X"87a88134",
X"863d0d04",
X"fd3d0d83",
X"a0805480",
X"5383e7b4",
X"085283e7",
X"b00851fd",
X"bf3f80d0",
X"805483b0",
X"805383e7",
X"b4085283",
X"e7b00851",
X"fdaa3fa0",
X"5483a080",
X"5383e7b4",
X"085283e7",
X"b00851fd",
X"973fa054",
X"83a48053",
X"83e7b408",
X"5283e7b0",
X"0851fd84",
X"3f905483",
X"a8805383",
X"e7b40852",
X"83e7b008",
X"51fcf13f",
X"83e7b833",
X"87a68134",
X"853d0d04",
X"803d0d90",
X"80900881",
X"0683e080",
X"0c823d0d",
X"04ff3d0d",
X"90809070",
X"0870fe06",
X"7607720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870812c",
X"810683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fd067610",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70822cbf",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"83067682",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870882c",
X"870683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"f1ff0676",
X"882b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"9008708b",
X"2cbf0683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f88fff",
X"06768b2b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70912cbf",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870fc",
X"87ffff06",
X"76912b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"992c8106",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870ffbf",
X"0a067699",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908080",
X"0870882c",
X"810683e0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"80087089",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8a2c8106",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708b2c81",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708c2c",
X"bf0683e0",
X"800c5182",
X"3d0d04fe",
X"3d0d7481",
X"e629872a",
X"9080a00c",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d848080",
X"53805288",
X"800a51ff",
X"b33f8180",
X"80538052",
X"82800a51",
X"c63f843d",
X"0d04803d",
X"0d8151fb",
X"fc3f7280",
X"2e903880",
X"51fdfe3f",
X"cd3f83e7",
X"bc3351fd",
X"f43f8151",
X"fc8d3f80",
X"51fc883f",
X"8051fbd9",
X"3f823d0d",
X"04fd3d0d",
X"75528054",
X"80ff7225",
X"8838810b",
X"ff801353",
X"54ffbf12",
X"51709926",
X"8638e012",
X"529e39ff",
X"9f125199",
X"71279538",
X"d012e013",
X"70545451",
X"89712788",
X"388f7327",
X"83388052",
X"73802e85",
X"38818012",
X"527181ff",
X"0683e080",
X"0c853d0d",
X"04803d0d",
X"84d8c051",
X"80717081",
X"05533470",
X"84e0c02e",
X"098106f0",
X"38823d0d",
X"04fe3d0d",
X"02970533",
X"51ff863f",
X"83e08008",
X"81ff0683",
X"e7c00854",
X"52807324",
X"9b3883e7",
X"e0081372",
X"83e7e408",
X"07535371",
X"733483e7",
X"c0088105",
X"83e7c00c",
X"843d0d04",
X"fa3d0d82",
X"800a1b55",
X"8057883d",
X"fc055479",
X"53745278",
X"51ffbbfe",
X"3f883d0d",
X"04fe3d0d",
X"83e7d808",
X"527451c2",
X"e23f83e0",
X"80088c38",
X"76537552",
X"83e7d808",
X"51c63f84",
X"3d0d04fe",
X"3d0d83e7",
X"d8085375",
X"527451ff",
X"bda03f83",
X"e080088d",
X"38775376",
X"5283e7d8",
X"0851ffa0",
X"3f843d0d",
X"04fe3d0d",
X"83e7d808",
X"51ffbc93",
X"3f83e080",
X"08818080",
X"2e098106",
X"8738b180",
X"80539b39",
X"83e7d808",
X"51ffbbf7",
X"3f83e080",
X"0880d080",
X"2e098106",
X"9238b1b0",
X"805383e0",
X"80085283",
X"e7d80851",
X"fed63f84",
X"3d0d0480",
X"3d0df9e2",
X"3f83e080",
X"08842980",
X"f6d40570",
X"0883e080",
X"0c51823d",
X"0d04ed3d",
X"0d804480",
X"43804280",
X"4180705a",
X"5bfdce3f",
X"800b83e7",
X"c00c800b",
X"83e7e40c",
X"80f4b851",
X"eaa73f81",
X"800b83e7",
X"e40c80f4",
X"bc51ea99",
X"3f80d00b",
X"83e7c00c",
X"7830707a",
X"07802570",
X"872b83e7",
X"e40c5155",
X"f8d33f83",
X"e0800852",
X"80f4c451",
X"e9f33f80",
X"f80b83e7",
X"c00c7881",
X"32703070",
X"72078025",
X"70872b83",
X"e7e40c51",
X"5656feef",
X"3f83e080",
X"085280f4",
X"d051e9c9",
X"3f81a00b",
X"83e7c00c",
X"78823270",
X"30707207",
X"80257087",
X"2b83e7e4",
X"0c515683",
X"e7d80852",
X"56ffb79d",
X"3f83e080",
X"085280f4",
X"d851e999",
X"3f81f00b",
X"83e7c00c",
X"810b83e7",
X"c45b5883",
X"e7c00882",
X"197a3270",
X"30707207",
X"80257087",
X"2b83e7e4",
X"0c51578e",
X"3d7055ff",
X"1b545757",
X"5799b13f",
X"79708405",
X"5b0851ff",
X"b6d33f74",
X"5483e080",
X"08537752",
X"80f4e051",
X"e8cb3fa8",
X"1783e7c0",
X"0c811858",
X"77852e09",
X"8106ffaf",
X"3883900b",
X"83e7c00c",
X"78873270",
X"30707207",
X"80257087",
X"2b83e7e4",
X"0c515656",
X"f7f73f80",
X"f4f05583",
X"e0800880",
X"2e8f3883",
X"e7d40851",
X"ffb5fe3f",
X"83e08008",
X"55745280",
X"f4f851e7",
X"f83f83e0",
X"0b83e7c0",
X"0c788832",
X"70307072",
X"07802570",
X"872b83e7",
X"e40c5157",
X"80f58452",
X"55e7d63f",
X"868da051",
X"f8f13f80",
X"52913d70",
X"52559cc3",
X"3f835274",
X"519cbc3f",
X"63557482",
X"fa386119",
X"59788025",
X"85387459",
X"90398879",
X"25853888",
X"59873978",
X"882682d9",
X"3878822b",
X"5580f390",
X"150804f5",
X"e43f83e0",
X"80086157",
X"5575812e",
X"09810689",
X"3883e080",
X"08105590",
X"3975ff2e",
X"09810688",
X"3883e080",
X"08812c55",
X"90752585",
X"38905588",
X"39748024",
X"83388155",
X"7451f5be",
X"3f828e39",
X"f5d03f83",
X"e0800861",
X"05557480",
X"25853880",
X"55883985",
X"75258338",
X"85557451",
X"f5c93f81",
X"ec396087",
X"3862802e",
X"81e33883",
X"e38c0883",
X"e3880cac",
X"f00b83e3",
X"900c83e7",
X"d80851d7",
X"8d3ffadd",
X"3f81c639",
X"60568076",
X"259838ac",
X"8f0b83e3",
X"900c83e7",
X"b8157008",
X"5255d6ee",
X"3f740852",
X"92397580",
X"25923883",
X"e7b81508",
X"51ffb3e7",
X"3f8052fd",
X"1951b839",
X"62802e81",
X"8c3883e7",
X"b8157008",
X"83e7c408",
X"720c83e7",
X"c40cfd1a",
X"70535155",
X"8bac3f83",
X"e0800856",
X"80518ba2",
X"3f83e080",
X"08527451",
X"87b93f75",
X"52805187",
X"b23f80d5",
X"39605580",
X"7525b638",
X"83e39408",
X"83e3880c",
X"acf00b83",
X"e3900c83",
X"e7d40851",
X"d5f83f83",
X"e7d40851",
X"d48e3f83",
X"e0800881",
X"ff067052",
X"55f4d73f",
X"74802e9d",
X"388155a1",
X"39748025",
X"943883e7",
X"d40851ff",
X"b2d93f80",
X"51f4bb3f",
X"84396287",
X"387a802e",
X"fa833880",
X"557483e0",
X"800c953d",
X"0d04fe3d",
X"0df4e73f",
X"83e08008",
X"802e8638",
X"8051818a",
X"39f4ec3f",
X"83e08008",
X"80fe38f5",
X"8c3f83e0",
X"8008802e",
X"b9388151",
X"f29b3f80",
X"51f4a23f",
X"ef8f3f80",
X"0b83e7c0",
X"0cf9ab3f",
X"83e08008",
X"53ff0b83",
X"e7c00cf0",
X"fb3f7280",
X"cb3883e7",
X"bc3351f3",
X"fc3f7251",
X"f1eb3f80",
X"c039f4b4",
X"3f83e080",
X"08802eb5",
X"388151f1",
X"d83f8051",
X"f3df3fee",
X"cc3fac8f",
X"0b83e390",
X"0c83e7c4",
X"0851d4aa",
X"3fff0b83",
X"e7c00cf0",
X"b73f83e7",
X"c4085280",
X"5185b03f",
X"8151f5a6",
X"3f843d0d",
X"04fc3d0d",
X"800b83e7",
X"bc348480",
X"805284a4",
X"808051ff",
X"b5923f83",
X"e0800880",
X"cd3888fb",
X"3f80f8a8",
X"51ffb9d1",
X"3f83e080",
X"0855b080",
X"805480c0",
X"805380f5",
X"8c5283e0",
X"800851f6",
X"fa3f83e7",
X"d8085380",
X"f59c5274",
X"51ffb49a",
X"3f83e080",
X"088438f7",
X"883f83e7",
X"bc3351f2",
X"d03f8151",
X"f4bc3f92",
X"ee3f8151",
X"f4b43f81",
X"51fdeb3f",
X"fa3983e0",
X"8c080283",
X"e08c0cfb",
X"3d0d0280",
X"f5a80b83",
X"e38c0c80",
X"f5ac0b83",
X"e3840c80",
X"f5b00b83",
X"e3940c83",
X"e08c08fc",
X"050c800b",
X"83e7c40b",
X"83e08c08",
X"f8050c83",
X"e08c08f4",
X"050cffb2",
X"e73f83e0",
X"80088605",
X"fc0683e0",
X"8c08f005",
X"0c0283e0",
X"8c08f005",
X"08310d83",
X"3d7083e0",
X"8c08f805",
X"08708405",
X"83e08c08",
X"f8050c0c",
X"51ffafaf",
X"3f83e08c",
X"08f40508",
X"810583e0",
X"8c08f405",
X"0c83e08c",
X"08f40508",
X"872e0981",
X"06ffab38",
X"84a88080",
X"51ebcf3f",
X"ff0b83e7",
X"c00c800b",
X"83e7e40c",
X"84d8c00b",
X"83e7e00c",
X"8151eef9",
X"3f8151ef",
X"9e3f8051",
X"ef993f81",
X"51efbf3f",
X"8151f094",
X"3f8251ef",
X"e23f8051",
X"f0b83f80",
X"51f0e23f",
X"80cfd552",
X"8051e0ae",
X"3ffda63f",
X"83e08c08",
X"fc05080d",
X"800b83e0",
X"800c873d",
X"0d83e08c",
X"0c04803d",
X"0d81ff51",
X"800b83e7",
X"f01234ff",
X"115170f4",
X"38823d0d",
X"04ff3d0d",
X"73703353",
X"51811133",
X"71347181",
X"1234833d",
X"0d04fb3d",
X"0d777956",
X"56807071",
X"55555271",
X"7525ac38",
X"72167033",
X"70147081",
X"ff065551",
X"51517174",
X"27893881",
X"127081ff",
X"06535171",
X"81147083",
X"ffff0655",
X"52547473",
X"24d63871",
X"83e0800c",
X"873d0d04",
X"fb3d0d77",
X"56d7f83f",
X"83e08008",
X"802ef638",
X"83ea8c08",
X"86057081",
X"ff065253",
X"d5fa3f81",
X"0b9088d4",
X"349088d4",
X"337081ff",
X"06515372",
X"8b38fac6",
X"3f8351f0",
X"963fea39",
X"80557416",
X"75822b54",
X"549088c0",
X"13337434",
X"81155574",
X"852e0981",
X"06e83881",
X"0b9088d4",
X"34753383",
X"e7f03481",
X"163383e7",
X"f1348216",
X"3383e7f2",
X"34831633",
X"83e7f334",
X"845283e7",
X"f051feba",
X"3f83e080",
X"0881ff06",
X"84173357",
X"5372762e",
X"0981068c",
X"38d6a13f",
X"83e08008",
X"802e9a38",
X"83ea8c08",
X"a82e0981",
X"06893886",
X"0b83ea8c",
X"0c8739a8",
X"0b83ea8c",
X"0c80e451",
X"ef913f87",
X"3d0d04f4",
X"3d0d7e60",
X"5955805d",
X"8075822b",
X"7183ea90",
X"120c83ea",
X"a4175b5b",
X"57767934",
X"77772e83",
X"b9387652",
X"7751ffad",
X"f53f8e3d",
X"fc055490",
X"5383e9f8",
X"527751ff",
X"adb03f7c",
X"5675902e",
X"09810683",
X"953883e9",
X"f851fd95",
X"3f83e9fa",
X"51fd8e3f",
X"83e9fc51",
X"fd873f76",
X"83ea880c",
X"7751ffaa",
X"fc3f0b0b",
X"80f3c852",
X"83e08008",
X"51cc9e3f",
X"83e08008",
X"812e0981",
X"0680d438",
X"7683eaa0",
X"0c820b83",
X"e9f834ff",
X"960b83e9",
X"f9347751",
X"ffadc03f",
X"83e08008",
X"5583e080",
X"08772588",
X"3883e080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"e9fa3474",
X"83e9fb34",
X"7683e9fc",
X"34ff800b",
X"83e9fd34",
X"81903983",
X"e9f83383",
X"e9f93371",
X"882b0756",
X"5b7483ff",
X"ff2e0981",
X"0680e838",
X"fe800b83",
X"eaa00c81",
X"0b83ea88",
X"0cff0b83",
X"e9f834ff",
X"0b83e9f9",
X"347751ff",
X"accd3f83",
X"e0800883",
X"eaa80c83",
X"e0800855",
X"83e08008",
X"80258838",
X"83e08008",
X"8f055574",
X"842c7083",
X"ffff0670",
X"882a5851",
X"557583e9",
X"fa347483",
X"e9fb3476",
X"83e9fc34",
X"ff800b83",
X"e9fd3481",
X"0b83ea87",
X"34a53974",
X"85962e09",
X"810680fe",
X"387583ea",
X"a00c7751",
X"ffac813f",
X"83ea8733",
X"83e08008",
X"07557483",
X"ea873483",
X"ea873381",
X"06557480",
X"2e833884",
X"5783e9fc",
X"3383e9fd",
X"3371882b",
X"07565c74",
X"81802e09",
X"8106a138",
X"83e9fa33",
X"83e9fb33",
X"71882b07",
X"565bad80",
X"75278738",
X"76820757",
X"9c397681",
X"07579639",
X"7482802e",
X"09810687",
X"38768307",
X"57873974",
X"81ff268a",
X"387783ea",
X"901b0c76",
X"79348e3d",
X"0d04803d",
X"0d728429",
X"83ea9005",
X"700883e0",
X"800c5182",
X"3d0d04fe",
X"3d0d800b",
X"83e9f40c",
X"800b83e9",
X"f00cff0b",
X"83e7ec0c",
X"a80b83ea",
X"8c0cae51",
X"d0c23f80",
X"0b83ea90",
X"54528073",
X"70840555",
X"0c811252",
X"71842e09",
X"8106ef38",
X"843d0d04",
X"fe3d0d74",
X"02840596",
X"05225353",
X"71802e96",
X"38727081",
X"05543351",
X"d0cd3fff",
X"127083ff",
X"ff065152",
X"e739843d",
X"0d04fe3d",
X"0d029205",
X"225382ac",
X"51eaa43f",
X"80c351d0",
X"aa3f8196",
X"51ea983f",
X"725283e7",
X"f051ffb4",
X"3f725283",
X"e7f051f8",
X"f13f83e0",
X"800881ff",
X"0651d087",
X"3f843d0d",
X"04ffb13d",
X"0d80d13d",
X"f80551f9",
X"9b3f83e9",
X"f4088105",
X"83e9f40c",
X"80cf3d33",
X"cf117081",
X"ff065156",
X"56748326",
X"88e23875",
X"8f06ff05",
X"567583e7",
X"ec082e9b",
X"38758326",
X"96387583",
X"e7ec0c75",
X"842983ea",
X"90057008",
X"53557551",
X"fa993f80",
X"762488be",
X"38758429",
X"83ea9005",
X"55740880",
X"2e88af38",
X"83e7ec08",
X"842983ea",
X"90057008",
X"02880582",
X"b9053352",
X"5b557480",
X"d22e84ac",
X"387480d2",
X"24903874",
X"bf2e9c38",
X"7480d02e",
X"81d13887",
X"ee397480",
X"d32e80cf",
X"387480d7",
X"2e81c038",
X"87dd3902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"5656cf83",
X"3f80c151",
X"cebd3ff6",
X"ed3f860b",
X"83e7f034",
X"815283e7",
X"f051cfe0",
X"3f8151fd",
X"e93f7489",
X"38860b83",
X"ea8c0c87",
X"39a80b83",
X"ea8c0cce",
X"d23f80c1",
X"51ce8c3f",
X"f6bc3f90",
X"0b83ea87",
X"33810656",
X"5674802e",
X"83389856",
X"83e9fc33",
X"83e9fd33",
X"71882b07",
X"56597481",
X"802e0981",
X"069c3883",
X"e9fa3383",
X"e9fb3371",
X"882b0756",
X"57ad8075",
X"278c3875",
X"81800756",
X"853975a0",
X"07567583",
X"e7f034ff",
X"0b83e7f1",
X"34e00b83",
X"e7f23480",
X"0b83e7f3",
X"34845283",
X"e7f051ce",
X"d73f8451",
X"869b3902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"5659cdc7",
X"3f7951ff",
X"a6d23f83",
X"e0800880",
X"2e8a3880",
X"ce51ccf3",
X"3f85f139",
X"80c151cc",
X"ea3fcddf",
X"3fcc943f",
X"83eaa008",
X"58837525",
X"9b3883e9",
X"fc3383e9",
X"fd337188",
X"2b07fc17",
X"71297a05",
X"8380055a",
X"51578d39",
X"74818029",
X"18ff8005",
X"58818057",
X"80567676",
X"2e9238cc",
X"c63f83e0",
X"800883e7",
X"f0173481",
X"1656eb39",
X"ccb53f83",
X"e0800881",
X"ff067753",
X"83e7f052",
X"56f4e73f",
X"83e08008",
X"81ff0655",
X"75752e09",
X"81068195",
X"389451e5",
X"e63fccaf",
X"3f80c151",
X"cbe93fcc",
X"de3f7752",
X"7951ffa4",
X"e53f805e",
X"80d13dfd",
X"f4055476",
X"5383e7f0",
X"527951ff",
X"a2f23f02",
X"82b90533",
X"55815974",
X"80d72e09",
X"810680c5",
X"38775279",
X"51ffa4b6",
X"3f80d13d",
X"fdf00554",
X"76538f3d",
X"70537a52",
X"58ffa3ee",
X"3f805676",
X"762ea238",
X"751883e7",
X"f0173371",
X"33707232",
X"70307080",
X"2570307f",
X"06811d5d",
X"5f515151",
X"525b55db",
X"3982ac51",
X"e4e13f78",
X"802e8638",
X"80c35184",
X"3980ce51",
X"cadd3fcb",
X"d23fca87",
X"3f83d839",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"05595580",
X"705d5980",
X"e451e4ab",
X"3fcaf43f",
X"80c151ca",
X"ae3f83ea",
X"8808792e",
X"82d63883",
X"eaa80880",
X"fc055580",
X"fd527451",
X"85a03f83",
X"e080085b",
X"778224b2",
X"38ff1870",
X"872b83ff",
X"ff800680",
X"f6f40583",
X"e7f05957",
X"55818055",
X"75708105",
X"57337770",
X"81055934",
X"ff157081",
X"ff065155",
X"74ea3882",
X"85397782",
X"e82e81a3",
X"387782e9",
X"2e098106",
X"81aa3878",
X"58778732",
X"70307072",
X"0780257a",
X"8a327030",
X"70720780",
X"25730753",
X"545a5157",
X"5575802e",
X"97387878",
X"269238a0",
X"0b83e7f0",
X"1a348119",
X"7081ff06",
X"5a55eb39",
X"81187081",
X"ff065955",
X"8a7827ff",
X"bc388f58",
X"83e7eb18",
X"3383e7f0",
X"1934ff18",
X"7081ff06",
X"59557784",
X"26ea3890",
X"58800b83",
X"e7f01934",
X"81187081",
X"ff067098",
X"2b525955",
X"748025e9",
X"3880c655",
X"7a858f24",
X"843880c2",
X"557483e7",
X"f03480f1",
X"0b83e7f3",
X"34810b83",
X"e7f4347a",
X"83e7f134",
X"7a882c55",
X"7483e7f2",
X"3480cb39",
X"82f07825",
X"80c43877",
X"80fd29fd",
X"97d30552",
X"7951ffa1",
X"913f80d1",
X"3dfdec05",
X"5480fd53",
X"83e7f052",
X"7951ffa0",
X"c93f7b81",
X"19595675",
X"80fc2483",
X"38785877",
X"882c5574",
X"83e8ed34",
X"7783e8ee",
X"347583e8",
X"ef348180",
X"5980cc39",
X"83eaa008",
X"57837825",
X"9b3883e9",
X"fc3383e9",
X"fd337188",
X"2b07fc1a",
X"71297905",
X"83800559",
X"51598d39",
X"77818029",
X"17ff8005",
X"57818059",
X"76527951",
X"ffa09f3f",
X"80d13dfd",
X"ec055478",
X"5383e7f0",
X"527951ff",
X"9fd83f78",
X"51f6c33f",
X"c7f53fc6",
X"aa3f8b39",
X"83e9f008",
X"810583e9",
X"f00c80d1",
X"3d0d04f6",
X"e43ffc39",
X"fc3d0d76",
X"78718429",
X"83ea9005",
X"70085153",
X"5353709e",
X"3880ce72",
X"3480cf0b",
X"81133480",
X"ce0b8213",
X"3480c50b",
X"83133470",
X"84133480",
X"e73983ea",
X"a4133354",
X"80d27234",
X"73822a70",
X"81065151",
X"80cf5370",
X"843880d7",
X"53728113",
X"34a00b82",
X"13347383",
X"06517081",
X"2e9e3870",
X"81248838",
X"70802e8f",
X"389f3970",
X"822e9238",
X"70832e92",
X"38933980",
X"d8558e39",
X"80d35589",
X"3980cd55",
X"843980c4",
X"55748313",
X"3480c40b",
X"84133480",
X"0b851334",
X"863d0d04",
X"fc3d0d76",
X"78535481",
X"53805587",
X"39711073",
X"10545273",
X"72265172",
X"802ea738",
X"70802e86",
X"38718025",
X"e8387280",
X"2e983871",
X"74268938",
X"73723175",
X"74075654",
X"72812a72",
X"812a5353",
X"e5397351",
X"78833874",
X"517083e0",
X"800c863d",
X"0d04fe3d",
X"0d805375",
X"527451ff",
X"a33f843d",
X"0d04fe3d",
X"0d815375",
X"527451ff",
X"933f843d",
X"0d04fb3d",
X"0d777955",
X"55805674",
X"76258638",
X"74305581",
X"56738025",
X"88387330",
X"76813257",
X"54805373",
X"527451fe",
X"e73f83e0",
X"80085475",
X"802e8738",
X"83e08008",
X"30547383",
X"e0800c87",
X"3d0d04fa",
X"3d0d787a",
X"57558057",
X"74772586",
X"38743055",
X"8157759f",
X"2c548153",
X"75743274",
X"31527451",
X"feaa3f83",
X"e0800854",
X"76802e87",
X"3883e080",
X"08305473",
X"83e0800c",
X"883d0d04",
X"fd3d0d75",
X"5480740c",
X"800b8415",
X"0c800b88",
X"150c800b",
X"8c150c87",
X"a6803370",
X"81ff0651",
X"51dd933f",
X"70812a81",
X"32718132",
X"71810671",
X"81063184",
X"170c5353",
X"70832a81",
X"3271822a",
X"81327181",
X"06718106",
X"31760c52",
X"5287a090",
X"33700981",
X"0688160c",
X"5183e080",
X"08802e80",
X"c23883e0",
X"8008812a",
X"70810683",
X"e0800881",
X"06318416",
X"0c5183e0",
X"8008832a",
X"83e08008",
X"822a7181",
X"06718106",
X"31760c52",
X"5283e080",
X"08842a81",
X"0688150c",
X"83e08008",
X"852a8106",
X"8c150c85",
X"3d0d04fe",
X"3d0d7476",
X"54527151",
X"fece3f72",
X"812ea238",
X"8173268d",
X"3872822e",
X"a8387283",
X"2e9c38e6",
X"397108e2",
X"38841208",
X"dd388812",
X"08d838a5",
X"39881208",
X"812e9e38",
X"91398812",
X"08812e95",
X"38710891",
X"38841208",
X"8c388c12",
X"08812e09",
X"8106ffb2",
X"38843d0d",
X"04000000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002a93",
X"00002ad4",
X"00002af6",
X"00002b1c",
X"00002b1c",
X"00002b1c",
X"00002b1c",
X"00002b8d",
X"00002bde",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"000039f4",
X"000039f8",
X"00003a00",
X"00003a0c",
X"00003a18",
X"00003a24",
X"00003a30",
X"00003a34",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
