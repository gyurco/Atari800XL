
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81df",
X"f4738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81e9",
X"800c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757581da",
X"a12d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7581d8b5",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80e88604",
X"fd3d0d75",
X"705254ae",
X"c33f83c0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"c0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83c0",
X"8008732e",
X"a13883c0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183c0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83c2d808",
X"248a38b5",
X"983fff0b",
X"83c2d80c",
X"800b83c0",
X"800c04ff",
X"3d0d7352",
X"83c0b408",
X"722e9b38",
X"d93f8183",
X"0b9088a0",
X"0c715196",
X"c93f8193",
X"0b9088a0",
X"0c7183c0",
X"b40c833d",
X"0d04f43d",
X"0d7e6062",
X"5c5a5580",
X"568154bc",
X"1508762e",
X"09810681",
X"92387451",
X"ffb93f79",
X"58757a25",
X"80f73883",
X"c3880870",
X"892a5783",
X"ff067884",
X"80723156",
X"56577378",
X"25833873",
X"557583c2",
X"d8082e84",
X"38fef33f",
X"83c2d808",
X"8025a638",
X"75892b51",
X"98fd3f83",
X"c388088f",
X"3dfc1155",
X"5c548152",
X"f81b5196",
X"e73f7614",
X"83c3880c",
X"7583c2d8",
X"0c745376",
X"527851b3",
X"b33f83c0",
X"800883c3",
X"88081683",
X"c3880c78",
X"7631761b",
X"5b595677",
X"8024ff8b",
X"38617a71",
X"0c547554",
X"75802e83",
X"38815473",
X"83c0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"853f7651",
X"fe993f86",
X"3dfc0553",
X"78527751",
X"968a3f79",
X"75710c54",
X"83c08008",
X"5483c080",
X"08802e83",
X"38815473",
X"83c0800c",
X"863d0d04",
X"fe3d0d75",
X"83c2d808",
X"53538072",
X"24953871",
X"732e9038",
X"80c30b90",
X"88a00c71",
X"9088a40c",
X"fdb43f80",
X"d30b9088",
X"a00c7451",
X"fdc13f80",
X"e30b9088",
X"a00c7251",
X"97b53f80",
X"f30b9088",
X"a00c83c0",
X"80085283",
X"c0800880",
X"2e833881",
X"527183c0",
X"800c843d",
X"0d04803d",
X"0d7280c0",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"3d0d72bc",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"c40b83c0",
X"800c04fd",
X"3d0d7577",
X"71547053",
X"5553a9e4",
X"3f82c813",
X"08bc150c",
X"82c01308",
X"80c0150c",
X"fcb43f73",
X"5193ab3f",
X"7383c0b4",
X"0c83c080",
X"085383c0",
X"8008802e",
X"83388153",
X"7283c080",
X"0c853d0d",
X"04fd3d0d",
X"75775553",
X"fc883f72",
X"802ea538",
X"bc130852",
X"7351a8ee",
X"3f83c080",
X"088f3877",
X"527251ff",
X"9a3f83c0",
X"8008538a",
X"3982cc13",
X"0853d839",
X"81537283",
X"c0800c85",
X"3d0d04fe",
X"3d0dff0b",
X"83c2d80c",
X"7483c0b8",
X"0c7583c2",
X"d40cafc6",
X"3f83c080",
X"0881ff06",
X"52815371",
X"993883c2",
X"f0518e94",
X"3f83c080",
X"085283c0",
X"8008802e",
X"83387252",
X"71537283",
X"c0800c84",
X"3d0d04fa",
X"3d0d787a",
X"82c41208",
X"82c41208",
X"70722459",
X"56565757",
X"73732e09",
X"81069138",
X"80c01652",
X"80c01751",
X"a6df3f83",
X"c0800855",
X"7483c080",
X"0c883d0d",
X"04f63d0d",
X"7c5b807b",
X"715c5457",
X"7a772e8c",
X"38811a82",
X"cc140854",
X"5a72f638",
X"805980d9",
X"397a5481",
X"5780707b",
X"7b315a57",
X"55ff1853",
X"74732580",
X"c13882cc",
X"14085273",
X"51ff8c3f",
X"800b83c0",
X"800825a1",
X"3882cc14",
X"0882cc11",
X"0882cc16",
X"0c7482cc",
X"120c5375",
X"802e8638",
X"7282cc17",
X"0c725480",
X"577382cc",
X"15088117",
X"575556ff",
X"b8398119",
X"59800bff",
X"1b545478",
X"73258338",
X"81547681",
X"32707506",
X"515372ff",
X"90388c3d",
X"0d04f73d",
X"0d7b7d5a",
X"5a82d052",
X"83c2d408",
X"5181c6bb",
X"3f83c080",
X"0857f9aa",
X"3f795283",
X"c2dc5195",
X"b73f83c0",
X"80085480",
X"5383c080",
X"08732e09",
X"81068283",
X"3883c0b8",
X"080b0b81",
X"e5c85370",
X"5256a69c",
X"3f0b0b81",
X"e5c85280",
X"c01651a6",
X"8f3f75bc",
X"170c7382",
X"c0170c81",
X"0b82c417",
X"0c810b82",
X"c8170c73",
X"82cc170c",
X"ff1782d0",
X"17555781",
X"913983c0",
X"c4337082",
X"2a708106",
X"51545572",
X"81803874",
X"812a8106",
X"587780f6",
X"3874842a",
X"810682c4",
X"150c83c0",
X"c4338106",
X"82c8150c",
X"79527351",
X"a5b63f73",
X"51a5cd3f",
X"83c08008",
X"1453af73",
X"70810555",
X"3472bc15",
X"0c83c0c5",
X"527251a5",
X"973f83c0",
X"bc0882c0",
X"150c83c0",
X"d25280c0",
X"1451a584",
X"3f78802e",
X"8d387351",
X"782d83c0",
X"8008802e",
X"99387782",
X"cc150c75",
X"802e8638",
X"7382cc17",
X"0c7382d0",
X"15ff1959",
X"55567680",
X"2e9b3883",
X"c0bc5283",
X"c2dc5194",
X"ad3f83c0",
X"80088a38",
X"83c0c533",
X"5372fed2",
X"3878802e",
X"893883c0",
X"b80851fc",
X"b83f83c0",
X"b8085372",
X"83c0800c",
X"8b3d0d04",
X"ff3d0d80",
X"527351fd",
X"b53f833d",
X"0d04f03d",
X"0d627052",
X"54f5d93f",
X"83c08008",
X"7453873d",
X"70535555",
X"f5f93ff6",
X"d93f7351",
X"d33f6353",
X"745283c0",
X"800851fa",
X"b83f923d",
X"0d047183",
X"c0800c04",
X"80c01283",
X"c0800c04",
X"803d0d72",
X"82c01108",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"7282cc11",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d7282c4",
X"110883c0",
X"800c5182",
X"3d0d04f9",
X"3d0d7983",
X"c0900857",
X"57817727",
X"81963876",
X"88170827",
X"818e3875",
X"33557482",
X"2e893874",
X"832eb338",
X"80fe3974",
X"54761083",
X"fe065376",
X"882a8c17",
X"08055289",
X"3dfc0551",
X"a9f43f83",
X"c0800880",
X"df38029d",
X"0533893d",
X"3371882b",
X"07565680",
X"d1398454",
X"76822b83",
X"fc065376",
X"872a8c17",
X"08055289",
X"3dfc0551",
X"a9c43f83",
X"c08008b0",
X"38029f05",
X"33028405",
X"9e053371",
X"982b7190",
X"2b07028c",
X"059d0533",
X"70882b72",
X"078d3d33",
X"7180ffff",
X"fe800607",
X"51525357",
X"58568339",
X"81557483",
X"c0800c89",
X"3d0d04fb",
X"3d0d83c0",
X"9008fe19",
X"881208fe",
X"05555654",
X"80567473",
X"278d3882",
X"14337571",
X"29941608",
X"05575375",
X"83c0800c",
X"873d0d04",
X"fc3d0d76",
X"52800b83",
X"c0900870",
X"33515253",
X"70832e09",
X"81069138",
X"95123394",
X"13337198",
X"2b71902b",
X"07555551",
X"9b12339a",
X"13337188",
X"2b077407",
X"83c0800c",
X"55863d0d",
X"04fc3d0d",
X"7683c090",
X"08555580",
X"75238815",
X"08537281",
X"2e883888",
X"14087326",
X"85388152",
X"b2397290",
X"38733352",
X"71832e09",
X"81068538",
X"90140853",
X"728c160c",
X"72802e8d",
X"387251fe",
X"d63f83c0",
X"80085285",
X"39901408",
X"52719016",
X"0c805271",
X"83c0800c",
X"863d0d04",
X"fa3d0d78",
X"83c09008",
X"71228105",
X"7083ffff",
X"06575457",
X"5573802e",
X"88389015",
X"08537286",
X"38835280",
X"e739738f",
X"06527180",
X"da388113",
X"90160c8c",
X"15085372",
X"9038830b",
X"84172257",
X"52737627",
X"80c638bf",
X"39821633",
X"ff057484",
X"2a065271",
X"b2387251",
X"fcb13f81",
X"527183c0",
X"800827a8",
X"38835283",
X"c0800888",
X"1708279c",
X"3883c080",
X"088c160c",
X"83c08008",
X"51fdbc3f",
X"83c08008",
X"90160c73",
X"75238052",
X"7183c080",
X"0c883d0d",
X"04f23d0d",
X"60626458",
X"5e5b7533",
X"5574a02e",
X"09810688",
X"38811670",
X"4456ef39",
X"62703356",
X"5674af2e",
X"09810684",
X"38811643",
X"800b881c",
X"0c627033",
X"5155749f",
X"2691387a",
X"51fdd23f",
X"83c08008",
X"56807d34",
X"83813993",
X"3d841c08",
X"7058595f",
X"8a55a076",
X"70810558",
X"34ff1555",
X"74ff2e09",
X"8106ef38",
X"80705a5c",
X"887f085f",
X"5a7b811d",
X"7081ff06",
X"60137033",
X"70af3270",
X"30a07327",
X"71802507",
X"5151525b",
X"535e5755",
X"7480e738",
X"76ae2e09",
X"81068338",
X"8155787a",
X"27750755",
X"74802e9f",
X"38798832",
X"703078ae",
X"32703070",
X"73079f2a",
X"53515751",
X"5675bb38",
X"88598b5a",
X"ffab3976",
X"982b5574",
X"80258738",
X"81df8417",
X"3357ff9f",
X"17557499",
X"268938e0",
X"177081ff",
X"06585578",
X"811a7081",
X"ff06721b",
X"535b5755",
X"767534fe",
X"f8397b1e",
X"7f0c8055",
X"76a02683",
X"38815574",
X"8b19347a",
X"51fc823f",
X"83c08008",
X"80f538a0",
X"547a2270",
X"852b83e0",
X"06545590",
X"1b08527c",
X"51a3ff3f",
X"83c08008",
X"5783c080",
X"08818138",
X"7c335574",
X"802e80f4",
X"388b1d33",
X"70832a70",
X"81065156",
X"5674b438",
X"8b7d841d",
X"0883c080",
X"08595b5b",
X"58ff1858",
X"77ff2e9a",
X"38797081",
X"055b3379",
X"7081055b",
X"33717131",
X"52565675",
X"802ee238",
X"86397580",
X"2e96387a",
X"51fbe53f",
X"ff863983",
X"c0800856",
X"83c08008",
X"b6388339",
X"7656841b",
X"088b1133",
X"515574a7",
X"388b1d33",
X"70842a70",
X"81065156",
X"56748938",
X"83569439",
X"81569039",
X"7c51fa94",
X"3f83c080",
X"08881c0c",
X"fd813975",
X"83c0800c",
X"903d0d04",
X"f83d0d7a",
X"7c595782",
X"5483fe53",
X"77527651",
X"a2c43f83",
X"5683c080",
X"0880ec38",
X"81173377",
X"3371882b",
X"07565682",
X"567482d4",
X"d52e0981",
X"0680d438",
X"7554b653",
X"77527651",
X"a2983f83",
X"c0800898",
X"38811733",
X"77337188",
X"2b0783c0",
X"80085256",
X"56748182",
X"c62eac38",
X"825480d2",
X"53775276",
X"51a1ef3f",
X"83c08008",
X"98388117",
X"33773371",
X"882b0783",
X"c0800852",
X"56567481",
X"82c62e83",
X"38815675",
X"83c0800c",
X"8a3d0d04",
X"eb3d0d67",
X"5a800b83",
X"c0900ca1",
X"913f83c0",
X"80088106",
X"55825674",
X"83ef3874",
X"75538f3d",
X"70535759",
X"feca3f83",
X"c0800881",
X"ff065776",
X"812e0981",
X"0680d438",
X"905483be",
X"53745275",
X"51a1833f",
X"83c08008",
X"80c9388f",
X"3d335574",
X"802e80c9",
X"3802bf05",
X"33028405",
X"be053371",
X"982b7190",
X"2b07028c",
X"05bd0533",
X"70882b72",
X"07953d33",
X"71077058",
X"7b575e52",
X"5e575957",
X"fdee3f83",
X"c0800881",
X"ff065776",
X"832e0981",
X"06863881",
X"5682f239",
X"76802e86",
X"38865682",
X"e839a454",
X"8d537852",
X"7551a09a",
X"3f815683",
X"c0800882",
X"d43802be",
X"05330284",
X"05bd0533",
X"71882b07",
X"595d77ab",
X"380280ce",
X"05330284",
X"0580cd05",
X"3371982b",
X"71902b07",
X"973d3370",
X"882b7207",
X"02940580",
X"cb053371",
X"0754525e",
X"57595602",
X"b7053378",
X"71290288",
X"05b60533",
X"028c05b5",
X"05337188",
X"2b07701d",
X"707f8c05",
X"0c5f5957",
X"595d8e3d",
X"33821b34",
X"02b90533",
X"903d3371",
X"882b075a",
X"5c78841b",
X"2302bb05",
X"33028405",
X"ba053371",
X"882b0756",
X"5c74ab38",
X"0280ca05",
X"33028405",
X"80c90533",
X"71982b71",
X"902b0796",
X"3d337088",
X"2b720702",
X"940580c7",
X"05337107",
X"51525357",
X"5e5c7476",
X"31783179",
X"842a903d",
X"33547171",
X"31535656",
X"81b7a03f",
X"83c08008",
X"82057088",
X"1c0c83c0",
X"8008e08a",
X"05565674",
X"83dffe26",
X"83388257",
X"83fff676",
X"27853883",
X"57893986",
X"5676802e",
X"80db3876",
X"7a347683",
X"2e098106",
X"b0380280",
X"d6053302",
X"840580d5",
X"05337198",
X"2b71902b",
X"07993d33",
X"70882b72",
X"07029405",
X"80d30533",
X"71077f90",
X"050c525e",
X"57585686",
X"39771b90",
X"1b0c841a",
X"228c1b08",
X"1971842a",
X"05941c0c",
X"5d800b81",
X"1b347983",
X"c0900c80",
X"567583c0",
X"800c973d",
X"0d04e93d",
X"0d83c090",
X"08568554",
X"75802e81",
X"8238800b",
X"81173499",
X"3de01146",
X"6a548a3d",
X"705458ec",
X"0551f6e5",
X"3f83c080",
X"085483c0",
X"800880df",
X"38893d33",
X"5473802e",
X"913802ab",
X"05337084",
X"2a810651",
X"5574802e",
X"86388354",
X"80c13976",
X"51f4893f",
X"83c08008",
X"a0170c02",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"9c1c0c52",
X"78981b0c",
X"53565957",
X"810b8117",
X"34745473",
X"83c0800c",
X"993d0d04",
X"f53d0d7d",
X"7f617283",
X"c090085a",
X"5d5d595c",
X"807b0c85",
X"5775802e",
X"81e03881",
X"16338106",
X"55845774",
X"802e81d2",
X"38913974",
X"81173486",
X"39800b81",
X"17348157",
X"81c0399c",
X"16089817",
X"08315574",
X"78278338",
X"74587780",
X"2e81a938",
X"98160870",
X"83ff0656",
X"577480cf",
X"38821633",
X"ff057789",
X"2a067081",
X"ff065a55",
X"78a03876",
X"8738a016",
X"08558d39",
X"a4160851",
X"f0e93f83",
X"c0800855",
X"817527ff",
X"a83874a4",
X"170ca416",
X"0851f283",
X"3f83c080",
X"085583c0",
X"8008802e",
X"ff893883",
X"c0800819",
X"a8170c98",
X"160883ff",
X"06848071",
X"31515577",
X"75278338",
X"77557483",
X"ffff0654",
X"98160883",
X"ff0653a8",
X"16085279",
X"577b8338",
X"7b577651",
X"9ac03f83",
X"c08008fe",
X"d0389816",
X"08159817",
X"0c741a78",
X"76317c08",
X"177d0c59",
X"5afed339",
X"80577683",
X"c0800c8d",
X"3d0d04fa",
X"3d0d7883",
X"c0900855",
X"56855573",
X"802e81e3",
X"38811433",
X"81065384",
X"5572802e",
X"81d5389c",
X"14085372",
X"76278338",
X"72569814",
X"0857800b",
X"98150c75",
X"802e81b9",
X"38821433",
X"70892b56",
X"5376802e",
X"b7387452",
X"ff165181",
X"b2a13f83",
X"c08008ff",
X"18765470",
X"53585381",
X"b2913f83",
X"c0800873",
X"26963874",
X"30707806",
X"7098170c",
X"777131a4",
X"17085258",
X"51538939",
X"a0140870",
X"a4160c53",
X"747627b9",
X"387251ee",
X"d63f83c0",
X"80085381",
X"0b83c080",
X"08278b38",
X"88140883",
X"c0800826",
X"8838800b",
X"811534b0",
X"3983c080",
X"08a4150c",
X"98140815",
X"98150c75",
X"753156c4",
X"39981408",
X"16709816",
X"0c735256",
X"efc53f83",
X"c080088c",
X"3883c080",
X"08811534",
X"81559439",
X"821433ff",
X"0576892a",
X"0683c080",
X"0805a815",
X"0c805574",
X"83c0800c",
X"883d0d04",
X"ef3d0d63",
X"56855583",
X"c0900880",
X"2e80d238",
X"933df405",
X"84170c64",
X"53883d70",
X"53765257",
X"f1cf3f83",
X"c0800855",
X"83c08008",
X"b438883d",
X"33547380",
X"2ea13802",
X"a7053370",
X"842a7081",
X"06515555",
X"83557380",
X"2e973876",
X"51eef53f",
X"83c08008",
X"88170c75",
X"51efa63f",
X"83c08008",
X"557483c0",
X"800c933d",
X"0d04e43d",
X"0d6ea13d",
X"08405e85",
X"5683c090",
X"08802e84",
X"85389e3d",
X"f405841f",
X"0c7e9838",
X"7d51eef5",
X"3f83c080",
X"085683ee",
X"39814181",
X"f6398341",
X"81f13993",
X"3d7f9605",
X"4159807f",
X"8295055e",
X"56756081",
X"ff053483",
X"41901e08",
X"762e81d3",
X"38a0547d",
X"2270852b",
X"83e00654",
X"58901e08",
X"52785196",
X"c93f83c0",
X"80084183",
X"c08008ff",
X"b8387833",
X"5c7b802e",
X"ffb4388b",
X"193370bf",
X"06718106",
X"52435574",
X"802e80de",
X"387b81bf",
X"0655748f",
X"2480d338",
X"9a193355",
X"7480cb38",
X"f31d7058",
X"5d815675",
X"8b2e0981",
X"0685388e",
X"568b3975",
X"9a2e0981",
X"0683389c",
X"56751970",
X"70810552",
X"33713381",
X"1a821a5f",
X"5b525b55",
X"74863879",
X"77348539",
X"80df7734",
X"777b5757",
X"7aa02e09",
X"8106c038",
X"81567b81",
X"e5327030",
X"709f2a51",
X"51557bae",
X"2e933874",
X"802e8e38",
X"61832a70",
X"81065155",
X"74802e97",
X"387d51ed",
X"df3f83c0",
X"80084183",
X"c0800887",
X"38901e08",
X"feaf3880",
X"60347580",
X"2e88387c",
X"527f518d",
X"eb3f6080",
X"2e863880",
X"0b901f0c",
X"60566083",
X"2e853860",
X"81d03889",
X"1f57901e",
X"08802e81",
X"a8388056",
X"75197033",
X"515574a0",
X"2ea03874",
X"852e0981",
X"06843881",
X"e5557477",
X"70810559",
X"34811670",
X"81ff0657",
X"55877627",
X"d7388819",
X"335574a0",
X"2ea938ae",
X"77708105",
X"59348856",
X"75197033",
X"515574a0",
X"2e953874",
X"77708105",
X"59348116",
X"7081ff06",
X"57558a76",
X"27e2388b",
X"19337f88",
X"05349f19",
X"339e1a33",
X"71982b71",
X"902b079d",
X"1c337088",
X"2b72079c",
X"1e337107",
X"640c5299",
X"1d33981e",
X"3371882b",
X"07535153",
X"57595674",
X"7f840523",
X"97193396",
X"1a337188",
X"2b075656",
X"747f8605",
X"23807734",
X"7d51ebf0",
X"3f83c080",
X"08833270",
X"30707207",
X"9f2c83c0",
X"80080652",
X"5656961f",
X"3355748a",
X"38891f52",
X"961f518b",
X"f73f7583",
X"c0800c9e",
X"3d0d04f4",
X"3d0d7e8f",
X"3dec1156",
X"56589053",
X"f0155277",
X"51e0b13f",
X"83c08008",
X"80d63878",
X"902e0981",
X"0680cd38",
X"02ab0533",
X"81e9880b",
X"81e98833",
X"5758568c",
X"3974762e",
X"8a388417",
X"70335657",
X"74f33876",
X"33705755",
X"74802eac",
X"38821722",
X"708a2b90",
X"3dec0556",
X"70555656",
X"96800a52",
X"7751dfe0",
X"3f83c080",
X"08863878",
X"752e8538",
X"80568539",
X"81173356",
X"7583c080",
X"0c8e3d0d",
X"04fc3d0d",
X"76705255",
X"8afe3f83",
X"c0800815",
X"ff055473",
X"752e8e38",
X"73335372",
X"ae2e8638",
X"ff1454ef",
X"39775281",
X"14518a96",
X"3f83c080",
X"08307083",
X"c0800807",
X"802583c0",
X"800c5386",
X"3d0d04fa",
X"3d0d7857",
X"80775256",
X"e6c23f83",
X"c0800883",
X"c0800833",
X"53547176",
X"2e80c738",
X"733383c0",
X"94173356",
X"53749138",
X"765183c3",
X"ac085271",
X"2d83c080",
X"0852ad39",
X"ff9f1352",
X"71992689",
X"38e01370",
X"81ff0654",
X"52747332",
X"70307072",
X"07802578",
X"05811770",
X"33545758",
X"545271ff",
X"bb388052",
X"7183c080",
X"0c883d0d",
X"04fc3d0d",
X"76705255",
X"e6803f83",
X"c0800854",
X"815383c0",
X"800880d0",
X"387451e5",
X"c33f83c0",
X"800881e5",
X"d85383c0",
X"80085253",
X"fea33f83",
X"c08008b0",
X"3881e5dc",
X"527251fe",
X"943f83c0",
X"8008a138",
X"81e5e052",
X"7251fe85",
X"3f83c080",
X"08923881",
X"e5e45272",
X"51fdf63f",
X"83c08008",
X"802e8338",
X"81547353",
X"7283c080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"e5903f81",
X"5383c080",
X"08983873",
X"51e4d93f",
X"83c3a008",
X"5283c080",
X"0851fdbd",
X"3f83c080",
X"08537283",
X"c0800c85",
X"3d0d04dd",
X"3d0da63d",
X"085f800b",
X"83c7e033",
X"555b737b",
X"2e85cc38",
X"86537a52",
X"83c09451",
X"a1c73f7e",
X"51daae3f",
X"83c08008",
X"33973d56",
X"54737b2e",
X"09810696",
X"3881eac8",
X"52745187",
X"db3f9a39",
X"7e527851",
X"dde13f85",
X"96397e51",
X"da8f3f83",
X"c0800852",
X"7451d9bf",
X"3f804480",
X"43804280",
X"41adbb52",
X"963d7052",
X"5ee0cb3f",
X"83c08008",
X"59800b83",
X"c0800855",
X"5c83c080",
X"087c2e94",
X"38811c74",
X"525ce3cd",
X"3f83c080",
X"085483c0",
X"8008ee38",
X"805aff40",
X"7909709f",
X"2c7b065b",
X"547b7a24",
X"8438ff1c",
X"5af61a70",
X"09709f2c",
X"72067bff",
X"125a5a52",
X"55558075",
X"25953876",
X"51e3923f",
X"83c08008",
X"76ff1858",
X"55577380",
X"24ed3874",
X"602e8638",
X"a2823f74",
X"4078ff1b",
X"70585e58",
X"807a2595",
X"387751e2",
X"e83f83c0",
X"800876ff",
X"18585558",
X"738024ed",
X"38800b83",
X"c7dc0c81",
X"800b83c8",
X"980c81e5",
X"e8518bdf",
X"3f800b83",
X"c8980c83",
X"c0945281",
X"e5f0518b",
X"ce3fa80b",
X"83c7dc0c",
X"76802e80",
X"e43883c7",
X"dc087779",
X"32703070",
X"72078025",
X"70872b83",
X"c8980c51",
X"56785356",
X"56e29b3f",
X"83c08008",
X"802e8838",
X"81e5fc51",
X"8b953f76",
X"51e1dd3f",
X"83c08008",
X"5281e8a8",
X"518b843f",
X"7651e1e5",
X"3f83c080",
X"0883c7dc",
X"08555775",
X"74258638",
X"a81656f7",
X"397583c7",
X"dc0c86f0",
X"7624ff98",
X"3887980b",
X"83c7dc0c",
X"77802ea9",
X"387751e1",
X"9b3f83c0",
X"80087852",
X"55e1bb3f",
X"81e68454",
X"83c08008",
X"853881e6",
X"80547453",
X"735281e5",
X"cc518aab",
X"3f805481",
X"e5d4518a",
X"a23f8114",
X"5473a82e",
X"098106ef",
X"38868da0",
X"519e803f",
X"8052913d",
X"705257ba",
X"933f8352",
X"7651ba8c",
X"3f645473",
X"ff2e0981",
X"069738ff",
X"1b700970",
X"9f2c7206",
X"52555b80",
X"0b83c094",
X"1c3481c2",
X"39807425",
X"ab387a85",
X"2e098106",
X"91388653",
X"805283c0",
X"94519dbd",
X"3f805b81",
X"a5397383",
X"c0941c34",
X"811b5b81",
X"99398076",
X"34819339",
X"63818f38",
X"62802e80",
X"fb387c54",
X"73ff2e96",
X"3878802e",
X"81893878",
X"51dffa3f",
X"83c08008",
X"ff155559",
X"e7397880",
X"2e80f438",
X"7851dff6",
X"3f83c080",
X"08802efb",
X"c7387851",
X"dfbe3f83",
X"c0800852",
X"81e5c851",
X"81e73f83",
X"c08008a3",
X"387d5183",
X"9f3f83c0",
X"80085574",
X"ff165654",
X"807425ae",
X"38741e70",
X"33555673",
X"af2eff8a",
X"38e93978",
X"51deff3f",
X"83c08008",
X"527d5182",
X"d73f8f39",
X"60882961",
X"10057a05",
X"62055afb",
X"c7396380",
X"2efb8a38",
X"80527651",
X"b89e3fa5",
X"3d0d04ff",
X"3d0d028f",
X"05337010",
X"81059088",
X"900c5283",
X"3d0d04ff",
X"3d0d028f",
X"05335290",
X"88840870",
X"892a7081",
X"06515151",
X"70802e86",
X"38afca3f",
X"ea397190",
X"88800c83",
X"3d0d0480",
X"3d0d9088",
X"8c087088",
X"2a708106",
X"51515170",
X"802e8638",
X"afa73fea",
X"39908888",
X"0883c080",
X"0c823d0d",
X"04908894",
X"0883c080",
X"0c04fd3d",
X"0d757754",
X"54807325",
X"94387370",
X"81055533",
X"5281e688",
X"5187883f",
X"ff1353e9",
X"39853d0d",
X"04fd3d0d",
X"75775354",
X"73335170",
X"89387133",
X"5170802e",
X"a1387333",
X"72335253",
X"72712785",
X"38ff5194",
X"39707327",
X"85388151",
X"8b398114",
X"81135354",
X"d3398051",
X"7083c080",
X"0c853d0d",
X"04fd3d0d",
X"75775454",
X"72337081",
X"ff065252",
X"70802ea3",
X"387181ff",
X"068114ff",
X"bf125354",
X"52709926",
X"8938a012",
X"7081ff06",
X"53517174",
X"70810556",
X"34d23980",
X"7434853d",
X"0d04ffbd",
X"3d0d80c6",
X"3d0852a5",
X"3d705254",
X"ffb33f80",
X"c73d0852",
X"853d7052",
X"53ffa63f",
X"72527351",
X"fedf3f80",
X"c53d0d04",
X"fe3d0d74",
X"76535371",
X"70810553",
X"33517073",
X"70810555",
X"3470f038",
X"843d0d04",
X"fe3d0d74",
X"52807233",
X"52537073",
X"2e8d3881",
X"12811471",
X"33535452",
X"70f53872",
X"83c0800c",
X"843d0d04",
X"f63d0d7c",
X"7e60625a",
X"5d5b5680",
X"59815585",
X"39747a29",
X"55745275",
X"51819f8f",
X"3f83c080",
X"087a27ed",
X"3874802e",
X"80e03874",
X"52755181",
X"9ef93f83",
X"c0800875",
X"53765254",
X"819f9f3f",
X"83c08008",
X"7a537552",
X"56819edf",
X"3f83c080",
X"08793070",
X"7b079f2a",
X"70778024",
X"07515154",
X"55728738",
X"83c08008",
X"c2387681",
X"18b01655",
X"58588974",
X"258b38b7",
X"14537a85",
X"3880d714",
X"53727834",
X"811959ff",
X"9c398077",
X"348c3d0d",
X"04f73d0d",
X"7b7d7f62",
X"029005bb",
X"05335759",
X"565a5ab0",
X"58728338",
X"a0587570",
X"70810552",
X"33715954",
X"55903980",
X"74258e38",
X"ff147770",
X"81055933",
X"545472ef",
X"3873ff15",
X"55538073",
X"25893877",
X"52795178",
X"2def3975",
X"33755753",
X"72802e90",
X"38725279",
X"51782d75",
X"70810557",
X"3353ed39",
X"8b3d0d04",
X"ee3d0d64",
X"66696970",
X"70810552",
X"335b4a5c",
X"5e5e7680",
X"2e82f938",
X"76a52e09",
X"810682e0",
X"38807041",
X"67707081",
X"05523371",
X"4a59575f",
X"76b02e09",
X"81068c38",
X"75708105",
X"57337648",
X"57815fd0",
X"17567589",
X"2680da38",
X"76675c59",
X"805c9339",
X"778a2480",
X"c3387b8a",
X"29187b70",
X"81055d33",
X"5a5cd019",
X"7081ff06",
X"58588977",
X"27a438ff",
X"9f197081",
X"ff06ffa9",
X"1b5a5156",
X"85762792",
X"38ffbf19",
X"7081ff06",
X"51567585",
X"268a38c9",
X"19587780",
X"25ffb938",
X"7a477b40",
X"7881ff06",
X"577680e4",
X"2e80e538",
X"7680e424",
X"a7387680",
X"d82e8186",
X"387680d8",
X"24903876",
X"802e81cc",
X"3876a52e",
X"81b63881",
X"b9397680",
X"e32e818c",
X"3881af39",
X"7680f52e",
X"9b387680",
X"f5248b38",
X"7680f32e",
X"81813881",
X"99397680",
X"f82e80ca",
X"38818f39",
X"913d7055",
X"5780538a",
X"5279841b",
X"7108535b",
X"56fbfd3f",
X"7655ab39",
X"79841b71",
X"08943d70",
X"5b5b525b",
X"56758025",
X"8c387530",
X"56ad7834",
X"0280c105",
X"57765480",
X"538a5275",
X"51fbd13f",
X"77557e54",
X"b839913d",
X"70557780",
X"d8327030",
X"70802556",
X"51585690",
X"5279841b",
X"7108535b",
X"57fbad3f",
X"7555db39",
X"79841b83",
X"1233545b",
X"56983979",
X"841b7108",
X"575b5680",
X"547f537c",
X"527d51fc",
X"9c3f8739",
X"76527d51",
X"7c2d6670",
X"33588105",
X"47fd8339",
X"943d0d04",
X"7283c09c",
X"0c7183c0",
X"a00c04fb",
X"3d0d883d",
X"70708405",
X"52085754",
X"755383c0",
X"9c085283",
X"c0a00851",
X"fcc63f87",
X"3d0d04ff",
X"3d0d7370",
X"08535102",
X"93053372",
X"34700881",
X"05710c83",
X"3d0d04fc",
X"3d0d873d",
X"88115578",
X"54bddb53",
X"51fc993f",
X"8052873d",
X"51d13f86",
X"3d0d04fc",
X"3d0d7655",
X"7483c3b8",
X"082eaf38",
X"80537451",
X"87cc3f83",
X"c0800881",
X"ff06ff14",
X"7081ff06",
X"7230709f",
X"2a515255",
X"53547280",
X"2e843871",
X"dd3873fe",
X"387483c3",
X"b80c863d",
X"0d04ff3d",
X"0dff0b83",
X"c3b80c84",
X"b43f8151",
X"87903f83",
X"c0800881",
X"ff065271",
X"ee3881d4",
X"3f7183c0",
X"800c833d",
X"0d04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"823f7280",
X"2ea03883",
X"c3cc1433",
X"75708105",
X"57348114",
X"7083ffff",
X"06ff1570",
X"83ffff06",
X"56525552",
X"dd39800b",
X"83c0800c",
X"863d0d04",
X"fc3d0d76",
X"787a1156",
X"53558053",
X"71742e93",
X"38721551",
X"703383c3",
X"cc133481",
X"12811454",
X"52ea3980",
X"0b83c080",
X"0c863d0d",
X"04fd3d0d",
X"905483c3",
X"b8085186",
X"fd3f83c0",
X"800881ff",
X"06ff1571",
X"30713070",
X"73079f2a",
X"729f2a06",
X"52555255",
X"5372db38",
X"853d0d04",
X"803d0d83",
X"c3c40883",
X"2b83c3c0",
X"08079080",
X"a80c823d",
X"0d04800b",
X"83c3c40c",
X"e33f0481",
X"0b83c3c4",
X"0cda3f04",
X"ed3f0471",
X"83c3bc0c",
X"04803d0d",
X"8051f43f",
X"810b83c3",
X"c40c860b",
X"83c3c00c",
X"ffba3f82",
X"3d0d0484",
X"0b83c3c0",
X"0cffad3f",
X"04860b83",
X"c3c00cff",
X"a33f0483",
X"0b83c3c0",
X"0cff993f",
X"04870b83",
X"c3c00cff",
X"8f3f0480",
X"3d0d028b",
X"05339080",
X"a40c9080",
X"a8087081",
X"06515170",
X"f5389080",
X"a4087081",
X"ff0683c0",
X"800c5182",
X"3d0d0480",
X"3d0d81ff",
X"51d13f83",
X"c0800881",
X"ff0683c0",
X"800c823d",
X"0d04803d",
X"0d73902b",
X"73079080",
X"b40c823d",
X"0d0404fb",
X"3d0d7802",
X"84059f05",
X"3370982b",
X"55575572",
X"80259b38",
X"7580ff06",
X"56805280",
X"f751e03f",
X"83c08008",
X"81ff0654",
X"73812680",
X"fb38fee1",
X"3fffa43f",
X"fed13fff",
X"9e3f7551",
X"fef13f74",
X"982a51fe",
X"ea3f7490",
X"2a7081ff",
X"065253fe",
X"de3f7488",
X"2a7081ff",
X"065253fe",
X"d23f7481",
X"ff0651fe",
X"ca3f8155",
X"7580c02e",
X"09810686",
X"38819555",
X"8d397580",
X"c82e0981",
X"06843881",
X"87557451",
X"fea93f8a",
X"55fecc3f",
X"83c08008",
X"81ff0670",
X"982b5454",
X"7280258c",
X"38ff1570",
X"81ff0656",
X"5374e238",
X"7383c080",
X"0c873d0d",
X"04fa3d0d",
X"fdb73ffd",
X"d83f8a54",
X"fe993fff",
X"147081ff",
X"06555373",
X"f3387374",
X"535580c0",
X"51feac3f",
X"83c08008",
X"81ff0654",
X"73812e09",
X"8106829f",
X"3883aa52",
X"80c851fe",
X"923f83c0",
X"800881ff",
X"06537281",
X"2e098106",
X"81a83874",
X"54873d74",
X"115456fd",
X"ce3f83c0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e5",
X"38029a05",
X"33537281",
X"2e098106",
X"81d93802",
X"9b053353",
X"80ce9054",
X"7281aa2e",
X"8d3881c7",
X"3980e451",
X"8d8d3fff",
X"14547380",
X"2e81b838",
X"820a5281",
X"e951fdab",
X"3f83c080",
X"0881ff06",
X"5372de38",
X"725280fa",
X"51fd983f",
X"83c08008",
X"81ff0653",
X"72819038",
X"72547316",
X"53fcdc3f",
X"83c08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e83887",
X"3d337086",
X"2a708106",
X"5154548c",
X"557280e3",
X"38845580",
X"de397452",
X"81e951fc",
X"d23f83c0",
X"800881ff",
X"06538255",
X"81e95681",
X"73278638",
X"735580c1",
X"5680ce90",
X"548a3980",
X"e4518bff",
X"3fff1454",
X"73802ea9",
X"38805275",
X"51fca03f",
X"83c08008",
X"81ff0653",
X"72e13884",
X"805280d0",
X"51fc8c3f",
X"83c08008",
X"81ff0653",
X"72802e83",
X"38805574",
X"83c3c834",
X"fb873ffb",
X"ca3f883d",
X"0d04fb3d",
X"0d775480",
X"0b83c3c8",
X"3370832a",
X"70810651",
X"55575572",
X"752e0981",
X"06853873",
X"892b5473",
X"5280d151",
X"fbc53f83",
X"c0800881",
X"ff065372",
X"bd3882b8",
X"c054fb8b",
X"3f83c080",
X"0881ff06",
X"537281ff",
X"2e098106",
X"8938ff14",
X"5473e738",
X"9f397281",
X"fe2e0981",
X"06963883",
X"c7cc5283",
X"c3cc51fa",
X"f53ffadb",
X"3ffad83f",
X"83398155",
X"fa8b3ffa",
X"ce3f7481",
X"ff0683c0",
X"800c873d",
X"0d04fb3d",
X"0d7783c3",
X"cc5654f9",
X"e63f83c3",
X"c8337083",
X"2a708106",
X"51545672",
X"85387389",
X"2b547352",
X"80d851fa",
X"c23f83c0",
X"800881ff",
X"06537280",
X"e73881ff",
X"51f9e03f",
X"81fe51f9",
X"da3f8480",
X"53747081",
X"05563351",
X"f9cd3fff",
X"137083ff",
X"ff065153",
X"72eb3872",
X"51f9bc3f",
X"7251f9b7",
X"3ff9dc3f",
X"83c08008",
X"9f0653a7",
X"88547285",
X"2e8c389e",
X"3980e451",
X"89bd3fff",
X"1454f9bf",
X"3f83c080",
X"0881ff06",
X"537281ff",
X"2e843873",
X"e438f8e5",
X"3ff9a83f",
X"800b83c0",
X"800c873d",
X"0d047183",
X"c7d00c88",
X"80800b83",
X"c7cc0c84",
X"80800b83",
X"c7d40c04",
X"f03d0d83",
X"80805683",
X"c7d00816",
X"83c7cc08",
X"17565474",
X"33743483",
X"c7d40816",
X"54807434",
X"81165675",
X"8380a02e",
X"098106db",
X"3883d080",
X"5683c7d0",
X"081683c7",
X"cc081756",
X"54743374",
X"3483c7d4",
X"08165480",
X"74348116",
X"567583d0",
X"902e0981",
X"06db3883",
X"a8805683",
X"c7d00816",
X"83c7cc08",
X"17565474",
X"33743483",
X"c7d40816",
X"54807434",
X"81165675",
X"83a8902e",
X"098106db",
X"38805683",
X"c7d00816",
X"83c7d408",
X"17555573",
X"33753481",
X"16567581",
X"80802e09",
X"8106e438",
X"89da3f89",
X"3d58a253",
X"81e18452",
X"77518194",
X"f93f8057",
X"8c805683",
X"c7d40816",
X"77195555",
X"73337534",
X"81168118",
X"585676a2",
X"2e098106",
X"e638860b",
X"87a88334",
X"800b87a8",
X"8234800b",
X"87809a34",
X"af0b8780",
X"9634bf0b",
X"87809734",
X"800b8780",
X"98349f0b",
X"87809934",
X"800b8780",
X"9b34f80b",
X"87a88934",
X"7687a880",
X"34820b87",
X"d08f3482",
X"0b87a881",
X"34840b87",
X"809f34ff",
X"0b87d08b",
X"34923d0d",
X"04fe3d0d",
X"805383c7",
X"d4081383",
X"c7d00814",
X"52527033",
X"72348113",
X"53728180",
X"802e0981",
X"06e43883",
X"80805383",
X"c7d40813",
X"83c7d008",
X"14525270",
X"33723481",
X"13537283",
X"80a02e09",
X"8106e438",
X"83d08053",
X"83c7d408",
X"1383c7d0",
X"08145252",
X"70337234",
X"81135372",
X"83d0902e",
X"098106e4",
X"3883a880",
X"5383c7d4",
X"081383c7",
X"d0081452",
X"52703372",
X"34811353",
X"7283a890",
X"2e098106",
X"e438843d",
X"0d04803d",
X"0d908090",
X"08810683",
X"c0800c82",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe067607",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"812c8106",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fd06",
X"76100772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087082",
X"2cbf0683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fe8306",
X"76822b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"882c8706",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f1ff",
X"0676882b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"708b2c81",
X"0683c080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870ef",
X"ff06768b",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870912c",
X"bf0683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fc87ffff",
X"0676912b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70992c81",
X"0683c080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870ff",
X"bf0a0676",
X"992b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"9008709a",
X"2c830683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70cf0a06",
X"769a2b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"9c2c8706",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f10a",
X"06769c2b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"9080bc08",
X"870683c0",
X"800c823d",
X"0d04ff3d",
X"0d9080bc",
X"700870f8",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"bc087084",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80bc7008",
X"70ef0676",
X"842b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"bc087085",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80bc7008",
X"70df0676",
X"852b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"bc087086",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80bc7008",
X"70ffbf06",
X"76862b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80800870",
X"882c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"70892c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708a2c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708b",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"8c2cbf06",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"70922c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"0870932c",
X"810683c0",
X"800c5182",
X"3d0d0471",
X"9080a00c",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727081",
X"055434ff",
X"1151f039",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708405",
X"540cff11",
X"51f03984",
X"3d0d04fe",
X"3d0d8880",
X"53805288",
X"800a51ff",
X"b43f8280",
X"53805282",
X"800a51c8",
X"3f800b87",
X"aa803484",
X"3d0d0480",
X"3d0d8151",
X"f9d53f72",
X"802e9038",
X"8051fbd6",
X"3fc93f81",
X"e9fc3351",
X"fbcc3f81",
X"51f9e63f",
X"8051f9e1",
X"3f8051f9",
X"b23f823d",
X"0d04fd3d",
X"0d755280",
X"5480ff72",
X"25883881",
X"0bff8013",
X"5354ffbf",
X"12517099",
X"268638e0",
X"1252b039",
X"ff9f1251",
X"997127a7",
X"38d012e0",
X"13545170",
X"89268538",
X"72529839",
X"728f2685",
X"3872528f",
X"3971ba2e",
X"09810685",
X"389a5283",
X"39805273",
X"802e8538",
X"81801252",
X"7181ff06",
X"83c0800c",
X"853d0d04",
X"803d0d84",
X"98c05180",
X"71708105",
X"53347084",
X"a0c02e09",
X"8106f038",
X"823d0d04",
X"fe3d0d02",
X"97053351",
X"fef43f83",
X"c0800881",
X"ff0683c7",
X"dc085452",
X"8073249b",
X"3883c894",
X"08137283",
X"c8980807",
X"53537173",
X"3483c7dc",
X"08810583",
X"c7dc0c84",
X"3d0d04fb",
X"3d0d8056",
X"873dfc05",
X"54785379",
X"527751ff",
X"b8aa3f87",
X"3d0d04fe",
X"3d0d83c7",
X"f8085274",
X"51ffbfae",
X"3f83c080",
X"088c3876",
X"53755283",
X"c7f80851",
X"ca3f843d",
X"0d04fe3d",
X"0d83c7f8",
X"08537552",
X"7451ffb9",
X"ec3f83c0",
X"80088d38",
X"77537652",
X"83c7f808",
X"51ffa43f",
X"843d0d04",
X"f73d0d9c",
X"d23f83c0",
X"800881ff",
X"06ff0557",
X"76833881",
X"5780e9ae",
X"3f83c080",
X"0883c080",
X"08565a87",
X"15335473",
X"802e80df",
X"38740881",
X"e1c02e09",
X"810680d3",
X"38800b91",
X"16335559",
X"73792e80",
X"c6387456",
X"9a163354",
X"73832e09",
X"8106a438",
X"a4167033",
X"55588052",
X"73519abc",
X"3f805380",
X"5273519a",
X"dc3f8114",
X"54767425",
X"83388054",
X"73783481",
X"1980d817",
X"91173356",
X"57597874",
X"2e098106",
X"ffbe3881",
X"c4158ca0",
X"1b555574",
X"742e0981",
X"06ff8838",
X"8b3d0d04",
X"f63d0d80",
X"e8a03f83",
X"c080087d",
X"83c08008",
X"58595b77",
X"83c7dc0c",
X"87163355",
X"74802e81",
X"a7387508",
X"547381e5",
X"a02e0981",
X"06933890",
X"16335387",
X"16335281",
X"e69051e6",
X"fe3f8188",
X"397381e1",
X"c02e0981",
X"0680fd38",
X"745281e6",
X"a451e6e7",
X"3f807091",
X"1833565b",
X"5973792e",
X"80e638a4",
X"1657f617",
X"33557980",
X"2e9138ff",
X"15547382",
X"268938a8",
X"187083c7",
X"dc0c5874",
X"812e0981",
X"06873881",
X"e6ac518d",
X"3974822e",
X"0981068a",
X"3881e6b4",
X"51e6a03f",
X"95397483",
X"2e098106",
X"8f387633",
X"81055281",
X"e6c051e6",
X"8a3f815a",
X"811980d8",
X"18911833",
X"56585978",
X"742e0981",
X"06ff9f38",
X"a81881c4",
X"178ca01d",
X"56575875",
X"742e0981",
X"06feb838",
X"8c3d0d04",
X"803d0d72",
X"842981ea",
X"80057008",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"72842981",
X"ea9c0570",
X"0883c080",
X"0c51823d",
X"0d04f73d",
X"0d81eab0",
X"51ffbbb0",
X"3f908090",
X"08599080",
X"bc085a78",
X"57795883",
X"c7e03355",
X"74802e80",
X"ca3883c7",
X"fc085381",
X"e7905283",
X"c0800851",
X"ffb5f63f",
X"83c08008",
X"b23883c0",
X"8008568b",
X"3dec1155",
X"558853f8",
X"155283c7",
X"fc0851ff",
X"b3de3f76",
X"93f88083",
X"0679ec87",
X"fffc0607",
X"705a9080",
X"900c7990",
X"80bc0c8b",
X"3d0d04f9",
X"3d0d81ea",
X"b051ffba",
X"bf3f9080",
X"90085790",
X"80bc0858",
X"83c7e033",
X"5574802e",
X"80c63883",
X"c7fc0853",
X"81e79052",
X"83c08008",
X"51ffb589",
X"3f83c080",
X"085583c0",
X"8008a938",
X"83c08008",
X"5283c7fc",
X"0851ffb3",
X"ab3f7456",
X"893df411",
X"55558853",
X"f8155283",
X"c7fc0851",
X"ffb1af3f",
X"ffb0e73f",
X"893d0d04",
X"fd3d0d83",
X"c7f80851",
X"ffb3db3f",
X"83c08008",
X"90802e09",
X"8106ad38",
X"805487c1",
X"80805383",
X"c0800852",
X"83c7f808",
X"51f9f03f",
X"87c18080",
X"143387c1",
X"90801534",
X"81145473",
X"90802e09",
X"8106e938",
X"853d0d04",
X"fd3d0d90",
X"80805286",
X"84808051",
X"ffb4b83f",
X"805483c0",
X"8008742e",
X"098106b4",
X"3883c880",
X"085180fa",
X"b93f81ea",
X"b051ffb8",
X"eb3f83c7",
X"f8085381",
X"e79c5283",
X"c0800851",
X"ffb3ca3f",
X"83c08008",
X"742e0981",
X"068438fe",
X"eb3f8154",
X"7383c080",
X"0c853d0d",
X"0481e7a8",
X"0b83c080",
X"0c04fc3d",
X"0d765473",
X"902e8182",
X"38739024",
X"8e387384",
X"2e983873",
X"862ea738",
X"82bf3973",
X"932e8199",
X"3873942e",
X"81d43882",
X"b0398481",
X"80805382",
X"80805283",
X"c7f40851",
X"f8b53f82",
X"ba398054",
X"84818080",
X"5380c080",
X"5283c7f4",
X"0851f89f",
X"3f848280",
X"805380c0",
X"805283c7",
X"f40851f8",
X"8e3f8481",
X"80801433",
X"8481c080",
X"15348482",
X"80801433",
X"8482c080",
X"15348114",
X"547380c0",
X"802e0981",
X"06dc3881",
X"ee398482",
X"80805381",
X"80805283",
X"c7f40851",
X"f7d53f80",
X"54848280",
X"80143384",
X"81808015",
X"34811454",
X"73818080",
X"2e098106",
X"e83881bf",
X"39848180",
X"805380c0",
X"805283c7",
X"f40851f7",
X"a63f8055",
X"84818080",
X"15547333",
X"8481c080",
X"16347333",
X"84828080",
X"16347333",
X"8482c080",
X"16348115",
X"557480c0",
X"802e0981",
X"06d63880",
X"fe398481",
X"808053a0",
X"805283c7",
X"f40851f6",
X"e63f8055",
X"84818080",
X"15547333",
X"8481a080",
X"16347333",
X"8481c080",
X"16347333",
X"8481e080",
X"16347333",
X"84828080",
X"16347333",
X"8482a080",
X"16347333",
X"8482c080",
X"16347333",
X"8482e080",
X"16348115",
X"5574a080",
X"2e098106",
X"ffb6389f",
X"39f5bd3f",
X"800b83c7",
X"dc0c800b",
X"83c8980c",
X"81e7ac51",
X"dfbd3f81",
X"b78dc051",
X"f3a53f86",
X"3d0d04fc",
X"3d0d7670",
X"5255ffb6",
X"9d3f83c0",
X"80085481",
X"5383c080",
X"0880c238",
X"7451ffb5",
X"df3f83c0",
X"800881e7",
X"c85383c0",
X"80085253",
X"cebf3f83",
X"c08008a1",
X"3881e7cc",
X"527251ce",
X"b03f83c0",
X"80089238",
X"81e7d052",
X"7251cea1",
X"3f83c080",
X"08802e83",
X"38815473",
X"537283c0",
X"800c863d",
X"0d04f03d",
X"0d80de8b",
X"0b83c3ac",
X"0c83c7f4",
X"0851d0cb",
X"3f83c7f4",
X"0851ffab",
X"943fff0b",
X"81e7cc53",
X"83c08008",
X"5256cde1",
X"3f83c080",
X"08802e9f",
X"38805892",
X"3dd81155",
X"559053f0",
X"155283c7",
X"f40851ff",
X"ad863f02",
X"bb053356",
X"81a53983",
X"c7f40851",
X"ffae833f",
X"83c08008",
X"5783c080",
X"08828080",
X"2e098106",
X"83388456",
X"83c08008",
X"8180802e",
X"09810680",
X"e138805c",
X"805b805a",
X"8059f3b4",
X"3f800b83",
X"c7dc0c80",
X"0b83c898",
X"0c81e7d4",
X"51ddb43f",
X"80d00b83",
X"c7dc0c81",
X"e7e451dd",
X"a63f80f8",
X"0b83c7dc",
X"0c81e7f8",
X"51dd983f",
X"758025a2",
X"38805289",
X"3d705255",
X"8d963f83",
X"5274518d",
X"8f3f7855",
X"74802583",
X"38905680",
X"7525dd38",
X"86567680",
X"c0802e09",
X"81068538",
X"93568c39",
X"76a0802e",
X"09810683",
X"38945675",
X"51faa73f",
X"923d0d04",
X"f63d0d80",
X"5a805980",
X"58805780",
X"705656f2",
X"ab3f800b",
X"83c7dc0c",
X"800b83c8",
X"980c81e8",
X"8c51dcab",
X"3f81800b",
X"83c8980c",
X"81e89051",
X"dc9d3f80",
X"d00b83c7",
X"dc0c7430",
X"70760780",
X"2570872b",
X"83c8980c",
X"5153eaf7",
X"3f83c080",
X"085281e8",
X"9851dbf7",
X"3f80f80b",
X"83c7dc0c",
X"74813270",
X"30707207",
X"80257087",
X"2b83c898",
X"0c515454",
X"f9a33f83",
X"c0800852",
X"81e8a451",
X"dbcd3f81",
X"a00b83c7",
X"dc0c7482",
X"32703070",
X"72078025",
X"70872b83",
X"c8980c51",
X"5483c7f8",
X"085254ff",
X"a88b3f83",
X"c0800852",
X"81e8ac51",
X"db9d3f81",
X"c80b83c7",
X"dc0c7483",
X"32703070",
X"72078025",
X"70872b83",
X"c8980c51",
X"5483c7f4",
X"085254ff",
X"a7db3f81",
X"e8b45383",
X"c0800880",
X"2e8f3883",
X"c7f40851",
X"ffa7c63f",
X"83c08008",
X"53725281",
X"e8bc51da",
X"d63f81f0",
X"0b83c7dc",
X"0c748432",
X"70307072",
X"07802570",
X"872b83c8",
X"980c5154",
X"81e8c452",
X"54dab43f",
X"82c00b83",
X"c7dc0c74",
X"85327030",
X"70720780",
X"2570872b",
X"83c8980c",
X"515481e8",
X"dc5254da",
X"923f800b",
X"83c8980c",
X"839051f2",
X"cb3f868d",
X"a051edef",
X"3f805287",
X"3d705253",
X"8a823f83",
X"52725189",
X"fb3f7953",
X"7281cb38",
X"77155574",
X"80258538",
X"72559039",
X"85752585",
X"38855587",
X"39748526",
X"81aa3874",
X"842981e1",
X"a8055372",
X"0804e8b3",
X"3f83c080",
X"08775553",
X"73812e09",
X"81068938",
X"83c08008",
X"10539039",
X"73ff2e09",
X"81068838",
X"83c08008",
X"812c5390",
X"73258538",
X"90538839",
X"72802483",
X"38815372",
X"51e88d3f",
X"80de39e8",
X"9f3f83c0",
X"80081753",
X"72802585",
X"38805388",
X"39877325",
X"83388753",
X"7251e899",
X"3fbe3976",
X"86387880",
X"2eb63883",
X"c3a40883",
X"c3a00caf",
X"990b83c3",
X"ac0c83c7",
X"f80851ca",
X"d23ff4e8",
X"3f9a3978",
X"802e9538",
X"f9e83f81",
X"53963978",
X"802e8938",
X"efce3f84",
X"39788738",
X"75802efb",
X"de388053",
X"7283c080",
X"0c8c3d0d",
X"04fd3d0d",
X"83c88451",
X"80e8c23f",
X"8053ebc9",
X"3f83c080",
X"08732e09",
X"81068338",
X"8153800b",
X"83c7e033",
X"53547174",
X"2e098106",
X"83388154",
X"72812e09",
X"81069838",
X"73730652",
X"71802e8f",
X"38f4c13f",
X"83c08008",
X"863883c0",
X"80085380",
X"0b83c7e0",
X"33535471",
X"812e0981",
X"06833871",
X"5472a638",
X"73810652",
X"71802e9d",
X"387283c7",
X"e4555273",
X"70840555",
X"0851ffa4",
X"8a3f8112",
X"5271882e",
X"098106eb",
X"387283c7",
X"e034e9e0",
X"3f83c080",
X"08802e86",
X"38805180",
X"da39e9e5",
X"3f83c080",
X"0880ce38",
X"e9f03f83",
X"c0800880",
X"2eaa3881",
X"51e5903f",
X"e1ca3f80",
X"0b83c7dc",
X"0cfa813f",
X"83c08008",
X"52ff0b83",
X"c7dc0ce3",
X"dc3f71a1",
X"387151e4",
X"ee3f9f39",
X"e9d13f83",
X"c0800880",
X"2e943881",
X"51e4dc3f",
X"e1963ff7",
X"d53fe3b9",
X"3f8151ea",
X"f23f853d",
X"0d04fd3d",
X"0d805283",
X"c8845180",
X"d6fd3f82",
X"80805380",
X"52818180",
X"8051e9f1",
X"3f80c080",
X"53805284",
X"81808051",
X"ea823f80",
X"54e9ae3f",
X"83c08008",
X"83388154",
X"7383c7e0",
X"347381ff",
X"06547380",
X"2e9238f2",
X"bf3f83c0",
X"80088938",
X"83c08008",
X"83c7e034",
X"8151ea93",
X"3ffda63f",
X"fc3983c0",
X"8c080283",
X"c08c0cfb",
X"3d0d0280",
X"d3c45383",
X"c08c08fc",
X"050c8051",
X"d58e3f81",
X"e8e40b83",
X"c3a40c81",
X"e7d00b83",
X"c39c0c81",
X"e7cc0b83",
X"c3b40c81",
X"e8e80b83",
X"c3b00c81",
X"e8ec0b83",
X"c3a80c80",
X"0b83c7e4",
X"0b83c08c",
X"08f8050c",
X"83c08c08",
X"f4050cff",
X"a5893f83",
X"c0800886",
X"05fc0683",
X"c08c08f0",
X"050c0283",
X"c08c08f0",
X"0508310d",
X"833d7083",
X"c08c08f8",
X"05087084",
X"0583c08c",
X"08f8050c",
X"0c51ffa1",
X"9a3f83c0",
X"8c08f405",
X"08810583",
X"c08c08f4",
X"050c83c0",
X"8c08f405",
X"08882e09",
X"8106ffab",
X"38869480",
X"8051deda",
X"3fff0b83",
X"c7dc0c80",
X"0b83c898",
X"0c8498c0",
X"0b83c894",
X"0c8151e2",
X"9a3f8151",
X"e2bf3f80",
X"51e2ba3f",
X"8151e2e0",
X"3f8251e3",
X"883f8051",
X"e3dd3f80",
X"51e4873f",
X"8051e4b0",
X"3f8051e4",
X"d83f8051",
X"e39c3fc8",
X"0b87809a",
X"34fd9b3f",
X"83c08c08",
X"fc05080d",
X"800b83c0",
X"800c873d",
X"0d83c08c",
X"0c04fa3d",
X"0d785580",
X"750c800b",
X"84160c80",
X"0b88160c",
X"800b8c16",
X"0c800b90",
X"160c83c8",
X"845180e3",
X"b03fe6a4",
X"3f83c080",
X"0887d088",
X"337081ff",
X"06515356",
X"71a73887",
X"d0803383",
X"c8a83487",
X"d0813383",
X"c8a43487",
X"d0823383",
X"c89c3487",
X"d0833383",
X"c8a034ff",
X"0b87d08b",
X"3487d089",
X"3387d08f",
X"3370822a",
X"70810670",
X"30707207",
X"7009709f",
X"2c77069e",
X"06575151",
X"56515154",
X"54807498",
X"06535371",
X"882e0981",
X"06833881",
X"53719832",
X"70307080",
X"25757131",
X"84190c51",
X"51528074",
X"86065353",
X"71822e09",
X"81068338",
X"81537186",
X"32703070",
X"80257571",
X"31780c51",
X"515283c8",
X"a8335281",
X"aa722784",
X"3881750c",
X"83c8a833",
X"5271bb26",
X"8438ff75",
X"0c83c8a4",
X"335281aa",
X"72278638",
X"810b8416",
X"0c83c8a4",
X"335271bb",
X"268638ff",
X"0b84160c",
X"83c89c33",
X"5281aa72",
X"27843881",
X"750c83c8",
X"9c335271",
X"bb268438",
X"ff750c83",
X"c8a03352",
X"81aa7227",
X"8638810b",
X"84160c83",
X"c8a03352",
X"71bb2686",
X"38ff0b84",
X"160c8057",
X"73942eaa",
X"38878090",
X"33878091",
X"33878092",
X"337081ff",
X"06727406",
X"06878093",
X"33710681",
X"06515254",
X"54547277",
X"2e098106",
X"83388157",
X"7688160c",
X"75802eb0",
X"3875812a",
X"70810677",
X"81063184",
X"170c5275",
X"832a7682",
X"2a718106",
X"71810631",
X"770c5353",
X"75842a81",
X"0688160c",
X"75852a81",
X"068c160c",
X"883d0d04",
X"fe3d0d74",
X"76545271",
X"51fccf3f",
X"72812ea2",
X"38817326",
X"8d387282",
X"2ea83872",
X"832e9c38",
X"e6397108",
X"e2388412",
X"08dd3888",
X"1208d838",
X"a5398812",
X"08812e9e",
X"38913988",
X"1208812e",
X"95387108",
X"91388412",
X"088c388c",
X"1208812e",
X"098106ff",
X"b238843d",
X"0d04fb3d",
X"0d780284",
X"059f0533",
X"5556800b",
X"81e3ac56",
X"5381732b",
X"74065271",
X"802e8338",
X"81527470",
X"82055622",
X"7073902b",
X"0790809c",
X"0c518113",
X"5372882e",
X"098106d9",
X"38805383",
X"c8b01333",
X"517081ff",
X"2eb83870",
X"1081e1cc",
X"05702253",
X"517181ff",
X"2ea83880",
X"73177033",
X"701081e1",
X"cc057022",
X"51515152",
X"5471712e",
X"91388114",
X"5473862e",
X"098106f1",
X"38719080",
X"9c0c8113",
X"5372862e",
X"098106ff",
X"b2388053",
X"72167033",
X"51517081",
X"ff2e9a38",
X"701081e1",
X"cc057022",
X"51517081",
X"ff2e8a38",
X"70848080",
X"0790809c",
X"0c811353",
X"72862e09",
X"8106d138",
X"80537216",
X"51703383",
X"c8b01434",
X"81135372",
X"862e0981",
X"06ec3887",
X"3d0d0404",
X"fe3d0d75",
X"02840593",
X"05338106",
X"52527088",
X"38719080",
X"940c8e39",
X"70812e09",
X"81068638",
X"71908098",
X"0c843d0d",
X"04fb3d0d",
X"78982b70",
X"982c7b98",
X"2b70982c",
X"0290059f",
X"05338106",
X"83c8cc11",
X"70337098",
X"2b70982c",
X"51585c5a",
X"56515551",
X"5470742e",
X"09810694",
X"3883c8ac",
X"12337098",
X"2b70982c",
X"51525670",
X"732eb138",
X"73753472",
X"83c8ac13",
X"3483c8ad",
X"3383c8cd",
X"3371982b",
X"71902b07",
X"83c8ac33",
X"70882b72",
X"0783c8cc",
X"33710790",
X"80b80c52",
X"59535452",
X"873d0d04",
X"fe3d0d74",
X"81113371",
X"3371882b",
X"0783c080",
X"0c535184",
X"3d0d0483",
X"c8b83383",
X"c0800c04",
X"83c08c08",
X"0283c08c",
X"0cf53d0d",
X"83c08c08",
X"88050883",
X"c08c088f",
X"053383c0",
X"8c089205",
X"22028c05",
X"73900583",
X"c08c08e8",
X"050c83c0",
X"8c08f805",
X"0c83c08c",
X"08f0050c",
X"83c08c08",
X"ec050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"f0050883",
X"c08c08e0",
X"050c83c0",
X"8c08fc05",
X"0c83c08c",
X"08f00508",
X"89278a38",
X"890b83c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"860587ff",
X"fc0683c0",
X"8c08e005",
X"0c0283c0",
X"8c08e005",
X"08310d85",
X"3d705583",
X"c08c08ec",
X"05085483",
X"c08c08f0",
X"05085383",
X"c08c08f4",
X"05085283",
X"c08c08e4",
X"050c80e1",
X"b73f83c0",
X"800881ff",
X"0683c08c",
X"08e40508",
X"83c08c08",
X"ec050c83",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08802e8c",
X"3883c08c",
X"08f80508",
X"0d89c839",
X"83c08c08",
X"f0050880",
X"2e89a638",
X"83c08c08",
X"ec050881",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"842ea938",
X"840b83c0",
X"8c08e005",
X"082588c7",
X"3883c08c",
X"08e00508",
X"852e859b",
X"3883c08c",
X"08e00508",
X"a12e87ad",
X"3888ac39",
X"800b83c0",
X"8c08ec05",
X"08850533",
X"83c08c08",
X"e0050c83",
X"c08c08fc",
X"050c83c0",
X"8c08e005",
X"08832e09",
X"81068883",
X"3883c08c",
X"08e80508",
X"81053383",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08812687",
X"e638810b",
X"83c08c08",
X"e0050880",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08fc050c",
X"83c08c08",
X"ec050882",
X"053383c0",
X"8c08e005",
X"08870534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088b0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08e005",
X"088c0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088d0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08e005",
X"088e0523",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088a0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"08057094",
X"0508fcff",
X"ff067194",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08ec0508",
X"86053383",
X"c08c08e0",
X"050c83c0",
X"8c08f405",
X"0c83c08c",
X"08e00508",
X"83c08c08",
X"fc05082e",
X"098106b6",
X"3883c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08fc0508",
X"83c08c08",
X"e005088b",
X"053483c0",
X"8c08ec05",
X"08870533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508812e",
X"8f3883c0",
X"8c08e005",
X"08822eb7",
X"38848c39",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"820b83c0",
X"8c08e005",
X"088a0534",
X"83d93983",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c83",
X"c08c08fc",
X"050883c0",
X"8c08e005",
X"088a0534",
X"83a13983",
X"c08c08fc",
X"0508802e",
X"83953883",
X"c08c08ec",
X"05088305",
X"33830683",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08832e09",
X"810682f3",
X"3883c08c",
X"08ec0508",
X"82053370",
X"982b83c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"83c08c08",
X"e0050880",
X"2582cc38",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"83c08c08",
X"ec050886",
X"053383c0",
X"8c08e005",
X"0880d605",
X"3483c08c",
X"08e00508",
X"840583c0",
X"8c08ec05",
X"08820533",
X"8f0683c0",
X"8c08e405",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"e4050883",
X"c08c08e0",
X"05083483",
X"c08c08ec",
X"05088405",
X"3383c08c",
X"08e00508",
X"81053480",
X"0b83c08c",
X"08e00508",
X"82053483",
X"c08c08e0",
X"050808ff",
X"83ff0682",
X"800783c0",
X"8c08e005",
X"080c83c0",
X"8c08e805",
X"08810533",
X"810583c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"83c08c08",
X"e8050881",
X"05348183",
X"3983c08c",
X"08fc0508",
X"802e80f7",
X"3883c08c",
X"08ec0508",
X"86053383",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08a22e09",
X"810680d7",
X"3883c08c",
X"08ec0508",
X"88053383",
X"c08c08ec",
X"05088705",
X"33718280",
X"290583c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c52",
X"83c08c08",
X"e4050c83",
X"c08c08f4",
X"050c83c0",
X"8c08e405",
X"0883c08c",
X"08e00508",
X"88052383",
X"c08c08ec",
X"05083383",
X"c08c08f0",
X"05087131",
X"7083ffff",
X"0683c08c",
X"08f0050c",
X"83c08c08",
X"e0050c83",
X"c08c08ec",
X"05080583",
X"c08c08ec",
X"050cf6d0",
X"3983c08c",
X"08f80508",
X"0d83c08c",
X"08f00508",
X"83c08c08",
X"e0050c83",
X"c08c08f8",
X"05080d83",
X"c08c08e0",
X"050883c0",
X"800c8d3d",
X"0d83c08c",
X"0c0483c0",
X"8c080283",
X"c08c0ce7",
X"3d0d83c0",
X"8c088805",
X"08028405",
X"83c08c08",
X"e8050c83",
X"c08c08d4",
X"050c800b",
X"83c8d434",
X"83c08c08",
X"d4050890",
X"0583c08c",
X"08c4050c",
X"800b83c0",
X"8c08c405",
X"0834800b",
X"83c08c08",
X"c4050881",
X"0534800b",
X"83c08c08",
X"c8050c83",
X"c08c08c8",
X"050880d8",
X"2983c08c",
X"08c40508",
X"0583c08c",
X"08ffb805",
X"0c800b83",
X"c08c08ff",
X"b8050880",
X"d8050c83",
X"c08c08ff",
X"b8050884",
X"0583c08c",
X"08ffb805",
X"0c83c08c",
X"08c80508",
X"83c08c08",
X"ffb80508",
X"34880b83",
X"c08c08ff",
X"b8050881",
X"0534800b",
X"83c08c08",
X"ffb80508",
X"82053483",
X"c08c08ff",
X"b8050808",
X"ffa1ff06",
X"a0800783",
X"c08c08ff",
X"b805080c",
X"83c08c08",
X"c8050881",
X"057081ff",
X"0683c08c",
X"08c8050c",
X"83c08c08",
X"ffb8050c",
X"810b83c0",
X"8c08c805",
X"0827fedb",
X"3883c08c",
X"08ec0570",
X"5483c08c",
X"08cc050c",
X"925283c0",
X"8c08d405",
X"085180d4",
X"de3f83c0",
X"800881ff",
X"067083c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffbc",
X"050890c9",
X"3883c08c",
X"08f40551",
X"f1ca3f83",
X"c0800883",
X"ffff0683",
X"c08c08f6",
X"055283c0",
X"8c08dc05",
X"0cf1b13f",
X"83c08008",
X"83ffff06",
X"83c08c08",
X"fd053383",
X"c08c08ff",
X"bc050883",
X"c08c08c8",
X"050c83c0",
X"8c08c005",
X"0c83c08c",
X"08d8050c",
X"83c08c08",
X"c8050883",
X"c08c08c0",
X"05082780",
X"fe3883c0",
X"8c08cc05",
X"085483c0",
X"8c08c805",
X"08538952",
X"83c08c08",
X"d4050851",
X"80d3e53f",
X"83c08008",
X"81ff0683",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"bc050883",
X"eb3883c0",
X"8c08ee05",
X"51f0b13f",
X"83c08008",
X"83ffff06",
X"5383c08c",
X"08c80508",
X"5283c08c",
X"08d40508",
X"51f0b53f",
X"83c08c08",
X"c8050881",
X"057081ff",
X"0683c08c",
X"08c8050c",
X"83c08c08",
X"ffb8050c",
X"fef23983",
X"c08c08c4",
X"05088105",
X"3383c08c",
X"08c0050c",
X"83c08c08",
X"c0050883",
X"9e3883c0",
X"8c08c005",
X"0883c08c",
X"08ffb805",
X"0c83c08c",
X"08dc0508",
X"88de2e09",
X"81068b38",
X"810b83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08d805",
X"08858e2e",
X"09810682",
X"c5388170",
X"83c08c08",
X"ffb80508",
X"0683c08c",
X"08ffb805",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"ffb80508",
X"802e829e",
X"3883c08c",
X"08c80508",
X"83c08c08",
X"c4050881",
X"053483c0",
X"8c08c005",
X"0883c08c",
X"08c40508",
X"87053483",
X"c08c08c0",
X"050883c0",
X"8c08c405",
X"088b0534",
X"83c08c08",
X"c0050883",
X"c08c08c4",
X"05088c05",
X"34830b83",
X"c08c08c4",
X"05088d05",
X"3483c08c",
X"08c00508",
X"83c08c08",
X"c405088e",
X"0523830b",
X"83c08c08",
X"c405088a",
X"053483c0",
X"8c08c405",
X"08940508",
X"83808007",
X"83c08c08",
X"c4050894",
X"050c83c8",
X"b8337083",
X"c08c08c8",
X"05080583",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"b8050883",
X"c8b83483",
X"c08c08ff",
X"bc050883",
X"c08c08c4",
X"05089405",
X"3483c08c",
X"08c80508",
X"83c08c08",
X"c4050880",
X"d6053483",
X"c08c08c8",
X"050883c0",
X"8c08c405",
X"08840534",
X"8e0b83c0",
X"8c08c405",
X"08850534",
X"83c08c08",
X"c0050883",
X"c08c08c4",
X"05088605",
X"3483c08c",
X"08c40508",
X"840508ff",
X"83ff0682",
X"800783c0",
X"8c08c405",
X"0884050c",
X"a23981db",
X"0b83c08c",
X"08ffb805",
X"0c8bc639",
X"83c08c08",
X"ffbc0508",
X"83c08c08",
X"ffb8050c",
X"8bb33983",
X"c08c08f1",
X"05335283",
X"c08c08d4",
X"05085180",
X"cfea3f80",
X"0b83c08c",
X"08c40508",
X"81053383",
X"c08c08ff",
X"b8050c83",
X"c08c08c8",
X"050c83c0",
X"8c08c805",
X"0883c08c",
X"08ffb805",
X"082789ba",
X"3883c08c",
X"08c80508",
X"80d82970",
X"83c08c08",
X"c4050805",
X"70880570",
X"83053383",
X"c08c08ff",
X"b8050c83",
X"c08c08cc",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08ffb805",
X"0886fd38",
X"83c08c08",
X"ffbc0508",
X"8d053383",
X"c08c08d0",
X"050c83c0",
X"8c08d005",
X"0886e138",
X"83c08c08",
X"cc050822",
X"02840571",
X"860587ff",
X"fc0683c0",
X"8c08ffb8",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08c0050c",
X"0283c08c",
X"08ffb805",
X"08310d89",
X"3d705983",
X"c08c08c0",
X"05085883",
X"c08c08ff",
X"bc050887",
X"05335783",
X"c08c08ff",
X"b8050ca2",
X"5583c08c",
X"08d00508",
X"54865381",
X"815283c0",
X"8c08d405",
X"085180c2",
X"9d3f83c0",
X"800881ff",
X"0683c08c",
X"08d0050c",
X"83c08c08",
X"d0050881",
X"c03883c0",
X"8c08ffbc",
X"05089605",
X"5383c08c",
X"08c00508",
X"5283c08c",
X"08ffb805",
X"0851a5d5",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"802e8185",
X"3883c08c",
X"08ffbc05",
X"08940583",
X"c08c08ff",
X"bc050896",
X"05337086",
X"2a83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08c0050c",
X"83c08c08",
X"ffb80508",
X"832e0981",
X"0680c638",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"cc050882",
X"053483c8",
X"b8337081",
X"0583c08c",
X"08ffb805",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffb805",
X"0883c8b8",
X"3483c08c",
X"08ffbc05",
X"0883c08c",
X"08c00508",
X"3483c08c",
X"08e00508",
X"0d83c08c",
X"08d00508",
X"81ff0683",
X"c08c08ff",
X"bc050c83",
X"c08c08ff",
X"bc0508fb",
X"e33883c0",
X"8c08c805",
X"0883ed38",
X"83c08c08",
X"c8050883",
X"c08c08ff",
X"b8050c83",
X"c08c08dc",
X"050880f9",
X"2e098106",
X"8b38810b",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"d8050891",
X"2e098106",
X"81813883",
X"c08c08ff",
X"b8050881",
X"0683c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"08802e80",
X"e238850b",
X"83c08c08",
X"c40508a6",
X"0534a00b",
X"83c08c08",
X"c40508a7",
X"0534850b",
X"83c08c08",
X"c40508a8",
X"053480c0",
X"0b83c08c",
X"08c40508",
X"a9053486",
X"0b83c08c",
X"08c40508",
X"aa053490",
X"0b83c08c",
X"08c40508",
X"ab053486",
X"0b83c08c",
X"08c40508",
X"ac0534a0",
X"0b83c08c",
X"08c40508",
X"ad053483",
X"c08c08dc",
X"050889d8",
X"32703070",
X"80255151",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"d8050883",
X"edec2e09",
X"810680ec",
X"38817083",
X"c08c08ff",
X"b8050806",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffbc050c",
X"83c08c08",
X"ffb80508",
X"802e80c4",
X"38840b83",
X"c08c08c4",
X"0508aa05",
X"3480c00b",
X"83c08c08",
X"c40508ab",
X"0534840b",
X"83c08c08",
X"c40508ac",
X"0534900b",
X"83c08c08",
X"c40508ad",
X"053483c0",
X"8c08ffbc",
X"050883c0",
X"8c08c405",
X"088c0534",
X"83c08c08",
X"dc050880",
X"f9327030",
X"70802551",
X"5183c08c",
X"08ffb805",
X"0c83c08c",
X"08d80508",
X"862e0981",
X"06ba3881",
X"7083c08c",
X"08ffb805",
X"080683c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb8",
X"0508802e",
X"933883c0",
X"8c08ffbc",
X"050883c0",
X"8c08c405",
X"088d0534",
X"83c08c08",
X"dc0508b4",
X"b4327030",
X"70802551",
X"5183c08c",
X"08ffb805",
X"0c83c08c",
X"08d80508",
X"90892e09",
X"81069938",
X"83c08c08",
X"ffb80508",
X"802e8d38",
X"820b83c0",
X"8c08c405",
X"088d0534",
X"83c08c08",
X"e4050883",
X"c08c08c4",
X"05080570",
X"84057083",
X"053383c0",
X"8c08ffb8",
X"050c83c0",
X"8c08cc05",
X"0c83c08c",
X"08c0050c",
X"80588057",
X"83c08c08",
X"ffb80508",
X"56805580",
X"548a53a1",
X"5283c08c",
X"08d40508",
X"51bbdf3f",
X"83c08008",
X"81ff0670",
X"30709f2a",
X"5183c08c",
X"08ffb805",
X"0c83c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffbc05",
X"08a02e8c",
X"3883c08c",
X"08ffb805",
X"08f6ed38",
X"83c08c08",
X"c005088b",
X"053383c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"0508802e",
X"b33883c0",
X"8c08cc05",
X"08830533",
X"83c08c08",
X"ffb8050c",
X"80588057",
X"83c08c08",
X"ffb80508",
X"56805580",
X"548b53a1",
X"5283c08c",
X"08d40508",
X"51badb3f",
X"83c08c08",
X"c8050881",
X"057081ff",
X"0683c08c",
X"08c40508",
X"81053352",
X"83c08c08",
X"c8050c83",
X"c08c08ff",
X"b8050cf6",
X"b539800b",
X"83c08c08",
X"c8050c83",
X"c08c08c8",
X"050880d8",
X"2983c08c",
X"08d40508",
X"05709a05",
X"3383c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffbc05",
X"08822e09",
X"8106bd38",
X"83c08c08",
X"ffb80508",
X"97053383",
X"c8d45983",
X"c08c08ff",
X"b8050c81",
X"5783c08c",
X"08ffb805",
X"085683c0",
X"8c08ffbc",
X"05085580",
X"548953a1",
X"5283c08c",
X"08d40508",
X"51b9b73f",
X"83c08c08",
X"c8050881",
X"057081ff",
X"0683c08c",
X"08c8050c",
X"83c08c08",
X"ffb8050c",
X"810b83c0",
X"8c08c805",
X"0827fee7",
X"38810b83",
X"c08c08c4",
X"05083480",
X"0b83c08c",
X"08ffb805",
X"0c83c08c",
X"08e80508",
X"0d83c08c",
X"08ffb805",
X"0883c080",
X"0c9b3d0d",
X"83c08c0c",
X"04f43d0d",
X"901f5980",
X"0b811a33",
X"555b7a74",
X"2781ad38",
X"7a80d829",
X"198a1133",
X"55557383",
X"2e098106",
X"81883894",
X"15335780",
X"527651df",
X"9b3f8053",
X"80527651",
X"dfbb3fad",
X"b93f83c0",
X"80085c80",
X"587781c4",
X"291c8711",
X"33555573",
X"802e80c0",
X"38740881",
X"e1c02e09",
X"8106b538",
X"80755b56",
X"7580d829",
X"1a9a1133",
X"55557383",
X"2e098106",
X"9238a415",
X"70335555",
X"76742787",
X"38ff1454",
X"73753481",
X"167081ff",
X"06575481",
X"7627d138",
X"81187081",
X"ff065954",
X"877827ff",
X"a43883c8",
X"b833ff05",
X"547383c8",
X"b834811b",
X"7081ff06",
X"811b335f",
X"5c547c7b",
X"26fed538",
X"800b83c0",
X"800c8e3d",
X"0d0483c0",
X"8c080283",
X"c08c0cda",
X"3d0d83c0",
X"8c088805",
X"08028405",
X"71900570",
X"337083c0",
X"8c08fef8",
X"050c83c0",
X"8c08fef4",
X"050c83c0",
X"8c08ff9c",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffb0",
X"050c83c0",
X"8c08fef4",
X"0508802e",
X"9a963880",
X"0b83c08c",
X"08ff9c05",
X"08810533",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"fef40508",
X"2599db38",
X"83c08c08",
X"ffa40508",
X"80d82983",
X"c08c08ff",
X"9c050805",
X"84057086",
X"053383c0",
X"8c08fef4",
X"050c83c0",
X"8c08ff88",
X"050c83c0",
X"8c08fef4",
X"0508802e",
X"98e138aa",
X"dd3f83c0",
X"8c08ff88",
X"050880d4",
X"050883c0",
X"80082698",
X"ca380283",
X"c08c08ff",
X"88050881",
X"053383c0",
X"8c08fef4",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08fef4",
X"050883c0",
X"8c08fc05",
X"2383c08c",
X"08fef405",
X"08860583",
X"fc0683c0",
X"8c08fef4",
X"050c0283",
X"c08c08fe",
X"f4050831",
X"0d853d70",
X"5583c08c",
X"08fc0554",
X"83c08c08",
X"ff880508",
X"5383c08c",
X"08ffb005",
X"085283c0",
X"8c08ff90",
X"050cb2ae",
X"3f83c080",
X"0881ff06",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"fef40508",
X"978f3883",
X"c08c08ff",
X"88050887",
X"053383c0",
X"8c08fef4",
X"050c83c0",
X"8c08fef4",
X"0508802e",
X"80d73883",
X"c08c08ff",
X"88050886",
X"053383c0",
X"8c08fef4",
X"050c83c0",
X"8c08fef4",
X"0508822e",
X"098106b5",
X"3883c08c",
X"08fc0522",
X"83c08c08",
X"fef4050c",
X"870b83c0",
X"8c08fef4",
X"05082799",
X"3883c08c",
X"08ff9005",
X"08820552",
X"83c08c08",
X"ff900508",
X"3351d8d6",
X"3f83c08c",
X"08ff8805",
X"08860533",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"fef40508",
X"832e0981",
X"0695f638",
X"83c08c08",
X"ff880508",
X"920583c0",
X"8c08ff88",
X"05088905",
X"3383c08c",
X"08fef405",
X"0c83c08c",
X"08ff9405",
X"0c83c08c",
X"08fef405",
X"08832eb7",
X"3883c08c",
X"08ff9405",
X"08820533",
X"83c08c08",
X"fc052283",
X"c08c08fe",
X"fc050c83",
X"c08c08fe",
X"f8050c83",
X"c08c08fe",
X"f8050883",
X"c08c08fe",
X"fc050826",
X"958f3880",
X"0b83c08c",
X"08ffb405",
X"0c800b83",
X"c08c08ff",
X"8c050c83",
X"c08c08fe",
X"f4050883",
X"2e098106",
X"83983883",
X"c08c08ff",
X"90050833",
X"83c08c08",
X"fef8050c",
X"83c08c08",
X"fef80508",
X"83c08c08",
X"ff8c0508",
X"2e098106",
X"82d93883",
X"c08c08ff",
X"90050881",
X"053383c0",
X"8c08fef4",
X"050c83c0",
X"8c08fef4",
X"0508942e",
X"09810682",
X"b638b053",
X"81e4b452",
X"83c08c08",
X"c8055180",
X"c7803f83",
X"c08c08fe",
X"f8050883",
X"c08c08ff",
X"8c050c83",
X"c08c08ff",
X"8c050810",
X"83c08c08",
X"ff8c0508",
X"0583c08c",
X"0805c805",
X"703383c0",
X"8c08ff90",
X"05080570",
X"33728105",
X"33710651",
X"5183c08c",
X"08fef405",
X"0c83c08c",
X"08fef805",
X"0c83c08c",
X"08fef405",
X"08802ea8",
X"3883c08c",
X"08fef805",
X"08820533",
X"81712b83",
X"c08c08ff",
X"b4050807",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"fef8050c",
X"83c08c08",
X"ff8c0508",
X"81057081",
X"ff0683c0",
X"8c08ff8c",
X"050c83c0",
X"8c08fef4",
X"050c83c0",
X"8c08ff8c",
X"0508902e",
X"098106fe",
X"e23883c0",
X"8c08ff90",
X"05088705",
X"3370982b",
X"83c08c08",
X"ff900508",
X"89053370",
X"982b7098",
X"2c73982c",
X"81800554",
X"515383c0",
X"8c08fefc",
X"050c83c0",
X"8c08fef8",
X"050c83c0",
X"8c08fef4",
X"050c83c0",
X"8c08fef8",
X"050883c0",
X"8c08f805",
X"2380ff0b",
X"83c08c08",
X"fef40508",
X"3183c08c",
X"08fef405",
X"0c83c08c",
X"08fef405",
X"0883c08c",
X"08fa0523",
X"84d73981",
X"800b83c0",
X"8c08f805",
X"2381800b",
X"83c08c08",
X"fa052384",
X"c03983c0",
X"8c08ff8c",
X"05081083",
X"c08c0805",
X"f80583c0",
X"8c08ff8c",
X"05088429",
X"83c08c08",
X"ff8c0508",
X"100583c0",
X"8c08ff94",
X"05080570",
X"84057033",
X"83c08c08",
X"ff900508",
X"05703383",
X"c08c08ff",
X"80050c83",
X"c08c08fe",
X"f4050c83",
X"c08c08fe",
X"f8050c83",
X"c08c08fe",
X"fc050c83",
X"c08c08ff",
X"84050c83",
X"c08c08ff",
X"80050883",
X"c08c08ff",
X"84050823",
X"83c08c08",
X"fef80508",
X"81053383",
X"c08c08fe",
X"f4050c83",
X"c08c08fe",
X"f4050890",
X"2e098106",
X"bf3883c0",
X"8c08fef8",
X"05083383",
X"c08c08ff",
X"90050805",
X"81057033",
X"70828029",
X"83c08c08",
X"ff800508",
X"05515183",
X"c08c08fe",
X"f4050c83",
X"c08c08fe",
X"f4050883",
X"c08c08ff",
X"84050823",
X"83c08c08",
X"fefc0508",
X"86052283",
X"c08c08fe",
X"f8050c83",
X"c08c08fe",
X"f80508a2",
X"3883c08c",
X"08fefc05",
X"08880522",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"fef40508",
X"81ff2e80",
X"e53883c0",
X"8c08ff84",
X"05082270",
X"83c08c08",
X"fef80508",
X"31708280",
X"29713183",
X"c08c08fe",
X"fc050888",
X"05227083",
X"c08c08fe",
X"f8050831",
X"70733553",
X"83c08c08",
X"fef8050c",
X"83c08c08",
X"fefc050c",
X"5183c08c",
X"08fef405",
X"0c83c08c",
X"08ff8005",
X"0c83c08c",
X"08fef405",
X"0883c08c",
X"08ff8405",
X"082383c0",
X"8c08ff8c",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ff8c050c",
X"83c08c08",
X"fef4050c",
X"810b83c0",
X"8c08ff8c",
X"050827fc",
X"dd38800b",
X"83c08c08",
X"ff8c050c",
X"83c08c08",
X"ff8c0508",
X"1083c08c",
X"08ff9405",
X"08057090",
X"05703383",
X"c08c08ff",
X"90050805",
X"70337281",
X"05337072",
X"06515351",
X"83c08c08",
X"fef8050c",
X"5183c08c",
X"08fef405",
X"0c83c08c",
X"08fef405",
X"08802e9d",
X"38900b83",
X"c08c08ff",
X"8c05082b",
X"83c08c08",
X"ffb40508",
X"0783c08c",
X"08ffb405",
X"0c83c08c",
X"08ff8c05",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"8c050c83",
X"c08c08fe",
X"f4050c97",
X"0b83c08c",
X"08ff8c05",
X"0827fef0",
X"3883c08c",
X"08f80522",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"fef40508",
X"bf269338",
X"83c08c08",
X"ffb40508",
X"820783c0",
X"8c08ffb4",
X"050c81c0",
X"0b83c08c",
X"08fef405",
X"08279338",
X"83c08c08",
X"ffb40508",
X"810783c0",
X"8c08ffb4",
X"050c83c0",
X"8c08fa05",
X"2283c08c",
X"08fef405",
X"0c83c08c",
X"08fef405",
X"08bf2693",
X"3883c08c",
X"08ffb405",
X"08880783",
X"c08c08ff",
X"b4050c81",
X"c00b83c0",
X"8c08fef4",
X"05082793",
X"3883c08c",
X"08ffb405",
X"08840783",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"88050890",
X"053383c0",
X"8c08ffb4",
X"050883c0",
X"8c08fef4",
X"050c83c0",
X"8c08ff94",
X"050c83c0",
X"8c08fef4",
X"050883c0",
X"8c08ff88",
X"05088c05",
X"082e85e9",
X"3883c08c",
X"08fef405",
X"0883c08c",
X"08ff8805",
X"088c050c",
X"83c08c08",
X"ff880508",
X"89053383",
X"c08c08fe",
X"f8050c83",
X"c08c08fe",
X"f8050880",
X"2e85a138",
X"83c08c08",
X"ffb40583",
X"c08c08fe",
X"f4050883",
X"c08c08fe",
X"f405088f",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08ff8005",
X"0c83c08c",
X"08ffa005",
X"0c83c08c",
X"08fef805",
X"08822e09",
X"810681c2",
X"38800b83",
X"c08c08fe",
X"f4050886",
X"2a708106",
X"5183c08c",
X"08fef405",
X"0c83c08c",
X"08fef805",
X"0c83c08c",
X"08fef405",
X"0883c08c",
X"08fef805",
X"082e8c38",
X"81c00b83",
X"c08c08fe",
X"f8050c83",
X"c08c08ff",
X"80050887",
X"2a708106",
X"5183c08c",
X"08fef405",
X"0c83c08c",
X"08fef405",
X"08802e94",
X"3883c08c",
X"08fef805",
X"08819032",
X"83c08c08",
X"fef8050c",
X"83c08c08",
X"ff800508",
X"842a7081",
X"065183c0",
X"8c08fef4",
X"050c83c0",
X"8c08fef4",
X"0508802e",
X"943883c0",
X"8c08fef8",
X"050880d0",
X"3283c08c",
X"08fef805",
X"0c83c08c",
X"08ff8005",
X"0883c08c",
X"08fef805",
X"083283c0",
X"8c08ff80",
X"050c800b",
X"83c08c08",
X"c0050c80",
X"0b83c08c",
X"08c40523",
X"800b81e3",
X"bc3383c0",
X"8c08fef4",
X"050c83c0",
X"8c08ff8c",
X"050c83c0",
X"8c08fef4",
X"050883c0",
X"8c08ff8c",
X"05082e82",
X"d73883c0",
X"8c08c005",
X"81e3bc0b",
X"83c08c08",
X"fefc050c",
X"83c08c08",
X"ff98050c",
X"83c08c08",
X"fefc0508",
X"3383c08c",
X"08fefc05",
X"08810533",
X"81722b81",
X"722b0770",
X"83c08c08",
X"ff800508",
X"065383c0",
X"8c08fef8",
X"050c83c0",
X"8c08ff84",
X"050c83c0",
X"8c08fef4",
X"050c83c0",
X"8c08fef4",
X"050883c0",
X"8c08fef8",
X"05082e09",
X"810681c1",
X"3883c08c",
X"08ff8c05",
X"08852680",
X"f73883c0",
X"8c08fefc",
X"05088205",
X"337081ff",
X"0683c08c",
X"08fef405",
X"0c83c08c",
X"08ff8405",
X"0c83c08c",
X"08fef405",
X"08802e80",
X"cb3883c0",
X"8c08ff8c",
X"050883c0",
X"8c08ff8c",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ff980508",
X"73055383",
X"c08c08ff",
X"8c050c83",
X"c08c08fe",
X"f8050c83",
X"c08c08fe",
X"f4050c83",
X"c08c08ff",
X"84050883",
X"c08c08fe",
X"f4050834",
X"83c08c08",
X"fefc0508",
X"83053383",
X"c08c08fe",
X"f4050c83",
X"c08c08fe",
X"f4050880",
X"2e9f3881",
X"0b83c08c",
X"08fef405",
X"082b83c0",
X"8c08ffa0",
X"05080807",
X"83c08c08",
X"ffa00508",
X"0c83c08c",
X"08fefc05",
X"08840570",
X"3383c08c",
X"08fef405",
X"0c83c08c",
X"08fefc05",
X"0c83c08c",
X"08fef405",
X"08fdc538",
X"83c08c08",
X"c0055280",
X"51c8ab3f",
X"83c08c08",
X"ffb40508",
X"5283c08c",
X"08ff9405",
X"0851c9f0",
X"3f83c08c",
X"08fb0533",
X"7081800a",
X"29810a05",
X"70982c55",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"f9053370",
X"81800a29",
X"810a0570",
X"982c5583",
X"c08c08fe",
X"f4050c83",
X"c08c08ff",
X"94050853",
X"83c08c08",
X"fefc050c",
X"83c08c08",
X"fef8050c",
X"c9c73f83",
X"c08c08ff",
X"88050888",
X"053383c0",
X"8c08fef4",
X"050c83c0",
X"8c08fef4",
X"0508802e",
X"84e73883",
X"c08c08ff",
X"88050890",
X"053383c0",
X"8c08fef4",
X"050c83c0",
X"8c08fef4",
X"05088126",
X"84c73880",
X"7081e3f4",
X"0b81e3f4",
X"0b810533",
X"83c08c08",
X"fef4050c",
X"83c08c08",
X"fef8050c",
X"83c08c08",
X"fefc050c",
X"83c08c08",
X"ff84050c",
X"83c08c08",
X"fef40508",
X"83c08c08",
X"ff840508",
X"2e81af38",
X"83c08c08",
X"fefc0508",
X"842983c0",
X"8c08fef8",
X"05080570",
X"3383c08c",
X"08ff9005",
X"08057033",
X"72810533",
X"70720651",
X"535183c0",
X"8c08fef8",
X"050c83c0",
X"8c08fef4",
X"050c83c0",
X"8c08fef4",
X"0508802e",
X"aa38810b",
X"83c08c08",
X"fefc0508",
X"2b83c08c",
X"08ff8405",
X"08077083",
X"ffff0683",
X"c08c08ff",
X"84050c83",
X"c08c08fe",
X"f4050c83",
X"c08c08fe",
X"fc050881",
X"057081ff",
X"0681e3f4",
X"71842971",
X"05708105",
X"33515383",
X"c08c08fe",
X"f8050c83",
X"c08c08fe",
X"fc050c83",
X"c08c08fe",
X"f4050c83",
X"c08c08fe",
X"f40508fe",
X"d33883c0",
X"8c08ff88",
X"05088a05",
X"2283c08c",
X"08ff9005",
X"0c83c08c",
X"08ff8405",
X"0883c08c",
X"08ff9005",
X"082e82b1",
X"38800b83",
X"c08c08ff",
X"b8050c80",
X"0b83c08c",
X"08ffbc05",
X"23807083",
X"c08c08ff",
X"b80583c0",
X"8c08ff8c",
X"050c83c0",
X"8c08fefc",
X"050c83c0",
X"8c08ff80",
X"050c81af",
X"3983c08c",
X"08ff8405",
X"0883c08c",
X"08fefc05",
X"082c7081",
X"065183c0",
X"8c08fef4",
X"050c83c0",
X"8c08fef4",
X"0508802e",
X"80e73883",
X"c08c08ff",
X"80050883",
X"c08c08ff",
X"80050881",
X"057081ff",
X"0683c08c",
X"08ff8c05",
X"08730583",
X"c08c08ff",
X"88050890",
X"053383c0",
X"8c08fefc",
X"05088429",
X"05535383",
X"c08c08ff",
X"80050c83",
X"c08c08fe",
X"f8050c83",
X"c08c08fe",
X"f4050c83",
X"c08c08fe",
X"f8050881",
X"e3f60533",
X"83c08c08",
X"fef40508",
X"3483c08c",
X"08fefc05",
X"08810570",
X"81ff0683",
X"c08c08fe",
X"fc050c83",
X"c08c08fe",
X"f4050c8f",
X"0b83c08c",
X"08fefc05",
X"082783c0",
X"8c08fef4",
X"050c83c0",
X"8c08ff80",
X"05088526",
X"8c3883c0",
X"8c08fef4",
X"0508fea9",
X"3883c08c",
X"08ffb805",
X"528051c2",
X"d13f83c0",
X"8c08ff84",
X"050883c0",
X"8c08ff88",
X"05088a05",
X"2383c08c",
X"08ff8805",
X"0880d205",
X"3383c08c",
X"08ff8805",
X"0880d405",
X"080583c0",
X"8c08ff88",
X"050880d4",
X"050c83c0",
X"8c08ffa8",
X"05080d83",
X"c08c08ff",
X"a4050881",
X"800a2981",
X"800a0570",
X"982c83c0",
X"8c08ff9c",
X"05088105",
X"3383c08c",
X"08fef805",
X"0c5183c0",
X"8c08ffa4",
X"050c83c0",
X"8c08fef8",
X"050883c0",
X"8c08ffa4",
X"050824e6",
X"a738800b",
X"83c08c08",
X"fef8050c",
X"83c08c08",
X"ffac0508",
X"0d83c08c",
X"08fef805",
X"0883c080",
X"0ca83d0d",
X"83c08c0c",
X"04e93d0d",
X"696c0288",
X"0580ea05",
X"225c5a5b",
X"80707141",
X"5e58ff78",
X"797a7b7c",
X"7d464c4a",
X"45405d43",
X"62993d34",
X"62028405",
X"80dd0534",
X"77792280",
X"ffff0654",
X"45727923",
X"79782e88",
X"87387a70",
X"81055c33",
X"70842a71",
X"8c067082",
X"2a5a5656",
X"8306ff1b",
X"7083ffff",
X"065c5456",
X"80547574",
X"2e91387a",
X"7081055c",
X"33ff1b70",
X"83ffff06",
X"5c545481",
X"76279b38",
X"7381ff06",
X"7b708105",
X"5d335574",
X"82802905",
X"ff1b7083",
X"ffff065c",
X"54548276",
X"27aa3873",
X"83ffff06",
X"7b708105",
X"5d337090",
X"2b72077d",
X"7081055f",
X"3370982b",
X"7207fe1f",
X"7083ffff",
X"06405252",
X"52525454",
X"7e802e80",
X"c4387686",
X"f738748a",
X"2e098106",
X"9438811f",
X"7081ff06",
X"811e7081",
X"ff065f52",
X"405386dc",
X"39748c2e",
X"09810686",
X"d338ff1f",
X"7081ff06",
X"ff1e7081",
X"ff065f52",
X"40537b63",
X"2586bd38",
X"ff4386b8",
X"3976812e",
X"83bb3876",
X"81248938",
X"76802e8d",
X"3886a539",
X"76822e84",
X"a638869c",
X"39f81553",
X"72842684",
X"95387284",
X"2981e4e4",
X"05537208",
X"0464802e",
X"80cd3878",
X"22838080",
X"06537283",
X"80802e09",
X"8106bc38",
X"80567564",
X"27a43875",
X"1e7083ff",
X"ff067710",
X"1b901172",
X"832a5851",
X"57515373",
X"75347287",
X"0681712b",
X"51537281",
X"16348116",
X"7081ff06",
X"57539776",
X"27cc387f",
X"84074080",
X"0b993d43",
X"56611670",
X"3370982b",
X"70982c51",
X"51515380",
X"732480fb",
X"38607329",
X"1e7083ff",
X"ff067a22",
X"83808006",
X"52585372",
X"8380802e",
X"09810680",
X"de386088",
X"32703070",
X"72078025",
X"63903270",
X"30707207",
X"80257307",
X"53545851",
X"55537380",
X"2ebd3876",
X"87065372",
X"b6387584",
X"29761005",
X"79118411",
X"79832a57",
X"57515373",
X"75346081",
X"16346586",
X"14236688",
X"14237587",
X"387f8107",
X"408d3975",
X"812e0981",
X"0685387f",
X"82074081",
X"167081ff",
X"06575381",
X"7627fee5",
X"38636129",
X"1e7083ff",
X"ff065f53",
X"80704642",
X"ff028405",
X"80dd0534",
X"ff0b993d",
X"3483f539",
X"811c7081",
X"ff065d53",
X"80427381",
X"2e098106",
X"8e387781",
X"800a2981",
X"800a0558",
X"80d33973",
X"802e8938",
X"73822e09",
X"81068d38",
X"7c81800a",
X"2981800a",
X"055da439",
X"815f83b8",
X"39ff1c70",
X"81ff065d",
X"537b6325",
X"8338ff43",
X"7c802e92",
X"387c8180",
X"0a2981ff",
X"0a055d7c",
X"982c5d83",
X"93397780",
X"2e923877",
X"81800a29",
X"81ff0a05",
X"5877982c",
X"5882fd39",
X"7753839e",
X"39748926",
X"80f43874",
X"842981e4",
X"f8055372",
X"08047387",
X"2e82e138",
X"73852e82",
X"db387388",
X"2e82d538",
X"738c2e82",
X"cf387389",
X"2e098106",
X"86388145",
X"82c23973",
X"812e0981",
X"0682b938",
X"62802582",
X"b3387b98",
X"2b70982c",
X"514382a8",
X"397383ff",
X"ff064682",
X"9f397383",
X"ffff0647",
X"82963973",
X"81ff0641",
X"828e3973",
X"811a3482",
X"87397381",
X"ff064481",
X"ff397e53",
X"82a03974",
X"812e81e3",
X"38748124",
X"89387480",
X"2e8d3881",
X"e7397482",
X"2e81d838",
X"81de3974",
X"567b8338",
X"81567453",
X"73862e09",
X"81069738",
X"75810653",
X"72802e8e",
X"38782282",
X"ffff06fe",
X"80800753",
X"b6397b83",
X"38815373",
X"822e0981",
X"06973872",
X"81065372",
X"802e8e38",
X"782281ff",
X"ff068180",
X"80075393",
X"397b9638",
X"fc145372",
X"81268e38",
X"7822ff80",
X"80075372",
X"792380e5",
X"39805573",
X"812e0981",
X"06833873",
X"55775377",
X"802e8938",
X"74810653",
X"7280ca38",
X"72d01554",
X"55728126",
X"83388155",
X"77802eb9",
X"38748106",
X"5372802e",
X"b0387822",
X"83808006",
X"53728380",
X"802e0981",
X"069f3873",
X"b02e0981",
X"06873861",
X"993d3491",
X"3973b12e",
X"09810689",
X"38610284",
X"0580dd05",
X"34618105",
X"538c3961",
X"74318105",
X"53843961",
X"14537283",
X"ffff0642",
X"79f7fb38",
X"7d832a53",
X"72821a34",
X"78228380",
X"80065372",
X"8380802e",
X"09810688",
X"3881537f",
X"872e8338",
X"80537283",
X"c0800c99",
X"3d0d04fd",
X"3d0d7583",
X"11338212",
X"3371982b",
X"71902b07",
X"81143370",
X"882b7207",
X"75337107",
X"83c0800c",
X"52535456",
X"5452853d",
X"0d04f63d",
X"0d02b705",
X"33028405",
X"bb053302",
X"8805bf05",
X"335b5b5b",
X"80588057",
X"78882b7a",
X"07568055",
X"7a548153",
X"a3527c51",
X"92c83f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f63d",
X"0d02b705",
X"33028405",
X"bb053302",
X"8805bf05",
X"335b5b5b",
X"80588057",
X"78882b7a",
X"07568055",
X"7a548353",
X"a3527c51",
X"928c3f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f73d",
X"0d02b305",
X"33028405",
X"b6052260",
X"5a585680",
X"55805480",
X"5381a352",
X"7b5191de",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8b3d0d04",
X"ee3d0d64",
X"90115c5c",
X"807b3480",
X"0b841c0c",
X"800b881c",
X"34810b89",
X"1c34880b",
X"8a1c3480",
X"0b8b1c34",
X"881b08c1",
X"06810788",
X"1c0c8f3d",
X"70545d88",
X"527b519c",
X"8e3f83c0",
X"800881ff",
X"06705b59",
X"7881a938",
X"903d335e",
X"81db5a7d",
X"892e0981",
X"06819938",
X"7c539252",
X"7b519be7",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"8182387c",
X"58885778",
X"56a95578",
X"54865381",
X"a0527b51",
X"90cc3f83",
X"c0800881",
X"ff06705b",
X"597880e0",
X"3802ba05",
X"337b347c",
X"5478537d",
X"527b519b",
X"cf3f83c0",
X"800881ff",
X"06705b59",
X"7880c138",
X"02bd0533",
X"527b519b",
X"e73f83c0",
X"800881ff",
X"06705b59",
X"78aa3881",
X"7b335a5a",
X"79792699",
X"38805479",
X"5388527b",
X"51fdbb3f",
X"811a7081",
X"ff067c33",
X"525b59e4",
X"39810b88",
X"1c34805a",
X"7983c080",
X"0c943d0d",
X"04800b83",
X"c0800c04",
X"f93d0d79",
X"028405ab",
X"05338e3d",
X"70545858",
X"58ffb7cc",
X"3f8a3d8a",
X"0551ffb7",
X"c33f7551",
X"fc8d3f83",
X"c0800884",
X"86812ebe",
X"3883c080",
X"08848681",
X"26993883",
X"c0800884",
X"82802e80",
X"e63883c0",
X"80088482",
X"812e9f38",
X"81b43983",
X"c0800880",
X"c082832e",
X"80f43883",
X"c0800880",
X"c086832e",
X"80e83881",
X"993983c0",
X"a4335580",
X"5674762e",
X"09810681",
X"8b387454",
X"76539152",
X"7751fbd6",
X"3f745476",
X"53905277",
X"51fbcb3f",
X"74547653",
X"84527751",
X"fbfc3f81",
X"0b83c0a4",
X"3481b156",
X"80de3980",
X"54765391",
X"527751fb",
X"a93f8054",
X"76539052",
X"7751fb9e",
X"3f800b83",
X"c0a43476",
X"52871833",
X"5197923f",
X"b5398054",
X"76539452",
X"7751fb82",
X"3f805476",
X"53905277",
X"51faf73f",
X"7551ffb5",
X"f73f83c0",
X"8008892a",
X"81065376",
X"52871833",
X"5190c93f",
X"800b83c0",
X"a4348056",
X"7583c080",
X"0c893d0d",
X"04f23d0d",
X"6090115a",
X"58800b88",
X"1a337159",
X"56567476",
X"2e82a538",
X"82ac3f84",
X"190883c0",
X"80082682",
X"95387833",
X"5a810b8e",
X"3d23903d",
X"f81155f4",
X"05539918",
X"5277518a",
X"e13f83c0",
X"800881ff",
X"06705755",
X"74772e09",
X"810681d9",
X"38863974",
X"5681d239",
X"81568257",
X"8e3d3377",
X"06557480",
X"2ebb3880",
X"0b8d3d34",
X"903df005",
X"54845375",
X"527751fa",
X"cd3f83c0",
X"800881ff",
X"0655749d",
X"387b5375",
X"527751fc",
X"e73f83c0",
X"800881ff",
X"06557481",
X"b12e818b",
X"3874ffb3",
X"38761081",
X"fc068117",
X"7081ff06",
X"58565787",
X"7627ffa8",
X"38815675",
X"7a2680eb",
X"38800b8d",
X"3d348c3d",
X"70555784",
X"53755277",
X"51f9f73f",
X"83c08008",
X"81ff0655",
X"7480c138",
X"7651ffb3",
X"f33f83c0",
X"80088287",
X"06557482",
X"812e0981",
X"06aa3802",
X"ae053381",
X"07557402",
X"8405ae05",
X"347b5375",
X"527751fb",
X"eb3f83c0",
X"800881ff",
X"06557481",
X"b12e9038",
X"74feb838",
X"81167081",
X"ff065755",
X"ff913980",
X"567581ff",
X"0656973f",
X"83c08008",
X"8fd00584",
X"1a0c7557",
X"7683c080",
X"0c903d0d",
X"0404803d",
X"0d9080a0",
X"08708a2c",
X"83c0800c",
X"51823d0d",
X"040483c8",
X"d80b83c0",
X"800c04fd",
X"3d0d7577",
X"5454800b",
X"83c8b834",
X"728a3890",
X"90800b84",
X"150c9039",
X"72812e09",
X"81068838",
X"9098800b",
X"84150c84",
X"140883c8",
X"d00c800b",
X"88150c80",
X"0b8c150c",
X"83c8d008",
X"53820b87",
X"80143487",
X"e851ff92",
X"b23f83c8",
X"d0085380",
X"0b881434",
X"83c8d008",
X"53810b87",
X"80143483",
X"c8d00853",
X"800b8c14",
X"3483c8d0",
X"0853800b",
X"a4143491",
X"7434800b",
X"83c0a834",
X"800b83c0",
X"ac34800b",
X"83c0b034",
X"80547381",
X"c42983c8",
X"dc055380",
X"0b831434",
X"81147081",
X"ff065553",
X"877427e6",
X"38853d0d",
X"04fe3d0d",
X"74768211",
X"3370bf06",
X"81712bff",
X"05565151",
X"52539071",
X"278338ff",
X"52765171",
X"712383c8",
X"d0085187",
X"13339012",
X"34800b83",
X"c0ac3480",
X"0b83c0b0",
X"34881333",
X"8a143352",
X"5271802e",
X"aa387081",
X"ff065184",
X"52708338",
X"70527183",
X"c0ac348a",
X"13337030",
X"70802584",
X"2b708807",
X"51515253",
X"7083c0b0",
X"34903970",
X"81ff0651",
X"70833898",
X"527183c0",
X"b034800b",
X"83c0800c",
X"843d0d04",
X"f13d0d61",
X"6568028c",
X"0580cb05",
X"33029005",
X"80ce0522",
X"02940580",
X"d6052242",
X"40415a40",
X"40fd8f3f",
X"83c08008",
X"a788055b",
X"8070715b",
X"5b528394",
X"3983c8d0",
X"08517d94",
X"123483c0",
X"ac338107",
X"55807054",
X"567f8626",
X"80ea387f",
X"842981e5",
X"ac0583c8",
X"d0085351",
X"70080480",
X"0b841334",
X"a1397733",
X"70307080",
X"25837131",
X"51515253",
X"70841334",
X"8d39810b",
X"841334b8",
X"39830b84",
X"13348170",
X"5456ad39",
X"810b8413",
X"34a23977",
X"33703070",
X"80258371",
X"31515152",
X"53708413",
X"34807833",
X"52527083",
X"38815271",
X"78348153",
X"74880755",
X"83c0b033",
X"83c8d008",
X"5257810b",
X"81d01234",
X"83c8d008",
X"51810b81",
X"9012347e",
X"802eae38",
X"72802ea9",
X"387eff1e",
X"52547083",
X"ffff0653",
X"7283ffff",
X"2e973873",
X"70810555",
X"3383c8d0",
X"08535170",
X"81c01334",
X"ff1351de",
X"3983c8d0",
X"08a81133",
X"53517688",
X"123483c8",
X"d0085174",
X"713481ff",
X"52913983",
X"c8d008a0",
X"11337081",
X"06515253",
X"708f38fb",
X"813f7a83",
X"c0800826",
X"e6388188",
X"39810ba0",
X"143483c8",
X"d008a811",
X"3380ff06",
X"70780752",
X"53517080",
X"2e80ed38",
X"71862a70",
X"81065151",
X"70802e91",
X"38807833",
X"52537083",
X"38815372",
X"783480e0",
X"3971842a",
X"70810651",
X"5170802e",
X"9b388119",
X"7083ffff",
X"067d3070",
X"9f2a5152",
X"5a51787c",
X"2e098106",
X"af38a439",
X"71832a70",
X"81065151",
X"70802e93",
X"38811a70",
X"81ff065b",
X"5179832e",
X"09810690",
X"388a3971",
X"a3065170",
X"802e8538",
X"71519239",
X"f9e83f7a",
X"83c08008",
X"26fce238",
X"7181bf06",
X"517083c0",
X"800c913d",
X"0d04f63d",
X"0d02b305",
X"33028405",
X"b7053302",
X"8805ba05",
X"22595959",
X"800b8c3d",
X"348c3dfc",
X"05568055",
X"80547653",
X"77527851",
X"fbf23f83",
X"c0800881",
X"ff0683c0",
X"800c8c3d",
X"0d04f33d",
X"0d7f6264",
X"028c0580",
X"c2052272",
X"22811533",
X"425f415e",
X"59598078",
X"237d5378",
X"33528151",
X"ffa03f83",
X"c0800881",
X"ff065675",
X"802e8638",
X"755481ad",
X"3983c8d0",
X"08a81133",
X"821b3370",
X"862a7081",
X"0673982b",
X"5351575c",
X"56577980",
X"25833881",
X"5673762e",
X"873881f0",
X"54818239",
X"818c1733",
X"7081ff06",
X"79227d71",
X"31902b70",
X"902c7009",
X"709f2c72",
X"06705252",
X"53515357",
X"57547574",
X"24833875",
X"55748480",
X"8029fc80",
X"80057090",
X"2c515574",
X"ff2e9438",
X"83c8d008",
X"81801133",
X"5154737c",
X"7081055e",
X"34db3977",
X"22760554",
X"73782379",
X"09709f2a",
X"70810682",
X"1c3381bf",
X"0671862b",
X"07515151",
X"5473821a",
X"347c7626",
X"8a387722",
X"547a7426",
X"febb3880",
X"547383c0",
X"800c8f3d",
X"0d04f93d",
X"0d7a5780",
X"0b893d23",
X"893dfc05",
X"53765279",
X"51f8da3f",
X"83c08008",
X"81ff0670",
X"57557496",
X"387c547b",
X"53883d22",
X"527651fd",
X"e53f83c0",
X"800881ff",
X"06567583",
X"c0800c89",
X"3d0d04f0",
X"3d0d6266",
X"02880580",
X"ce052241",
X"5d5e8002",
X"840580d2",
X"05227f81",
X"0533ff11",
X"5a5d5a5d",
X"81da5876",
X"bf2680e9",
X"3878802e",
X"80e1387a",
X"58787b27",
X"83387858",
X"821e3370",
X"872a585a",
X"76923d34",
X"923dfc05",
X"5677557b",
X"547e537d",
X"33528251",
X"f8de3f83",
X"c0800881",
X"ff065d80",
X"0b923d33",
X"585a7680",
X"2e833881",
X"5a821e33",
X"80ff067a",
X"872b0757",
X"76821f34",
X"7c913878",
X"78317083",
X"ffff0679",
X"1e5e5a57",
X"ff9b397c",
X"587783c0",
X"800c923d",
X"0d04f83d",
X"0d7b0284",
X"05b20522",
X"5858800b",
X"8a3d238a",
X"3dfc0553",
X"77527a51",
X"f6f73f83",
X"c0800881",
X"ff067057",
X"55749638",
X"7d547653",
X"893d2252",
X"7751feaf",
X"3f83c080",
X"0881ff06",
X"567583c0",
X"800c8a3d",
X"0d04ec3d",
X"0d666e02",
X"880580df",
X"0533028c",
X"0580e305",
X"33029005",
X"80e70533",
X"02940580",
X"eb053302",
X"980580ee",
X"05224143",
X"415f5c40",
X"570280f2",
X"0522963d",
X"23963df0",
X"05538417",
X"70537752",
X"59f6863f",
X"83c08008",
X"81ff0658",
X"7781e538",
X"777a8180",
X"06584080",
X"77258338",
X"81407994",
X"3d347b02",
X"840580c9",
X"05347c02",
X"840580ca",
X"05347d02",
X"840580cb",
X"05347a95",
X"3d347a88",
X"2a577602",
X"840580cd",
X"0534953d",
X"22577602",
X"840580ce",
X"05347688",
X"2a577602",
X"840580cf",
X"05347792",
X"3d34963d",
X"ec115757",
X"8855f417",
X"54923d22",
X"53775277",
X"51f6953f",
X"83c08008",
X"81ff0658",
X"7780ed38",
X"7e802e80",
X"cb38923d",
X"22790858",
X"587f802e",
X"9c387681",
X"80800779",
X"0c7e5496",
X"3dfc0553",
X"7783ffff",
X"06527851",
X"f9fc3f99",
X"39768280",
X"8007790c",
X"7e54953d",
X"22537783",
X"ffff0652",
X"7851fc8f",
X"3f83c080",
X"0881ff06",
X"58779d38",
X"923d2253",
X"80527f30",
X"70802584",
X"71315351",
X"57f9873f",
X"83c08008",
X"81ff0658",
X"7783c080",
X"0c963d0d",
X"04f63d0d",
X"7c028405",
X"b705335b",
X"5b805880",
X"57805680",
X"55795485",
X"5380527a",
X"51fda33f",
X"83c08008",
X"81ff0659",
X"78853879",
X"871c3478",
X"83c0800c",
X"8c3d0d04",
X"f93d0d02",
X"a7053302",
X"8405ab05",
X"33028805",
X"af053358",
X"5957800b",
X"83c8df33",
X"54547274",
X"2e9f3881",
X"147081ff",
X"06555373",
X"872681b6",
X"387381c4",
X"2983c8dc",
X"05831133",
X"515372e3",
X"387381c4",
X"2983c8d8",
X"0555800b",
X"87163476",
X"88163475",
X"8a163477",
X"89163480",
X"750c83c8",
X"d0088c16",
X"0c800b84",
X"1634880b",
X"85163480",
X"0b861634",
X"841508ff",
X"a1ff06a0",
X"80078416",
X"0c811470",
X"81ff0653",
X"537451fe",
X"bc3f83c0",
X"800881ff",
X"06705553",
X"7280cd38",
X"8a397308",
X"750c7254",
X"80c23972",
X"81eaa455",
X"5681eaa4",
X"08802eb2",
X"38758429",
X"14700876",
X"53700851",
X"5454722d",
X"83c08008",
X"81ff0653",
X"72802ece",
X"38811670",
X"81ff0681",
X"eaa47184",
X"29115356",
X"57537208",
X"d0388054",
X"7383c080",
X"0c893d0d",
X"04f93d0d",
X"7957800b",
X"84180883",
X"c8d00c58",
X"f08c3f88",
X"170883c0",
X"80082783",
X"ed38effe",
X"3f83c080",
X"08810588",
X"180c83c8",
X"d008b811",
X"337081ff",
X"06515154",
X"73812ea4",
X"38738124",
X"88387378",
X"2e8a38b8",
X"3973822e",
X"9538b139",
X"763381f0",
X"06547390",
X"2ea63891",
X"7734a139",
X"73587633",
X"81f00654",
X"73902e09",
X"81069138",
X"efac3f83",
X"c0800881",
X"c8058c18",
X"0ca07734",
X"80567581",
X"c42983c8",
X"df113355",
X"5573802e",
X"aa3883c8",
X"d8157008",
X"56547480",
X"2e9d3888",
X"1508802e",
X"96388c14",
X"0883c8d0",
X"082e0981",
X"06893873",
X"51881508",
X"54732d81",
X"167081ff",
X"06575487",
X"7627ffba",
X"38763354",
X"73b02e81",
X"993873b0",
X"248f3873",
X"912eab38",
X"73a02e80",
X"f53882a6",
X"397380d0",
X"2e81e438",
X"7380d024",
X"8b387380",
X"c02e8199",
X"38828f39",
X"7381802e",
X"81fb3882",
X"85398056",
X"7581c429",
X"83c8dc11",
X"83113356",
X"59557380",
X"2ea83883",
X"c8d81570",
X"08565474",
X"802e9b38",
X"8c140883",
X"c8d0082e",
X"0981068e",
X"38735184",
X"15085473",
X"2d800b83",
X"19348116",
X"7081ff06",
X"57548776",
X"27ffb938",
X"92773481",
X"b539edc6",
X"3f8c1708",
X"83c08008",
X"2781a738",
X"b0773481",
X"a13983c8",
X"d0085480",
X"0b8c1534",
X"83c8d008",
X"54840b88",
X"153480c0",
X"7734ed9a",
X"3f83c080",
X"08b2058c",
X"180c80fa",
X"39ed8b3f",
X"8c170883",
X"c0800827",
X"80ec3883",
X"c8d00854",
X"810b8c15",
X"3483c8d0",
X"0854800b",
X"88153483",
X"c8d00854",
X"880ba015",
X"34ecdf3f",
X"83c08008",
X"94058c18",
X"0c80d077",
X"34bc3983",
X"c8d008a0",
X"11337083",
X"2a708106",
X"51515555",
X"73802ea6",
X"38880ba0",
X"1634ecb2",
X"3f8c1708",
X"83c08008",
X"279438ff",
X"8077348e",
X"39775380",
X"528051fa",
X"8b3fff90",
X"773483c8",
X"d008a011",
X"3370832a",
X"70810651",
X"51555573",
X"802e8638",
X"880ba016",
X"34893d0d",
X"04f43d0d",
X"02bb0533",
X"028405bf",
X"05335d5d",
X"800b83c8",
X"dc0b83c8",
X"d80b8c11",
X"72718814",
X"755c5a5b",
X"5f5c595b",
X"58831533",
X"5372802e",
X"81883873",
X"33537c73",
X"2e098106",
X"80fc3881",
X"1433537b",
X"732e0981",
X"0680ef38",
X"750883c8",
X"d0082e09",
X"810680e2",
X"38805675",
X"81c42983",
X"c8e01170",
X"33831e33",
X"5b575553",
X"74782e09",
X"81069738",
X"83c8e413",
X"0879082e",
X"0981068a",
X"38811433",
X"527451fe",
X"f83f8116",
X"7081ff06",
X"57538776",
X"27c53880",
X"77085454",
X"72742e91",
X"38765184",
X"13085372",
X"2d83c080",
X"0881ff06",
X"54800b83",
X"1b347353",
X"a9398118",
X"81c41681",
X"c41681c4",
X"1981c41f",
X"81c41e81",
X"c41d6081",
X"c405415d",
X"5e5f5956",
X"56588778",
X"25feca38",
X"80537283",
X"c0800c8e",
X"3d0d04f8",
X"3d0d02ae",
X"05227d59",
X"57805681",
X"55805486",
X"53818052",
X"7a51f4ee",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8a3d0d04",
X"f73d0d02",
X"b2052202",
X"8405b705",
X"33605a5b",
X"57805682",
X"55795486",
X"53818052",
X"7b51f4be",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8b3d0d04",
X"f83d0d02",
X"af053359",
X"80588057",
X"80568055",
X"78548953",
X"80527a51",
X"f4943f83",
X"c0800881",
X"ff0683c0",
X"800c8a3d",
X"0d04ffb8",
X"3d0d80cb",
X"3d087053",
X"81e8f052",
X"56febeb6",
X"3f83c080",
X"0880f338",
X"7551feb8",
X"a13f83ff",
X"ff0b83c0",
X"80082580",
X"e1387551",
X"feb8a03f",
X"83c08008",
X"5583c080",
X"0880cf38",
X"82805383",
X"c0800852",
X"8a3d7052",
X"57fefbd9",
X"3f745275",
X"51feb790",
X"3f805980",
X"ca3dfdfc",
X"05548280",
X"53765275",
X"51feb596",
X"3f811555",
X"7488802e",
X"098106e1",
X"38805275",
X"51feb6e8",
X"3f800b83",
X"d4fc0c75",
X"83d4f80c",
X"8739800b",
X"83d4f80c",
X"80ca3d0d",
X"04ff3d0d",
X"73700853",
X"51029305",
X"33723470",
X"08810571",
X"0c833d0d",
X"04ffb83d",
X"0d80cb3d",
X"70708405",
X"52085856",
X"83d4f808",
X"802e80fa",
X"388a3d70",
X"5a765577",
X"5481d6a1",
X"5380cb3d",
X"fdfc0552",
X"55fee3b4",
X"3f805280",
X"ca3dfdfc",
X"0551ffad",
X"3f83d4fc",
X"085283d4",
X"f80851fe",
X"b5ee3f80",
X"587451fe",
X"e0f63f80",
X"ca3dfdf8",
X"055483c0",
X"80085374",
X"5283d4f8",
X"0851feb3",
X"e93f83d4",
X"fc081883",
X"d4fc0c80",
X"ca3dfdf8",
X"05548153",
X"81e8fc52",
X"83d4f808",
X"51feb3ca",
X"3f83d4fc",
X"081883d4",
X"fc0c80ca",
X"3d0d0483",
X"c08c0802",
X"83c08c0c",
X"fd3d0d80",
X"5383c08c",
X"088c0508",
X"5283c08c",
X"08880508",
X"5183d43f",
X"83c08008",
X"7083c080",
X"0c54853d",
X"0d83c08c",
X"0c0483c0",
X"8c080283",
X"c08c0cfd",
X"3d0d8153",
X"83c08c08",
X"8c050852",
X"83c08c08",
X"88050851",
X"83a13f83",
X"c0800870",
X"83c0800c",
X"54853d0d",
X"83c08c0c",
X"0483c08c",
X"080283c0",
X"8c0cf93d",
X"0d800b83",
X"c08c08fc",
X"050c83c0",
X"8c088805",
X"088025b9",
X"3883c08c",
X"08880508",
X"3083c08c",
X"0888050c",
X"800b83c0",
X"8c08f405",
X"0c83c08c",
X"08fc0508",
X"8a38810b",
X"83c08c08",
X"f4050c83",
X"c08c08f4",
X"050883c0",
X"8c08fc05",
X"0c83c08c",
X"088c0508",
X"8025b938",
X"83c08c08",
X"8c050830",
X"83c08c08",
X"8c050c80",
X"0b83c08c",
X"08f0050c",
X"83c08c08",
X"fc05088a",
X"38810b83",
X"c08c08f0",
X"050c83c0",
X"8c08f005",
X"0883c08c",
X"08fc050c",
X"805383c0",
X"8c088c05",
X"085283c0",
X"8c088805",
X"085181df",
X"3f83c080",
X"087083c0",
X"8c08f805",
X"0c5483c0",
X"8c08fc05",
X"08802e90",
X"3883c08c",
X"08f80508",
X"3083c08c",
X"08f8050c",
X"83c08c08",
X"f8050870",
X"83c0800c",
X"54893d0d",
X"83c08c0c",
X"0483c08c",
X"080283c0",
X"8c0cfb3d",
X"0d800b83",
X"c08c08fc",
X"050c83c0",
X"8c088805",
X"08802599",
X"3883c08c",
X"08880508",
X"3083c08c",
X"0888050c",
X"810b83c0",
X"8c08fc05",
X"0c83c08c",
X"088c0508",
X"80259038",
X"83c08c08",
X"8c050830",
X"83c08c08",
X"8c050c81",
X"5383c08c",
X"088c0508",
X"5283c08c",
X"08880508",
X"51bd3f83",
X"c0800870",
X"83c08c08",
X"f8050c54",
X"83c08c08",
X"fc050880",
X"2e903883",
X"c08c08f8",
X"05083083",
X"c08c08f8",
X"050c83c0",
X"8c08f805",
X"087083c0",
X"800c5487",
X"3d0d83c0",
X"8c0c0483",
X"c08c0802",
X"83c08c0c",
X"fd3d0d81",
X"0b83c08c",
X"08fc050c",
X"800b83c0",
X"8c08f805",
X"0c83c08c",
X"088c0508",
X"83c08c08",
X"88050827",
X"b93883c0",
X"8c08fc05",
X"08802eae",
X"38800b83",
X"c08c088c",
X"050824a2",
X"3883c08c",
X"088c0508",
X"1083c08c",
X"088c050c",
X"83c08c08",
X"fc050810",
X"83c08c08",
X"fc050cff",
X"b83983c0",
X"8c08fc05",
X"08802e80",
X"e13883c0",
X"8c088c05",
X"0883c08c",
X"08880508",
X"26ad3883",
X"c08c0888",
X"050883c0",
X"8c088c05",
X"083183c0",
X"8c088805",
X"0c83c08c",
X"08f80508",
X"83c08c08",
X"fc050807",
X"83c08c08",
X"f8050c83",
X"c08c08fc",
X"0508812a",
X"83c08c08",
X"fc050c83",
X"c08c088c",
X"0508812a",
X"83c08c08",
X"8c050cff",
X"953983c0",
X"8c089005",
X"08802e93",
X"3883c08c",
X"08880508",
X"7083c08c",
X"08f4050c",
X"51913983",
X"c08c08f8",
X"05087083",
X"c08c08f4",
X"050c5183",
X"c08c08f4",
X"050883c0",
X"800c853d",
X"0d83c08c",
X"0c0483c0",
X"8c080283",
X"c08c0cff",
X"3d0d800b",
X"83c08c08",
X"fc050c83",
X"c08c0888",
X"05088106",
X"ff117009",
X"7083c08c",
X"088c0508",
X"0683c08c",
X"08fc0508",
X"1183c08c",
X"08fc050c",
X"83c08c08",
X"88050881",
X"2a83c08c",
X"0888050c",
X"83c08c08",
X"8c050810",
X"83c08c08",
X"8c050c51",
X"51515183",
X"c08c0888",
X"0508802e",
X"8438ffab",
X"3983c08c",
X"08fc0508",
X"7083c080",
X"0c51833d",
X"0d83c08c",
X"0c04fc3d",
X"0d767079",
X"7b555555",
X"558f7227",
X"8c387275",
X"07830651",
X"70802ea9",
X"38ff1252",
X"71ff2e98",
X"38727081",
X"05543374",
X"70810556",
X"34ff1252",
X"71ff2e09",
X"8106ea38",
X"7483c080",
X"0c863d0d",
X"04745172",
X"70840554",
X"08717084",
X"05530c72",
X"70840554",
X"08717084",
X"05530c72",
X"70840554",
X"08717084",
X"05530c72",
X"70840554",
X"08717084",
X"05530cf0",
X"1252718f",
X"26c93883",
X"72279538",
X"72708405",
X"54087170",
X"8405530c",
X"fc125271",
X"8326ed38",
X"7054ff81",
X"39000000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"70704740",
X"0c704268",
X"0c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"000031fa",
X"0000323b",
X"0000325b",
X"0000327f",
X"0000328b",
X"00003295",
X"00003e8e",
X"00004831",
X"000048fa",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3a00",
X"0c0c3b00",
X"0a0a0005",
X"0b0b0005",
X"06060005",
X"07070004",
X"04044500",
X"05054400",
X"0e0f2900",
X"08080004",
X"09090004",
X"0a0f4300",
X"090f4200",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"02010302",
X"02020204",
X"01020800",
X"03800403",
X"20050310",
X"06034007",
X"03010803",
X"02090480",
X"0a05800b",
X"02200c02",
X"100d0240",
X"0e02800f",
X"000057b9",
X"00005ac0",
X"000058cc",
X"00005ac0",
X"00005909",
X"0000595a",
X"00005999",
X"000059a2",
X"00005ac0",
X"00005ac0",
X"00005ac0",
X"00005ac0",
X"000059ab",
X"000059b3",
X"000059ba",
X"00005bc0",
X"00005cb9",
X"00005dcd",
X"000060bf",
X"000060da",
X"000060c6",
X"000060da",
X"000060e1",
X"000060ec",
X"000060f3",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"41545800",
X"63686f6f",
X"73652000",
X"66696c65",
X"20202573",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"25782e48",
X"75622e20",
X"25642070",
X"6f727473",
X"00000000",
X"25782e48",
X"49440000",
X"204d6f75",
X"73650000",
X"204b6579",
X"626f6172",
X"64000000",
X"204a6f79",
X"73746963",
X"6b3a2564",
X"00000000",
X"52474200",
X"5343414e",
X"444f5542",
X"4c450000",
X"53564944",
X"454f0000",
X"48444d49",
X"00000000",
X"44564900",
X"56474100",
X"434f4d50",
X"4f534954",
X"45000000",
X"4e545343",
X"00000000",
X"50414c00",
X"73657474",
X"696e6773",
X"00000000",
X"35323030",
X"2e726f6d",
X"00000000",
X"31364b00",
X"556e6b6e",
X"6f776e20",
X"74797065",
X"206f6620",
X"63617274",
X"72696467",
X"65210000",
X"41353200",
X"43415200",
X"42494e00",
X"31366b20",
X"63617274",
X"20747970",
X"65000000",
X"4c656674",
X"20666f72",
X"206f6e65",
X"20636869",
X"70000000",
X"52696768",
X"7420666f",
X"72207477",
X"6f206368",
X"69700000",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a257300",
X"526f7461",
X"74652055",
X"5342206a",
X"6f797374",
X"69636b73",
X"00000000",
X"45786974",
X"00000000",
X"524f4d00",
X"4d454d00",
X"52504400",
X"2f757362",
X"2e6c6f67",
X"00000000",
X"0a000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"00000000",
X"00007350",
X"00007354",
X"00007360",
X"00007368",
X"00007370",
X"00007374",
X"00007378",
X"00007384",
X"0000738c",
X"000072a0",
X"000070c0",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"35323030",
X"00000000",
X"2f617461",
X"72353230",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
