
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f0",
X"b8738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80f3",
X"f00c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580ef",
X"fa2d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580efb9",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80d98f04",
X"f93d0d80",
X"0b83e080",
X"0c893d0d",
X"04fc3d0d",
X"76705255",
X"b3933f83",
X"e0800815",
X"ff055473",
X"752e8e38",
X"73335372",
X"ae2e8638",
X"ff1454ef",
X"39775281",
X"1451b2ab",
X"3f83e080",
X"08307083",
X"e0800807",
X"802583e0",
X"800c5386",
X"3d0d04fc",
X"3d0d7670",
X"525599cc",
X"3f83e080",
X"08548153",
X"83e08008",
X"80c73874",
X"51998f3f",
X"83e08008",
X"0b0b80f1",
X"f85383e0",
X"80085253",
X"ff8f3f83",
X"e08008a5",
X"380b0b80",
X"f1fc5272",
X"51fefe3f",
X"83e08008",
X"94380b0b",
X"80f28052",
X"7251feed",
X"3f83e080",
X"08802e83",
X"38815473",
X"537283e0",
X"800c863d",
X"0d04fd3d",
X"0d757052",
X"5498e53f",
X"815383e0",
X"80089838",
X"735198ae",
X"3f83e0a0",
X"085283e0",
X"800851fe",
X"b43f83e0",
X"80085372",
X"83e0800c",
X"853d0d04",
X"e03d0da3",
X"3d087052",
X"5e8ed33f",
X"83e08008",
X"33943d56",
X"54739438",
X"80f6f452",
X"745184c7",
X"397d5278",
X"5191d63f",
X"84d1397d",
X"518ebb3f",
X"83e08008",
X"5274518d",
X"eb3f83e0",
X"a8085293",
X"3d70525d",
X"94c63f83",
X"e0800859",
X"800b83e0",
X"8008555b",
X"83e08008",
X"7b2e9438",
X"811b7452",
X"5b97c83f",
X"83e08008",
X"5483e080",
X"08ee3880",
X"5aff7a43",
X"7a427a41",
X"5f790970",
X"9f2c7b06",
X"5b547a7a",
X"248438ff",
X"1b5af61a",
X"7009709f",
X"2c72067b",
X"ff125a5a",
X"52555580",
X"75259538",
X"76519787",
X"3f83e080",
X"0876ff18",
X"58555773",
X"8024ed38",
X"747f2e87",
X"3880c299",
X"3f745f78",
X"ff1b7058",
X"5d58807a",
X"25953877",
X"5196dc3f",
X"83e08008",
X"76ff1858",
X"55587380",
X"24ed3880",
X"0b83e7bc",
X"0c800b83",
X"e7dc0c0b",
X"0b80f284",
X"518bae3f",
X"81800b83",
X"e7dc0c0b",
X"0b80f28c",
X"518b9e3f",
X"a80b83e7",
X"bc0c7680",
X"2e80e838",
X"83e7bc08",
X"77793270",
X"30707207",
X"80257087",
X"2b83e7dc",
X"0c515678",
X"53565696",
X"8f3f83e0",
X"8008802e",
X"8a380b0b",
X"80f29451",
X"8ae33f76",
X"5195cf3f",
X"83e08008",
X"520b0b80",
X"f3a0518a",
X"d03f7651",
X"95d53f83",
X"e0800883",
X"e7bc0855",
X"57757425",
X"8638a816",
X"56f73975",
X"83e7bc0c",
X"86f07624",
X"ff943887",
X"980b83e7",
X"bc0c7780",
X"2eb73877",
X"51958b3f",
X"83e08008",
X"78525595",
X"ab3f0b0b",
X"80f29c54",
X"83e08008",
X"8f388739",
X"807634fd",
X"95390b0b",
X"80f29854",
X"74537352",
X"0b0b80f1",
X"ec5189e9",
X"3f80540b",
X"0b80f3ec",
X"5189de3f",
X"81145473",
X"a82e0981",
X"06ed3886",
X"8da051be",
X"9b3f8052",
X"903d7052",
X"5480def6",
X"3f835273",
X"5180deee",
X"3f61802e",
X"80ff387b",
X"5473ff2e",
X"96387880",
X"2e818038",
X"785194ab",
X"3f83e080",
X"08ff1555",
X"59e73978",
X"802e80eb",
X"38785194",
X"a73f83e0",
X"8008802e",
X"fc833878",
X"5193ef3f",
X"83e08008",
X"520b0b80",
X"f1f451ab",
X"cd3f83e0",
X"8008a438",
X"7c51ad85",
X"3f83e080",
X"085574ff",
X"16565480",
X"7425fbee",
X"38741d70",
X"33555673",
X"af2efec8",
X"38e83978",
X"5193ad3f",
X"83e08008",
X"527c51ac",
X"bc3ffbce",
X"397f8829",
X"6010057a",
X"0561055a",
X"fbff39a2",
X"3d0d0480",
X"3d0d9080",
X"f8337081",
X"ff067084",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d38a8",
X"0b9080f8",
X"34b80b90",
X"80f83470",
X"83e0800c",
X"823d0d04",
X"803d0d90",
X"80f83370",
X"81ff0670",
X"852a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"980b9080",
X"f834b80b",
X"9080f834",
X"7083e080",
X"0c823d0d",
X"04930b90",
X"80fc34ff",
X"0b9080e8",
X"3404ff3d",
X"0d028f05",
X"3352800b",
X"9080fc34",
X"8a51bbf0",
X"3fdf3f80",
X"f80b9080",
X"e034800b",
X"9080c834",
X"fa125271",
X"9080c034",
X"800b9080",
X"d8347190",
X"80d03490",
X"80f85280",
X"7234b872",
X"34833d0d",
X"04803d0d",
X"028b0533",
X"51709080",
X"f434febf",
X"3f83e080",
X"08802ef6",
X"38823d0d",
X"04803d0d",
X"853980c5",
X"ac3ffed8",
X"3f83e080",
X"08802ef2",
X"389080f4",
X"337081ff",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0da30b90",
X"80fc34ff",
X"0b9080e8",
X"349080f8",
X"51a87134",
X"b8713482",
X"3d0d0480",
X"3d0d9080",
X"fc337081",
X"c0067030",
X"70802583",
X"e0800c51",
X"5151823d",
X"0d04803d",
X"0d9080f8",
X"337081ff",
X"0670832a",
X"81327081",
X"06515151",
X"5170802e",
X"e838b00b",
X"9080f834",
X"b80b9080",
X"f834823d",
X"0d04803d",
X"0d9080ac",
X"08810683",
X"e0800c82",
X"3d0d04fd",
X"3d0d7577",
X"54548073",
X"25943873",
X"70810555",
X"335280f2",
X"a05185a1",
X"3fff1353",
X"e939853d",
X"0d04f63d",
X"0d7c7e60",
X"625a5d5b",
X"56805981",
X"55853974",
X"7a295574",
X"52755180",
X"dbd73f83",
X"e080087a",
X"27ed3874",
X"802e80e0",
X"38745275",
X"5180dbc1",
X"3f83e080",
X"08755376",
X"525480db",
X"c43f83e0",
X"80087a53",
X"75525680",
X"dba73f83",
X"e0800879",
X"30707b07",
X"9f2a7077",
X"80240751",
X"51545572",
X"873883e0",
X"8008c238",
X"768118b0",
X"16555858",
X"8974258b",
X"38b71453",
X"7a853880",
X"d7145372",
X"78348119",
X"59ff9c39",
X"8077348c",
X"3d0d04f7",
X"3d0d7b7d",
X"7f620290",
X"05bb0533",
X"5759565a",
X"5ab05872",
X"8338a058",
X"75707081",
X"05523371",
X"59545590",
X"39807425",
X"8e38ff14",
X"77708105",
X"59335454",
X"72ef3873",
X"ff155553",
X"80732589",
X"38775279",
X"51782def",
X"39753375",
X"57537280",
X"2e903872",
X"52795178",
X"2d757081",
X"05573353",
X"ed398b3d",
X"0d04ee3d",
X"0d646669",
X"69707081",
X"0552335b",
X"4a5c5e5e",
X"76802e82",
X"f93876a5",
X"2e098106",
X"82e03880",
X"70416770",
X"70810552",
X"33714a59",
X"575f76b0",
X"2e098106",
X"8c387570",
X"81055733",
X"76485781",
X"5fd01756",
X"75892680",
X"da387667",
X"5c59805c",
X"9339778a",
X"2480c338",
X"7b8a2918",
X"7b708105",
X"5d335a5c",
X"d0197081",
X"ff065858",
X"897727a4",
X"38ff9f19",
X"7081ff06",
X"ffa91b5a",
X"51568576",
X"279238ff",
X"bf197081",
X"ff065156",
X"7585268a",
X"38c91958",
X"778025ff",
X"b9387a47",
X"7b407881",
X"ff065776",
X"80e42e80",
X"e5387680",
X"e424a738",
X"7680d82e",
X"81863876",
X"80d82490",
X"3876802e",
X"81cc3876",
X"a52e81b6",
X"3881b939",
X"7680e32e",
X"818c3881",
X"af397680",
X"f52e9b38",
X"7680f524",
X"8b387680",
X"f32e8181",
X"38819939",
X"7680f82e",
X"80ca3881",
X"8f39913d",
X"70555780",
X"538a5279",
X"841b7108",
X"535b56fb",
X"fd3f7655",
X"ab397984",
X"1b710894",
X"3d705b5b",
X"525b5675",
X"80258c38",
X"753056ad",
X"78340280",
X"c1055776",
X"5480538a",
X"527551fb",
X"d13f7755",
X"7e54b839",
X"913d7055",
X"7780d832",
X"70307080",
X"25565158",
X"56905279",
X"841b7108",
X"535b57fb",
X"ad3f7555",
X"db397984",
X"1b831233",
X"545b5698",
X"3979841b",
X"7108575b",
X"5680547f",
X"537c527d",
X"51fc9c3f",
X"87397652",
X"7d517c2d",
X"66703358",
X"810547fd",
X"8339943d",
X"0d047283",
X"e0900c71",
X"83e0940c",
X"04fb3d0d",
X"883d7070",
X"84055208",
X"57547553",
X"83e09008",
X"5283e094",
X"0851fcc6",
X"3f873d0d",
X"04ff3d0d",
X"73700853",
X"51029305",
X"33723470",
X"08810571",
X"0c833d0d",
X"04fc3d0d",
X"873d8811",
X"55785498",
X"dd5351fc",
X"993f8052",
X"873d51d1",
X"3f863d0d",
X"04fd3d0d",
X"75705254",
X"a3c33f83",
X"e0800814",
X"5372742e",
X"9238ff13",
X"70335353",
X"71af2e09",
X"8106ee38",
X"81135372",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"77705354",
X"54c73f83",
X"e0800873",
X"2ea13883",
X"e0800873",
X"3152ff12",
X"5271ff2e",
X"8f387270",
X"81055433",
X"74708105",
X"5634eb39",
X"ff145480",
X"7434853d",
X"0d04803d",
X"0d7251ff",
X"903f823d",
X"0d047183",
X"e0800c04",
X"803d0d72",
X"51807134",
X"810bbc12",
X"0c800b80",
X"c0120c82",
X"3d0d0480",
X"0b83e2d4",
X"08248a38",
X"a4ad3fff",
X"0b83e2d4",
X"0c800b83",
X"e0800c04",
X"ff3d0d73",
X"5283e0b0",
X"08722e8d",
X"38d93f71",
X"5196983f",
X"7183e0b0",
X"0c833d0d",
X"04f43d0d",
X"7e60625c",
X"5a558154",
X"bc150881",
X"91387451",
X"cf3f7958",
X"807a2580",
X"f73883e3",
X"84087089",
X"2a5783ff",
X"06788480",
X"72315656",
X"57737825",
X"83387355",
X"7583e2d4",
X"082e8438",
X"ff893f83",
X"e2d40880",
X"25a63875",
X"892b5198",
X"db3f83e3",
X"84088f3d",
X"fc11555c",
X"548152f8",
X"1b5196c5",
X"3f761483",
X"e3840c75",
X"83e2d40c",
X"74537652",
X"7851a2de",
X"3f83e080",
X"0883e384",
X"081683e3",
X"840c7876",
X"31761b5b",
X"59567780",
X"24ff8b38",
X"617a710c",
X"54755475",
X"802e8338",
X"81547383",
X"e0800c8e",
X"3d0d04fc",
X"3d0dfe9b",
X"3f7651fe",
X"af3f863d",
X"fc055378",
X"52775195",
X"e83f7975",
X"710c5483",
X"e0800854",
X"83e08008",
X"802e8338",
X"81547383",
X"e0800c86",
X"3d0d04fe",
X"3d0d7583",
X"e2d40853",
X"53807224",
X"89387173",
X"2e8438fd",
X"d63f7451",
X"fdea3f72",
X"5197ad3f",
X"83e08008",
X"5283e080",
X"08802e83",
X"38815271",
X"83e0800c",
X"843d0d04",
X"803d0d72",
X"80c01108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"72bc1108",
X"83e0800c",
X"51823d0d",
X"0480c40b",
X"83e0800c",
X"04fd3d0d",
X"75777154",
X"70535553",
X"9f9b3f82",
X"c81308bc",
X"150c82c0",
X"130880c0",
X"150cfceb",
X"3f735193",
X"aa3f7383",
X"e0b00c83",
X"e0800853",
X"83e08008",
X"802e8338",
X"81537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"5553fcbf",
X"3f72802e",
X"a538bc13",
X"08527351",
X"9ea53f83",
X"e080088f",
X"38775272",
X"51ff9a3f",
X"83e08008",
X"538a3982",
X"cc130853",
X"d8398153",
X"7283e080",
X"0c853d0d",
X"04fe3d0d",
X"ff0b83e2",
X"d40c7483",
X"e0b40c75",
X"83e2d00c",
X"9f923f83",
X"e0800881",
X"ff065281",
X"53719938",
X"83e2ec51",
X"8e943f83",
X"e0800852",
X"83e08008",
X"802e8338",
X"72527153",
X"7283e080",
X"0c843d0d",
X"04fa3d0d",
X"787a82c4",
X"120882c4",
X"12087072",
X"24595656",
X"57577373",
X"2e098106",
X"913880c0",
X"165280c0",
X"17519c96",
X"3f83e080",
X"08557483",
X"e0800c88",
X"3d0d04f6",
X"3d0d7c5b",
X"807b715c",
X"54577a77",
X"2e8c3881",
X"1a82cc14",
X"08545a72",
X"f6388059",
X"80d9397a",
X"54815780",
X"707b7b31",
X"5a5755ff",
X"18537473",
X"2580c138",
X"82cc1408",
X"527351ff",
X"8c3f800b",
X"83e08008",
X"25a13882",
X"cc140882",
X"cc110882",
X"cc160c74",
X"82cc120c",
X"5375802e",
X"86387282",
X"cc170c72",
X"54805773",
X"82cc1508",
X"81175755",
X"56ffb839",
X"81195980",
X"0bff1b54",
X"54787325",
X"83388154",
X"76813270",
X"75065153",
X"72ff9038",
X"8c3d0d04",
X"f73d0d7b",
X"7d5a5a82",
X"d05283e2",
X"d0085180",
X"cedf3f83",
X"e0800857",
X"f9e13f79",
X"5283e2d8",
X"5195b43f",
X"83e08008",
X"54805383",
X"e0800873",
X"2e098106",
X"82833883",
X"e0b4080b",
X"0b80f1f4",
X"53705256",
X"9bd33f0b",
X"0b80f1f4",
X"5280c016",
X"519bc63f",
X"75bc170c",
X"7382c017",
X"0c810b82",
X"c4170c81",
X"0b82c817",
X"0c7382cc",
X"170cff17",
X"82d01755",
X"57819139",
X"83e0c033",
X"70822a70",
X"81065154",
X"55728180",
X"3874812a",
X"81065877",
X"80f63874",
X"842a8106",
X"82c4150c",
X"83e0c033",
X"810682c8",
X"150c7952",
X"73519aed",
X"3f73519b",
X"843f83e0",
X"80081453",
X"af737081",
X"05553472",
X"bc150c83",
X"e0c15272",
X"519ace3f",
X"83e0b808",
X"82c0150c",
X"83e0ce52",
X"80c01451",
X"9abb3f78",
X"802e8d38",
X"7351782d",
X"83e08008",
X"802e9938",
X"7782cc15",
X"0c75802e",
X"86387382",
X"cc170c73",
X"82d015ff",
X"19595556",
X"76802e9b",
X"3883e0b8",
X"5283e2d8",
X"5194aa3f",
X"83e08008",
X"8a3883e0",
X"c1335372",
X"fed23878",
X"802e8938",
X"83e0b408",
X"51fcb83f",
X"83e0b408",
X"537283e0",
X"800c8b3d",
X"0d04ff3d",
X"0d805273",
X"51fdb53f",
X"833d0d04",
X"f03d0d62",
X"705254f6",
X"903f83e0",
X"80087453",
X"873d7053",
X"5555f6b0",
X"3ff7903f",
X"7351d33f",
X"63537452",
X"83e08008",
X"51fab83f",
X"923d0d04",
X"7183e080",
X"0c0480c0",
X"1283e080",
X"0c04803d",
X"0d7282c0",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"cc110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"82c41108",
X"83e0800c",
X"51823d0d",
X"04f93d0d",
X"7983e098",
X"08575781",
X"77278196",
X"38768817",
X"0827818e",
X"38753355",
X"74822e89",
X"3874832e",
X"b33880fe",
X"39745476",
X"1083fe06",
X"5376882a",
X"8c170805",
X"52893dfc",
X"055199c0",
X"3f83e080",
X"0880df38",
X"029d0533",
X"893d3371",
X"882b0756",
X"5680d139",
X"84547682",
X"2b83fc06",
X"5376872a",
X"8c170805",
X"52893dfc",
X"05519990",
X"3f83e080",
X"08b03802",
X"9f053302",
X"84059e05",
X"3371982b",
X"71902b07",
X"028c059d",
X"05337088",
X"2b72078d",
X"3d337180",
X"fffffe80",
X"06075152",
X"53575856",
X"83398155",
X"7483e080",
X"0c893d0d",
X"04fb3d0d",
X"83e09808",
X"fe198812",
X"08fe0555",
X"56548056",
X"7473278d",
X"38821433",
X"75712994",
X"16080557",
X"537583e0",
X"800c873d",
X"0d04fc3d",
X"0d765280",
X"0b83e098",
X"08703351",
X"52537083",
X"2e098106",
X"91389512",
X"33941333",
X"71982b71",
X"902b0755",
X"55519b12",
X"339a1333",
X"71882b07",
X"740783e0",
X"800c5586",
X"3d0d04fc",
X"3d0d7683",
X"e0980855",
X"55807523",
X"88150853",
X"72812e88",
X"38881408",
X"73268538",
X"8152b239",
X"72903873",
X"33527183",
X"2e098106",
X"85389014",
X"0853728c",
X"160c7280",
X"2e8d3872",
X"51fed63f",
X"83e08008",
X"52853990",
X"14085271",
X"90160c80",
X"527183e0",
X"800c863d",
X"0d04fa3d",
X"0d7883e0",
X"98087122",
X"81057083",
X"ffff0657",
X"54575573",
X"802e8838",
X"90150853",
X"72863883",
X"5280e739",
X"738f0652",
X"7180da38",
X"81139016",
X"0c8c1508",
X"53729038",
X"830b8417",
X"22575273",
X"762780c6",
X"38bf3982",
X"1633ff05",
X"74842a06",
X"5271b238",
X"7251fcb1",
X"3f815271",
X"83e08008",
X"27a83883",
X"5283e080",
X"08881708",
X"279c3883",
X"e080088c",
X"160c83e0",
X"800851fd",
X"bc3f83e0",
X"80089016",
X"0c737523",
X"80527183",
X"e0800c88",
X"3d0d04f2",
X"3d0d6062",
X"64585e5b",
X"75335574",
X"a02e0981",
X"06883881",
X"16704456",
X"ef396270",
X"33565674",
X"af2e0981",
X"06843881",
X"1643800b",
X"881c0c62",
X"70335155",
X"749f2691",
X"387a51fd",
X"d23f83e0",
X"80085680",
X"7d348381",
X"39933d84",
X"1c087058",
X"595f8a55",
X"a0767081",
X"055834ff",
X"155574ff",
X"2e098106",
X"ef388070",
X"5a5c887f",
X"085f5a7b",
X"811d7081",
X"ff066013",
X"703370af",
X"327030a0",
X"73277180",
X"25075151",
X"525b535e",
X"57557480",
X"e73876ae",
X"2e098106",
X"83388155",
X"787a2775",
X"07557480",
X"2e9f3879",
X"88327030",
X"78ae3270",
X"30707307",
X"9f2a5351",
X"57515675",
X"bb388859",
X"8b5affab",
X"3976982b",
X"55748025",
X"873880ef",
X"c8173357",
X"ff9f1755",
X"74992689",
X"38e01770",
X"81ff0658",
X"5578811a",
X"7081ff06",
X"721b535b",
X"57557675",
X"34fef839",
X"7b1e7f0c",
X"805576a0",
X"26833881",
X"55748b19",
X"347a51fc",
X"823f83e0",
X"800880f5",
X"38a0547a",
X"2270852b",
X"83e00654",
X"55901b08",
X"527c5193",
X"cb3f83e0",
X"80085783",
X"e0800881",
X"81387c33",
X"5574802e",
X"80f4388b",
X"1d337083",
X"2a708106",
X"51565674",
X"b4388b7d",
X"841d0883",
X"e0800859",
X"5b5b58ff",
X"185877ff",
X"2e9a3879",
X"7081055b",
X"33797081",
X"055b3371",
X"71315256",
X"5675802e",
X"e2388639",
X"75802e96",
X"387a51fb",
X"e53fff86",
X"3983e080",
X"085683e0",
X"8008b638",
X"83397656",
X"841b088b",
X"11335155",
X"74a7388b",
X"1d337084",
X"2a708106",
X"51565674",
X"89388356",
X"94398156",
X"90397c51",
X"fa943f83",
X"e0800888",
X"1c0cfd81",
X"397583e0",
X"800c903d",
X"0d04f83d",
X"0d7a7c59",
X"57825483",
X"fe537752",
X"76519290",
X"3f835683",
X"e0800880",
X"ec388117",
X"33773371",
X"882b0756",
X"56825674",
X"82d4d52e",
X"09810680",
X"d4387554",
X"b6537752",
X"765191e4",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"ac388254",
X"80d25377",
X"52765191",
X"bb3f83e0",
X"80089838",
X"81173377",
X"3371882b",
X"0783e080",
X"08525656",
X"748182c6",
X"2e833881",
X"567583e0",
X"800c8a3d",
X"0d04eb3d",
X"0d675a80",
X"0b83e098",
X"0c90dd3f",
X"83e08008",
X"81065582",
X"567483ee",
X"38747553",
X"8f3d7053",
X"5759feca",
X"3f83e080",
X"0881ff06",
X"5776812e",
X"09810680",
X"d4389054",
X"83be5374",
X"52755190",
X"cf3f83e0",
X"800880c9",
X"388f3d33",
X"5574802e",
X"80c93802",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"70587b57",
X"5e525e57",
X"5957fdee",
X"3f83e080",
X"0881ff06",
X"5776832e",
X"09810686",
X"38815682",
X"f1397680",
X"2e863886",
X"5682e739",
X"a4548d53",
X"78527551",
X"8fe63f81",
X"5683e080",
X"0882d338",
X"02be0533",
X"028405bd",
X"05337188",
X"2b07595d",
X"77ab3802",
X"80ce0533",
X"02840580",
X"cd053371",
X"982b7190",
X"2b07973d",
X"3370882b",
X"72070294",
X"0580cb05",
X"33710754",
X"525e5759",
X"5602b705",
X"33787129",
X"028805b6",
X"0533028c",
X"05b50533",
X"71882b07",
X"701d707f",
X"8c050c5f",
X"5957595d",
X"8e3d3382",
X"1b3402b9",
X"0533903d",
X"3371882b",
X"075a5c78",
X"841b2302",
X"bb053302",
X"8405ba05",
X"3371882b",
X"07565c74",
X"ab380280",
X"ca053302",
X"840580c9",
X"05337198",
X"2b71902b",
X"07963d33",
X"70882b72",
X"07029405",
X"80c70533",
X"71075152",
X"53575e5c",
X"74763178",
X"3179842a",
X"903d3354",
X"71713153",
X"5656bfc5",
X"3f83e080",
X"08820570",
X"881c0c83",
X"e08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83e0980c",
X"80567583",
X"e0800c97",
X"3d0d04e9",
X"3d0d83e0",
X"98085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e63f83e0",
X"80085483",
X"e0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f48a",
X"3f83e080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383e080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83e09808",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0ea3f",
X"83e08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"843f83e0",
X"80085583",
X"e0800880",
X"2eff8938",
X"83e08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"518a8d3f",
X"83e08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83e0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83e09808",
X"55568555",
X"73802e81",
X"e1388114",
X"33810653",
X"84557280",
X"2e81d338",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b7388214",
X"3370892b",
X"56537680",
X"2eb53874",
X"52ff1651",
X"bac73f83",
X"e08008ff",
X"18765470",
X"535853ba",
X"b83f83e0",
X"80087326",
X"96387430",
X"70780670",
X"98170c77",
X"7131a417",
X"08525851",
X"538939a0",
X"140870a4",
X"160c5374",
X"7627b938",
X"7251eed9",
X"3f83e080",
X"0853810b",
X"83e08008",
X"278b3888",
X"140883e0",
X"80082688",
X"38800b81",
X"1534b039",
X"83e08008",
X"a4150c98",
X"14081598",
X"150c7575",
X"3156c439",
X"98140816",
X"7098160c",
X"735256ef",
X"c83f83e0",
X"80088c38",
X"83e08008",
X"81153481",
X"55943982",
X"1433ff05",
X"76892a06",
X"83e08008",
X"05a8150c",
X"80557483",
X"e0800c88",
X"3d0d04ef",
X"3d0d6356",
X"855583e0",
X"9808802e",
X"80d23893",
X"3df40584",
X"170c6453",
X"883d7053",
X"765257f1",
X"d23f83e0",
X"80085583",
X"e08008b4",
X"38883d33",
X"5473802e",
X"a13802a7",
X"05337084",
X"2a708106",
X"51555583",
X"5573802e",
X"97387651",
X"eef83f83",
X"e0800888",
X"170c7551",
X"efa93f83",
X"e0800855",
X"7483e080",
X"0c933d0d",
X"04e43d0d",
X"6ea13d08",
X"405e8556",
X"83e09808",
X"802e8485",
X"389e3df4",
X"05841f0c",
X"7e98387d",
X"51eef83f",
X"83e08008",
X"5683ee39",
X"814181f6",
X"39834181",
X"f139933d",
X"7f960541",
X"59807f82",
X"95055e56",
X"756081ff",
X"05348341",
X"901e0876",
X"2e81d338",
X"a0547d22",
X"70852b83",
X"e0065458",
X"901e0852",
X"78518698",
X"3f83e080",
X"084183e0",
X"8008ffb8",
X"3878335c",
X"7b802eff",
X"b4388b19",
X"3370bf06",
X"71810652",
X"43557480",
X"2e80de38",
X"7b81bf06",
X"55748f24",
X"80d3389a",
X"19335574",
X"80cb38f3",
X"1d70585d",
X"8156758b",
X"2e098106",
X"85388e56",
X"8b39759a",
X"2e098106",
X"83389c56",
X"75197070",
X"81055233",
X"7133811a",
X"821a5f5b",
X"525b5574",
X"86387977",
X"34853980",
X"df773477",
X"7b57577a",
X"a02e0981",
X"06c03881",
X"567b81e5",
X"32703070",
X"9f2a5151",
X"557bae2e",
X"93387480",
X"2e8e3861",
X"832a7081",
X"06515574",
X"802e9738",
X"7d51ede2",
X"3f83e080",
X"084183e0",
X"80088738",
X"901e08fe",
X"af388060",
X"3475802e",
X"88387c52",
X"7f5183a5",
X"3f60802e",
X"8638800b",
X"901f0c60",
X"5660832e",
X"85386081",
X"d038891f",
X"57901e08",
X"802e81a8",
X"38805675",
X"19703351",
X"5574a02e",
X"a0387485",
X"2e098106",
X"843881e5",
X"55747770",
X"81055934",
X"81167081",
X"ff065755",
X"877627d7",
X"38881933",
X"5574a02e",
X"a938ae77",
X"70810559",
X"34885675",
X"19703351",
X"5574a02e",
X"95387477",
X"70810559",
X"34811670",
X"81ff0657",
X"558a7627",
X"e2388b19",
X"337f8805",
X"349f1933",
X"9e1a3371",
X"982b7190",
X"2b079d1c",
X"3370882b",
X"72079c1e",
X"33710764",
X"0c52991d",
X"33981e33",
X"71882b07",
X"53515357",
X"5956747f",
X"84052397",
X"1933961a",
X"3371882b",
X"07565674",
X"7f860523",
X"8077347d",
X"51ebf33f",
X"83e08008",
X"83327030",
X"7072079f",
X"2c83e080",
X"08065256",
X"56961f33",
X"55748a38",
X"891f5296",
X"1f5181b1",
X"3f7583e0",
X"800c9e3d",
X"0d04fd3d",
X"0d757753",
X"54733351",
X"70893871",
X"33517080",
X"2ea13873",
X"33723352",
X"53727127",
X"8538ff51",
X"94397073",
X"27853881",
X"518b3981",
X"14811353",
X"54d33980",
X"517083e0",
X"800c853d",
X"0d04fd3d",
X"0d757754",
X"54723370",
X"81ff0652",
X"5270802e",
X"a3387181",
X"ff068114",
X"ffbf1253",
X"54527099",
X"268938a0",
X"127081ff",
X"06535171",
X"74708105",
X"5634d239",
X"80743485",
X"3d0d04ff",
X"bd3d0d80",
X"c63d0852",
X"a53d7052",
X"54ffb33f",
X"80c73d08",
X"52853d70",
X"5253ffa6",
X"3f725273",
X"51fedf3f",
X"80c53d0d",
X"04fe3d0d",
X"74765353",
X"71708105",
X"53335170",
X"73708105",
X"553470f0",
X"38843d0d",
X"04fe3d0d",
X"74528072",
X"33525370",
X"732e8d38",
X"81128114",
X"71335354",
X"5270f538",
X"7283e080",
X"0c843d0d",
X"04fc3d0d",
X"76557483",
X"e398082e",
X"af388053",
X"745187c1",
X"3f83e080",
X"0881ff06",
X"ff147081",
X"ff067230",
X"709f2a51",
X"52555354",
X"72802e84",
X"3871dd38",
X"73fe3874",
X"83e3980c",
X"863d0d04",
X"ff3d0dff",
X"0b83e398",
X"0c84a53f",
X"81518785",
X"3f83e080",
X"0881ff06",
X"5271ee38",
X"81d33f71",
X"83e0800c",
X"833d0d04",
X"fc3d0d76",
X"028405a2",
X"05220288",
X"05a60522",
X"7a545555",
X"55ff823f",
X"72802ea0",
X"3883e3ac",
X"14337570",
X"81055734",
X"81147083",
X"ffff06ff",
X"157083ff",
X"ff065652",
X"5552dd39",
X"800b83e0",
X"800c863d",
X"0d04fc3d",
X"0d76787a",
X"11565355",
X"80537174",
X"2e933872",
X"15517033",
X"83e3ac13",
X"34811281",
X"145452ea",
X"39800b83",
X"e0800c86",
X"3d0d04fd",
X"3d0d9054",
X"83e39808",
X"5186f43f",
X"83e08008",
X"81ff06ff",
X"15713071",
X"30707307",
X"9f2a729f",
X"2a065255",
X"52555372",
X"db38853d",
X"0d04803d",
X"0d83e3a4",
X"081083e3",
X"9c080790",
X"80a80c82",
X"3d0d0480",
X"0b83e3a4",
X"0ce43f04",
X"810b83e3",
X"a40cdb3f",
X"04ed3f04",
X"7183e3a0",
X"0c04803d",
X"0d8051f4",
X"3f810b83",
X"e3a40c81",
X"0b83e39c",
X"0cffbb3f",
X"823d0d04",
X"803d0d72",
X"30707407",
X"802583e3",
X"9c0c51ff",
X"a53f823d",
X"0d04803d",
X"0d028b05",
X"339080a4",
X"0c9080a8",
X"08708106",
X"515170f5",
X"389080a4",
X"087081ff",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d81ff51",
X"d13f83e0",
X"800881ff",
X"0683e080",
X"0c823d0d",
X"04803d0d",
X"73902b73",
X"079080b4",
X"0c823d0d",
X"0404fb3d",
X"0d780284",
X"059f0533",
X"70982b55",
X"57557280",
X"259b3875",
X"80ff0656",
X"805280f7",
X"51e03f83",
X"e0800881",
X"ff065473",
X"812680ff",
X"388051fe",
X"e73fffa2",
X"3f8151fe",
X"df3fff9a",
X"3f7551fe",
X"ed3f7498",
X"2a51fee6",
X"3f74902a",
X"7081ff06",
X"5253feda",
X"3f74882a",
X"7081ff06",
X"5253fece",
X"3f7481ff",
X"0651fec6",
X"3f815575",
X"80c02e09",
X"81068638",
X"8195558d",
X"397580c8",
X"2e098106",
X"84388187",
X"557451fe",
X"a53f8a55",
X"fec83f83",
X"e0800881",
X"ff067098",
X"2b545472",
X"80258c38",
X"ff157081",
X"ff065653",
X"74e23873",
X"83e0800c",
X"873d0d04",
X"fa3d0dfd",
X"c53f8051",
X"fdda3f8a",
X"54fe933f",
X"ff147081",
X"ff065553",
X"73f33873",
X"74535580",
X"c051fea6",
X"3f83e080",
X"0881ff06",
X"5473812e",
X"09810682",
X"9f3883aa",
X"5280c851",
X"fe8c3f83",
X"e0800881",
X"ff065372",
X"812e0981",
X"0681a838",
X"7454873d",
X"74115456",
X"fdc83f83",
X"e0800873",
X"34811470",
X"81ff0655",
X"53837427",
X"e538029a",
X"05335372",
X"812e0981",
X"0681d938",
X"029b0533",
X"5380ce90",
X"547281aa",
X"2e8d3881",
X"c73980e4",
X"518a893f",
X"ff145473",
X"802e81b8",
X"38820a52",
X"81e951fd",
X"a53f83e0",
X"800881ff",
X"065372de",
X"38725280",
X"fa51fd92",
X"3f83e080",
X"0881ff06",
X"53728190",
X"38725473",
X"1653fcd6",
X"3f83e080",
X"08733481",
X"147081ff",
X"06555383",
X"7427e838",
X"873d3370",
X"862a7081",
X"06515454",
X"8c557280",
X"e3388455",
X"80de3974",
X"5281e951",
X"fccc3f83",
X"e0800881",
X"ff065382",
X"5581e956",
X"81732786",
X"38735580",
X"c15680ce",
X"90548a39",
X"80e45188",
X"fb3fff14",
X"5473802e",
X"a9388052",
X"7551fc9a",
X"3f83e080",
X"0881ff06",
X"5372e138",
X"84805280",
X"d051fc86",
X"3f83e080",
X"0881ff06",
X"5372802e",
X"83388055",
X"7483e3a8",
X"348051fb",
X"873ffbc2",
X"3f883d0d",
X"04fb3d0d",
X"7754800b",
X"83e3a833",
X"70832a70",
X"81065155",
X"57557275",
X"2e098106",
X"85387389",
X"2b547352",
X"80d151fb",
X"bd3f83e0",
X"800881ff",
X"065372bd",
X"3882b8c0",
X"54fb833f",
X"83e08008",
X"81ff0653",
X"7281ff2e",
X"09810689",
X"38ff1454",
X"73e7389f",
X"397281fe",
X"2e098106",
X"963883e7",
X"ac5283e3",
X"ac51faed",
X"3ffad33f",
X"fad03f83",
X"39815580",
X"51fa893f",
X"fac43f74",
X"81ff0683",
X"e0800c87",
X"3d0d04fb",
X"3d0d7783",
X"e3ac5654",
X"8151f9ec",
X"3f83e3a8",
X"3370832a",
X"70810651",
X"54567285",
X"3873892b",
X"54735280",
X"d851fab6",
X"3f83e080",
X"0881ff06",
X"537280e4",
X"3881ff51",
X"f9d43f81",
X"fe51f9ce",
X"3f848053",
X"74708105",
X"563351f9",
X"c13fff13",
X"7083ffff",
X"06515372",
X"eb387251",
X"f9b03f72",
X"51f9ab3f",
X"f9d03f83",
X"e080089f",
X"0653a788",
X"5472852e",
X"8c389939",
X"80e45186",
X"b33fff14",
X"54f9b33f",
X"83e08008",
X"81ff2e84",
X"3873e938",
X"8051f8e4",
X"3ff99f3f",
X"800b83e0",
X"800c873d",
X"0d047183",
X"e7b00c88",
X"80800b83",
X"e7ac0c84",
X"80800b83",
X"e7b40c04",
X"fd3d0d77",
X"70175577",
X"05ff1a53",
X"5371ff2e",
X"94387370",
X"81055533",
X"51707370",
X"81055534",
X"ff1252e9",
X"39853d0d",
X"04fc3d0d",
X"87a68155",
X"743383e7",
X"b834a054",
X"83a08053",
X"83e7b008",
X"5283e7ac",
X"0851ffb8",
X"3fa05483",
X"a4805383",
X"e7b00852",
X"83e7ac08",
X"51ffa53f",
X"905483a8",
X"805383e7",
X"b0085283",
X"e7ac0851",
X"ff923fa0",
X"53805283",
X"e7b40883",
X"a0800551",
X"858b3fa0",
X"53805283",
X"e7b40883",
X"a4800551",
X"84fb3f90",
X"53805283",
X"e7b40883",
X"a8800551",
X"84eb3fff",
X"753483a0",
X"80548053",
X"83e7b008",
X"5283e7b4",
X"0851fecc",
X"3f80d080",
X"5483b080",
X"5383e7b0",
X"085283e7",
X"b40851fe",
X"b73f8691",
X"3fa25480",
X"5383e7b4",
X"088c8005",
X"5280f4ec",
X"51fea13f",
X"860b87a8",
X"8334800b",
X"87a88234",
X"800b87a0",
X"9a34af0b",
X"87a09634",
X"bf0b87a0",
X"9734800b",
X"87a09834",
X"9f0b87a0",
X"9934800b",
X"87a09b34",
X"e00b87a8",
X"8934a20b",
X"87a88034",
X"830b87a4",
X"8f34820b",
X"87a88134",
X"863d0d04",
X"fd3d0d83",
X"a0805480",
X"5383e7b4",
X"085283e7",
X"b00851fd",
X"bf3f80d0",
X"805483b0",
X"805383e7",
X"b4085283",
X"e7b00851",
X"fdaa3fa0",
X"5483a080",
X"5383e7b4",
X"085283e7",
X"b00851fd",
X"973fa054",
X"83a48053",
X"83e7b408",
X"5283e7b0",
X"0851fd84",
X"3f905483",
X"a8805383",
X"e7b40852",
X"83e7b008",
X"51fcf13f",
X"83e7b833",
X"87a68134",
X"853d0d04",
X"803d0d90",
X"80900881",
X"0683e080",
X"0c823d0d",
X"04ff3d0d",
X"90809070",
X"0870fe06",
X"7607720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870812c",
X"810683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fd067610",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70822cbf",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"83067682",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870882c",
X"870683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"f1ff0676",
X"882b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"9008708b",
X"2cbf0683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f88fff",
X"06768b2b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70912cbf",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870fc",
X"87ffff06",
X"76912b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80800870",
X"882c8106",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"70892c81",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708a2c",
X"810683e0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708b",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"fe3d0d74",
X"81e62987",
X"2a9080a0",
X"0c843d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727081",
X"055434ff",
X"1151f039",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708405",
X"540cff11",
X"51f03984",
X"3d0d04fe",
X"3d0d8480",
X"80538052",
X"88800a51",
X"ffb33f81",
X"80805380",
X"5282800a",
X"51c63f84",
X"3d0d0480",
X"3d0d8151",
X"fcbf3f72",
X"802e8338",
X"d23f8151",
X"fcdd3f80",
X"51fcd83f",
X"8051fca9",
X"3f823d0d",
X"04fd3d0d",
X"75528054",
X"80ff7225",
X"8838810b",
X"ff801353",
X"54ffbf12",
X"51709926",
X"8638e012",
X"529e39ff",
X"9f125199",
X"71279538",
X"d012e013",
X"70545451",
X"89712788",
X"388f7327",
X"83388052",
X"73802e85",
X"38818012",
X"527181ff",
X"0683e080",
X"0c853d0d",
X"04803d0d",
X"84d8c051",
X"80717081",
X"05533470",
X"84e0c02e",
X"098106f0",
X"38823d0d",
X"04fe3d0d",
X"02970533",
X"51ff863f",
X"83e08008",
X"81ff0683",
X"e7bc0854",
X"52807324",
X"9b3883e7",
X"d8081372",
X"83e7dc08",
X"07535371",
X"733483e7",
X"bc088105",
X"83e7bc0c",
X"843d0d04",
X"fa3d0d82",
X"800a1b55",
X"8057883d",
X"fc055479",
X"53745278",
X"51cca43f",
X"883d0d04",
X"fe3d0d83",
X"e7d40852",
X"7451d388",
X"3f83e080",
X"088c3876",
X"53755283",
X"e7d40851",
X"c73f843d",
X"0d04fe3d",
X"0d83e7d4",
X"08537552",
X"7451cdc7",
X"3f83e080",
X"088d3877",
X"53765283",
X"e7d40851",
X"ffa23f84",
X"3d0d04fe",
X"3d0d83e7",
X"d40851cc",
X"bb3f83e0",
X"80088180",
X"802e0981",
X"068738b1",
X"8080539a",
X"3983e7d4",
X"0851cca0",
X"3f83e080",
X"0880d080",
X"2e098106",
X"9238b1b0",
X"805383e0",
X"80085283",
X"e7d40851",
X"feda3f84",
X"3d0d0480",
X"3d0dfab6",
X"3f83e080",
X"08842980",
X"f5900570",
X"0883e080",
X"0c51823d",
X"0d04ee3d",
X"0d804380",
X"42804180",
X"705a5bfd",
X"d43f800b",
X"83e7bc0c",
X"800b83e7",
X"dc0c80f2",
X"ec51c78d",
X"3f81800b",
X"83e7dc0c",
X"80f2f051",
X"c6ff3f80",
X"d00b83e7",
X"bc0c7830",
X"707a0780",
X"2570872b",
X"83e7dc0c",
X"5155f9a9",
X"3f83e080",
X"085280f2",
X"f851c6d9",
X"3f80f80b",
X"83e7bc0c",
X"78813270",
X"30707207",
X"80257087",
X"2b83e7dc",
X"0c515656",
X"fef13f83",
X"e0800852",
X"80f38451",
X"c6af3f81",
X"a00b83e7",
X"bc0c7882",
X"32703070",
X"72078025",
X"70872b83",
X"e7dc0c51",
X"5683e7d4",
X"085256c7",
X"c93f83e0",
X"80085280",
X"f38c51c6",
X"803f81f0",
X"0b83e7bc",
X"0c810b83",
X"e7c05b58",
X"83e7bc08",
X"82197a32",
X"70307072",
X"07802570",
X"872b83e7",
X"dc0c5157",
X"8e3d7055",
X"ff1b5457",
X"57579991",
X"3f797084",
X"055b0851",
X"c7803f74",
X"5483e080",
X"08537752",
X"80f39451",
X"c5b33fa8",
X"1783e7bc",
X"0c811858",
X"77852e09",
X"8106ffb0",
X"3883900b",
X"83e7bc0c",
X"78873270",
X"30707207",
X"80257087",
X"2b83e7dc",
X"0c515656",
X"f8cf3f80",
X"f3a45583",
X"e0800880",
X"2e8e3883",
X"e7d00851",
X"c6ac3f83",
X"e0800855",
X"745280f3",
X"ac51c4e1",
X"3f83e00b",
X"83e7bc0c",
X"78883270",
X"30707207",
X"80257087",
X"2b83e7dc",
X"0c515780",
X"f3b85255",
X"c4bf3f86",
X"8da051f9",
X"873f8052",
X"913d7052",
X"5599e33f",
X"83527451",
X"99dc3f61",
X"19597880",
X"25853880",
X"59903988",
X"79258538",
X"88598739",
X"78882682",
X"db387882",
X"2b5580f1",
X"c8150804",
X"f6c33f83",
X"e0800861",
X"57557581",
X"2e098106",
X"893883e0",
X"80081055",
X"903975ff",
X"2e098106",
X"883883e0",
X"8008812c",
X"55907525",
X"85389055",
X"88397480",
X"24833881",
X"557451f6",
X"9d3f8290",
X"39f6af3f",
X"83e08008",
X"61055574",
X"80258538",
X"80558839",
X"87752583",
X"38875574",
X"51f6a83f",
X"81ee3960",
X"87386280",
X"2e81e538",
X"83e0a408",
X"83e0a00c",
X"8aea0b83",
X"e0a80c83",
X"e7d40851",
X"ffb5dd3f",
X"fae93f81",
X"c7396056",
X"80762599",
X"388a830b",
X"83e0a80c",
X"83e7b415",
X"70085255",
X"ffb5bd3f",
X"74085291",
X"39758025",
X"913883e7",
X"b4150851",
X"c49a3f80",
X"52fd1951",
X"b8396280",
X"2e818d38",
X"83e7b415",
X"700883e7",
X"c008720c",
X"83e7c00c",
X"fd1a7053",
X"51558b81",
X"3f83e080",
X"08568051",
X"8af73f83",
X"e0800852",
X"7451878f",
X"3f755280",
X"5187883f",
X"80d63960",
X"55807525",
X"b83883e0",
X"ac0883e0",
X"a00c8aea",
X"0b83e0a8",
X"0c83e7d0",
X"0851ffb4",
X"c73f83e7",
X"d00851ff",
X"b2d63f83",
X"e0800881",
X"ff067052",
X"55f5b33f",
X"74802e9c",
X"388155a0",
X"39748025",
X"933883e7",
X"d00851c3",
X"8b3f8051",
X"f5983f84",
X"39628738",
X"7a802efa",
X"8a388055",
X"7483e080",
X"0c943d0d",
X"04fe3d0d",
X"f5963f83",
X"e0800880",
X"2e863880",
X"5180f739",
X"f59b3f83",
X"e0800880",
X"eb38f5bb",
X"3f83e080",
X"08802eaa",
X"388151f2",
X"f83feff1",
X"3f800b83",
X"e7bc0cf9",
X"b93f83e0",
X"800853ff",
X"0b83e7bc",
X"0cf1dd3f",
X"72be3872",
X"51f2d63f",
X"bc39f4f2",
X"3f83e080",
X"08802eb1",
X"388151f2",
X"c43fefbd",
X"3f8a830b",
X"83e0a80c",
X"83e7c008",
X"51ffb38c",
X"3fff0b83",
X"e7bc0cf1",
X"a73f83e7",
X"c0085280",
X"5185983f",
X"8151f5d3",
X"3f843d0d",
X"04fc3d0d",
X"84808052",
X"84a48080",
X"51c5de3f",
X"83e08008",
X"80c33888",
X"e93f80f6",
X"e451ca9e",
X"3f83e080",
X"0855b080",
X"805480c0",
X"805380f3",
X"c05283e0",
X"800851f7",
X"a13f83e7",
X"d4085380",
X"f3d05274",
X"51c4e83f",
X"83e08008",
X"8438f7af",
X"3f8151f4",
X"fa3f92f5",
X"3f8151f4",
X"f23ffe91",
X"3ffc3983",
X"e08c0802",
X"83e08c0c",
X"fb3d0d02",
X"80f3dc0b",
X"83e0a40c",
X"80f3e00b",
X"83e09c0c",
X"80f3e40b",
X"83e0ac0c",
X"83e08c08",
X"fc050c80",
X"0b83e7c0",
X"0b83e08c",
X"08f8050c",
X"83e08c08",
X"f4050cc3",
X"c03f83e0",
X"80088605",
X"fc0683e0",
X"8c08f005",
X"0c0283e0",
X"8c08f005",
X"08310d83",
X"3d7083e0",
X"8c08f805",
X"08708405",
X"83e08c08",
X"f8050c0c",
X"51c0893f",
X"83e08c08",
X"f4050881",
X"0583e08c",
X"08f4050c",
X"83e08c08",
X"f4050886",
X"2e098106",
X"ffad3884",
X"a8808051",
X"ecd43fff",
X"0b83e7bc",
X"0c800b83",
X"e7dc0c84",
X"d8c00b83",
X"e7d80c81",
X"51effe3f",
X"8151f0a3",
X"3f8051f0",
X"9e3f8151",
X"f0c43f81",
X"51f1993f",
X"8251f0e7",
X"3f8051f1",
X"bd3f80cf",
X"8d528051",
X"ffbdc73f",
X"fdbf3f83",
X"e08c08fc",
X"05080d80",
X"0b83e080",
X"0c873d0d",
X"83e08c0c",
X"04803d0d",
X"81ff5180",
X"0b83e7e8",
X"1234ff11",
X"5170f438",
X"823d0d04",
X"ff3d0d73",
X"70335351",
X"81113371",
X"34718112",
X"34833d0d",
X"04fb3d0d",
X"77795656",
X"80707155",
X"55527175",
X"25ac3872",
X"16703370",
X"147081ff",
X"06555151",
X"51717427",
X"89388112",
X"7081ff06",
X"53517181",
X"147083ff",
X"ff065552",
X"54747324",
X"d6387183",
X"e0800c87",
X"3d0d04fc",
X"3d0d7655",
X"ffb6f33f",
X"83e08008",
X"802ef538",
X"83ea8408",
X"86057081",
X"ff065253",
X"ffb4f33f",
X"8439fb81",
X"3fffb6d2",
X"3f83e080",
X"08812ef2",
X"38805473",
X"1553ffb5",
X"b83f83e0",
X"80087334",
X"81145473",
X"852e0981",
X"06e93884",
X"39fad63f",
X"ffb6a73f",
X"83e08008",
X"802ef238",
X"743383e7",
X"e8348115",
X"3383e7e9",
X"34821533",
X"83e7ea34",
X"83153383",
X"e7eb3484",
X"5283e7e8",
X"51feba3f",
X"83e08008",
X"81ff0684",
X"16335653",
X"72752e09",
X"81068d38",
X"ffb59c3f",
X"83e08008",
X"802e9a38",
X"83ea8408",
X"a82e0981",
X"06893886",
X"0b83ea84",
X"0c8739a8",
X"0b83ea84",
X"0c80e451",
X"efd63f86",
X"3d0d04f4",
X"3d0d7e60",
X"5955805d",
X"8075822b",
X"7183ea88",
X"120c83ea",
X"9c175b5b",
X"57767934",
X"77772e83",
X"b8387652",
X"7751ffbe",
X"d23f8e3d",
X"fc055490",
X"5383e9f0",
X"527751ff",
X"be8d3f7c",
X"5675902e",
X"09810683",
X"943883e9",
X"f051fd94",
X"3f83e9f2",
X"51fd8d3f",
X"83e9f451",
X"fd863f76",
X"83ea800c",
X"7751ffbb",
X"d93f80f1",
X"fc5283e0",
X"800851ff",
X"ab933f83",
X"e0800881",
X"2e098106",
X"80d43876",
X"83ea980c",
X"820b83e9",
X"f034ff96",
X"0b83e9f1",
X"347751ff",
X"be9e3f83",
X"e0800855",
X"83e08008",
X"77258838",
X"83e08008",
X"8f055574",
X"842c7083",
X"ffff0670",
X"882a5851",
X"557583e9",
X"f2347483",
X"e9f33476",
X"83e9f434",
X"ff800b83",
X"e9f53481",
X"903983e9",
X"f03383e9",
X"f1337188",
X"2b07565b",
X"7483ffff",
X"2e098106",
X"80e838fe",
X"800b83ea",
X"980c810b",
X"83ea800c",
X"ff0b83e9",
X"f034ff0b",
X"83e9f134",
X"7751ffbd",
X"ab3f83e0",
X"800883ea",
X"a00c83e0",
X"80085583",
X"e0800880",
X"25883883",
X"e080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583e9f2",
X"347483e9",
X"f3347683",
X"e9f434ff",
X"800b83e9",
X"f534810b",
X"83e9ff34",
X"a5397485",
X"962e0981",
X"0680fe38",
X"7583ea98",
X"0c7751ff",
X"bcdf3f83",
X"e9ff3383",
X"e0800807",
X"557483e9",
X"ff3483e9",
X"ff338106",
X"5574802e",
X"83388457",
X"83e9f433",
X"83e9f533",
X"71882b07",
X"565c7481",
X"802e0981",
X"06a13883",
X"e9f23383",
X"e9f33371",
X"882b0756",
X"5bad8075",
X"27873876",
X"8207579c",
X"39768107",
X"57963974",
X"82802e09",
X"81068738",
X"76830757",
X"87397481",
X"ff268a38",
X"7783ea88",
X"1b0c7679",
X"348e3d0d",
X"04803d0d",
X"72842983",
X"ea880570",
X"0883e080",
X"0c51823d",
X"0d04fe3d",
X"0d800b83",
X"e9ec0c80",
X"0b83e9e8",
X"0cff0b83",
X"e7e40ca8",
X"0b83ea84",
X"0cae51ff",
X"afbc3f80",
X"0b83ea88",
X"54528073",
X"70840555",
X"0c811252",
X"71842e09",
X"8106ef38",
X"843d0d04",
X"fe3d0d74",
X"02840596",
X"05225353",
X"71802e97",
X"38727081",
X"05543351",
X"ffafc63f",
X"ff127083",
X"ffff0651",
X"52e63984",
X"3d0d04fe",
X"3d0d0292",
X"05225382",
X"ac51eae8",
X"3f80c351",
X"ffafa23f",
X"819651ea",
X"db3f7252",
X"83e7e851",
X"ffb23f72",
X"5283e7e8",
X"51f8ee3f",
X"83e08008",
X"81ff0651",
X"ffaefe3f",
X"843d0d04",
X"ffb13d0d",
X"80d13df8",
X"0551f997",
X"3f83e9ec",
X"08810583",
X"e9ec0c80",
X"cf3d33cf",
X"117081ff",
X"06515656",
X"74832688",
X"ed38758f",
X"06ff0556",
X"7583e7e4",
X"082e9b38",
X"75832696",
X"387583e7",
X"e40c7584",
X"2983ea88",
X"05700853",
X"557551fa",
X"963f8076",
X"2488c938",
X"75842983",
X"ea880555",
X"7408802e",
X"88ba3883",
X"e7e40884",
X"2983ea88",
X"05700802",
X"880582b9",
X"0533525b",
X"557480d2",
X"2e84b138",
X"7480d224",
X"903874bf",
X"2e9c3874",
X"80d02e81",
X"d73887f8",
X"397480d3",
X"2e80d238",
X"7480d72e",
X"81c63887",
X"e7390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290556",
X"56ffadfa",
X"3f80c151",
X"ffadb23f",
X"f6e73f86",
X"0b83e7e8",
X"34815283",
X"e7e851ff",
X"aed53f81",
X"51fde43f",
X"74893886",
X"0b83ea84",
X"0c8739a8",
X"0b83ea84",
X"0cffadc6",
X"3f80c151",
X"ffacfe3f",
X"f6b33f90",
X"0b83e9ff",
X"33810656",
X"5674802e",
X"83389856",
X"83e9f433",
X"83e9f533",
X"71882b07",
X"56597481",
X"802e0981",
X"069c3883",
X"e9f23383",
X"e9f33371",
X"882b0756",
X"57ad8075",
X"278c3875",
X"81800756",
X"853975a0",
X"07567583",
X"e7e834ff",
X"0b83e7e9",
X"34e00b83",
X"e7ea3480",
X"0b83e7eb",
X"34845283",
X"e7e851ff",
X"adc93f84",
X"51869e39",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"055659ff",
X"acb83f79",
X"51ffb7a5",
X"3f83e080",
X"08802e8b",
X"3880ce51",
X"ffabe23f",
X"85f23980",
X"c151ffab",
X"d83fffac",
X"cd3fffab",
X"803f83ea",
X"98085883",
X"75259b38",
X"83e9f433",
X"83e9f533",
X"71882b07",
X"fc177129",
X"7a058380",
X"055a5157",
X"8d397481",
X"802918ff",
X"80055881",
X"80578056",
X"76762e93",
X"38ffabb1",
X"3f83e080",
X"0883e7e8",
X"17348116",
X"56ea39ff",
X"ab9f3f83",
X"e0800881",
X"ff067753",
X"83e7e852",
X"56f4d63f",
X"83e08008",
X"81ff0655",
X"75752e09",
X"8106818a",
X"38ffab9e",
X"3f80c151",
X"ffaad63f",
X"ffabcb3f",
X"77527951",
X"ffb5b43f",
X"805e80d1",
X"3dfdf405",
X"54765383",
X"e7e85279",
X"51ffb3c1",
X"3f0282b9",
X"05335581",
X"587480d7",
X"2e098106",
X"bd3880d1",
X"3dfdf005",
X"5476538f",
X"3d70537a",
X"5259ffb4",
X"c63f8056",
X"76762ea2",
X"38751983",
X"e7e81733",
X"71337072",
X"32703070",
X"80257030",
X"7e06811d",
X"5d5e5151",
X"51525b55",
X"db3982ac",
X"51e5a13f",
X"77802e86",
X"3880c351",
X"843980ce",
X"51ffa9d1",
X"3fffaac6",
X"3fffa8f9",
X"3f83dd39",
X"0282bb05",
X"33028405",
X"82ba0533",
X"71828029",
X"05595580",
X"705d59ff",
X"a9ec3f80",
X"c151ffa9",
X"a43f83ea",
X"8008792e",
X"82de3883",
X"eaa00880",
X"fc055580",
X"fd527451",
X"86d73f83",
X"e080085b",
X"778224b2",
X"38ff1870",
X"872b83ff",
X"ff800680",
X"f5b00583",
X"e7e85957",
X"55818055",
X"75708105",
X"57337770",
X"81055934",
X"ff157081",
X"ff065155",
X"74ea3882",
X"8d397782",
X"e82e81ab",
X"387782e9",
X"2e098106",
X"81b23880",
X"f3e851ff",
X"afa73f78",
X"58778732",
X"70307072",
X"0780257a",
X"8a327030",
X"70720780",
X"25730753",
X"545a5157",
X"5575802e",
X"97387878",
X"269238a0",
X"0b83e7e8",
X"1a348119",
X"7081ff06",
X"5a55eb39",
X"81187081",
X"ff065955",
X"8a7827ff",
X"bc388f58",
X"83e7e318",
X"3383e7e8",
X"1934ff18",
X"7081ff06",
X"59557784",
X"26ea3890",
X"58800b83",
X"e7e81934",
X"81187081",
X"ff067098",
X"2b525955",
X"748025e9",
X"3880c655",
X"7a858f24",
X"843880c2",
X"557483e7",
X"e83480f1",
X"0b83e7eb",
X"34810b83",
X"e7ec347a",
X"83e7e934",
X"7a882c55",
X"7483e7ea",
X"3480cb39",
X"82f07825",
X"80c43877",
X"80fd29fd",
X"97d30552",
X"7951ffb1",
X"e23f80d1",
X"3dfdec05",
X"5480fd53",
X"83e7e852",
X"7951ffb1",
X"9a3f7b81",
X"19595675",
X"80fc2483",
X"38785877",
X"882c5574",
X"83e8e534",
X"7783e8e6",
X"347583e8",
X"e7348180",
X"5980cc39",
X"83ea9808",
X"57837825",
X"9b3883e9",
X"f43383e9",
X"f5337188",
X"2b07fc1a",
X"71297905",
X"83800559",
X"51598d39",
X"77818029",
X"17ff8005",
X"57818059",
X"76527951",
X"ffb0f03f",
X"80d13dfd",
X"ec055478",
X"5383e7e8",
X"527951ff",
X"b0a93f78",
X"51f6b83f",
X"ffa6e33f",
X"ffa5963f",
X"8b3983e9",
X"e8088105",
X"83e9e80c",
X"80d13d0d",
X"04f6d93f",
X"eb9f3ff9",
X"39fc3d0d",
X"76787184",
X"2983ea88",
X"05700851",
X"53535370",
X"9e3880ce",
X"723480cf",
X"0b811334",
X"80ce0b82",
X"133480c5",
X"0b831334",
X"70841334",
X"80e73983",
X"ea9c1333",
X"5480d272",
X"3473822a",
X"70810651",
X"5180cf53",
X"70843880",
X"d7537281",
X"1334a00b",
X"82133473",
X"83065170",
X"812e9e38",
X"70812488",
X"3870802e",
X"8f389f39",
X"70822e92",
X"3870832e",
X"92389339",
X"80d8558e",
X"3980d355",
X"893980cd",
X"55843980",
X"c4557483",
X"133480c4",
X"0b841334",
X"800b8513",
X"34863d0d",
X"04fd3d0d",
X"75538073",
X"0c800b84",
X"140c800b",
X"88140c87",
X"a6803370",
X"81ff0670",
X"812a8132",
X"71813271",
X"81067181",
X"06318418",
X"0c555670",
X"832a8132",
X"71822a81",
X"32718106",
X"71810631",
X"770c5254",
X"515187a0",
X"90337009",
X"81068815",
X"0c51853d",
X"0d04fe3d",
X"0d747654",
X"527151ff",
X"a03f7281",
X"2ea23881",
X"73268d38",
X"72822eab",
X"3872832e",
X"9f38e639",
X"7108e238",
X"841208dd",
X"38881208",
X"d838a039",
X"88120881",
X"2e098106",
X"cc389439",
X"88120881",
X"2e8d3871",
X"08893884",
X"1208802e",
X"ffb73884",
X"3d0d04fc",
X"3d0d7678",
X"53548153",
X"80558739",
X"71107310",
X"54527372",
X"26517280",
X"2ea73870",
X"802e8638",
X"718025e8",
X"3872802e",
X"98387174",
X"26893873",
X"72317574",
X"07565472",
X"812a7281",
X"2a5353e5",
X"39735178",
X"83387451",
X"7083e080",
X"0c863d0d",
X"04fe3d0d",
X"80537552",
X"7451ffa3",
X"3f843d0d",
X"04fe3d0d",
X"81537552",
X"7451ff93",
X"3f843d0d",
X"04fb3d0d",
X"77795555",
X"80567476",
X"25863874",
X"30558156",
X"73802588",
X"38733076",
X"81325754",
X"80537352",
X"7451fee7",
X"3f83e080",
X"08547580",
X"2e873883",
X"e0800830",
X"547383e0",
X"800c873d",
X"0d04fa3d",
X"0d787a57",
X"55805774",
X"77258638",
X"74305581",
X"57759f2c",
X"54815375",
X"74327431",
X"527451fe",
X"aa3f83e0",
X"80085476",
X"802e8738",
X"83e08008",
X"30547383",
X"e0800c88",
X"3d0d0400",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002a3c",
X"00002a7d",
X"00002a9f",
X"00002ac6",
X"00002ac6",
X"00002ac6",
X"00002ac6",
X"00002b37",
X"00002b89",
X"25732025",
X"73000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"6e616d65",
X"20000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00003928",
X"0000392c",
X"00003934",
X"00003940",
X"0000394c",
X"00003958",
X"00003964",
X"00003968",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
