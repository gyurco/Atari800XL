
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f2",
X"d4738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80f5",
X"cc0c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580ed",
X"842d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580eb98",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"97b30480",
X"3d0d80f6",
X"f0087008",
X"810683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d80f6",
X"f0087008",
X"70fe0676",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80f6f008",
X"70087081",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80f6f008",
X"700870fd",
X"06761007",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"f6f00870",
X"0870822c",
X"bf0683e0",
X"800c5151",
X"823d0d04",
X"ff3d0d80",
X"f6f00870",
X"0870fe83",
X"0676822b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80f6f008",
X"70087088",
X"2c870683",
X"e0800c51",
X"51823d0d",
X"04ff3d0d",
X"80f6f008",
X"700870f1",
X"ff067688",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d80f6f0",
X"08700870",
X"8b2cbf06",
X"83e0800c",
X"5151823d",
X"0d04ff3d",
X"0d80f6f0",
X"08700870",
X"f88fff06",
X"768b2b07",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"f7800870",
X"0870882c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"f7800870",
X"0870892c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"f7800870",
X"08708a2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"f7800870",
X"08708b2c",
X"810683e0",
X"800c5151",
X"823d0d04",
X"fd3d0d75",
X"81e62987",
X"2a80f6e0",
X"0854730c",
X"853d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d848080",
X"53805288",
X"800a51ff",
X"b33f8180",
X"80538052",
X"82800a51",
X"c63f843d",
X"0d04803d",
X"0d8151fc",
X"ce3f7280",
X"2e8338d2",
X"3f8151fc",
X"f03f8051",
X"fceb3f80",
X"51fcb83f",
X"823d0d04",
X"fd3d0d75",
X"52805480",
X"ff722588",
X"38810bff",
X"80135354",
X"ffbf1251",
X"70992686",
X"38e01252",
X"9e39ff9f",
X"12519971",
X"279538d0",
X"12e01370",
X"54545189",
X"71278838",
X"8f732783",
X"38805273",
X"802e8538",
X"81801252",
X"7181ff06",
X"83e0800c",
X"853d0d04",
X"803d0d86",
X"b8c05180",
X"71708105",
X"53347086",
X"c0c02e09",
X"8106f038",
X"823d0d04",
X"fe3d0d02",
X"97053351",
X"ff863f83",
X"e0800881",
X"ff0683e0",
X"9c085452",
X"8073249b",
X"3883e0b8",
X"08137283",
X"e0bc0807",
X"53537173",
X"3483e09c",
X"08810583",
X"e09c0c84",
X"3d0d04fa",
X"3d0d8280",
X"0a1b5580",
X"57883dfc",
X"05547953",
X"74527851",
X"b7ae3f88",
X"3d0d04fe",
X"3d0d83e0",
X"b0085274",
X"51bde83f",
X"83e08008",
X"8c387653",
X"755283e0",
X"b00851c7",
X"3f843d0d",
X"04fe3d0d",
X"83e0b008",
X"53755274",
X"51b8af3f",
X"83e08008",
X"8d387753",
X"765283e0",
X"b00851ff",
X"a23f843d",
X"0d04fe3d",
X"0d83e0b4",
X"0851b7af",
X"3f83e080",
X"08818080",
X"2e098106",
X"883883c1",
X"8080539b",
X"3983e0b4",
X"0851b793",
X"3f83e080",
X"0880d080",
X"2e098106",
X"933883c1",
X"b0805383",
X"e0800852",
X"83e0b408",
X"51fed83f",
X"843d0d04",
X"803d0dfa",
X"cc3f83e0",
X"80088726",
X"80cd3883",
X"e0800884",
X"2980f2e4",
X"05517008",
X"040b0b80",
X"f3cc51b7",
X"390b0b80",
X"f3d051af",
X"390b0b80",
X"f3d851a7",
X"390b0b80",
X"f3e4519f",
X"390b0b80",
X"f3f05197",
X"390b0b80",
X"f3fc518f",
X"390b0b80",
X"f4885187",
X"390b0b80",
X"f48c5170",
X"83e0800c",
X"823d0d04",
X"ee3d0d80",
X"43804280",
X"4180705a",
X"5bfd893f",
X"800b83e0",
X"9c0c800b",
X"83e0bc0c",
X"0b0b80f4",
X"9051b19d",
X"3f81800b",
X"83e0bc0c",
X"0b0b80f4",
X"9451b18d",
X"3f80d00b",
X"83e09c0c",
X"7830707a",
X"07802570",
X"872b83e0",
X"bc0c5155",
X"f8ee3f83",
X"e0800852",
X"0b0b80f4",
X"9c51b0e5",
X"3f80f80b",
X"83e09c0c",
X"78813270",
X"30707207",
X"80257087",
X"2b83e0bc",
X"0c515656",
X"fea23f83",
X"e0800852",
X"0b0b80f4",
X"a851b0b9",
X"3f81a00b",
X"83e09c0c",
X"78823270",
X"30707207",
X"80257087",
X"2b83e0bc",
X"0c515683",
X"e0b40852",
X"56b1ff3f",
X"83e08008",
X"520b0b80",
X"f4b051b0",
X"883f81f0",
X"0b83e09c",
X"0c810b83",
X"e0a05b58",
X"83e09c08",
X"82197a32",
X"70307072",
X"07802570",
X"872b83e0",
X"bc0c5157",
X"8e3d7055",
X"ff1b5457",
X"5757a5e6",
X"3f797084",
X"055b0851",
X"b1b43f74",
X"5483e080",
X"08537752",
X"0b0b80f4",
X"b851afb9",
X"3fa81783",
X"e09c0c81",
X"18587785",
X"2e098106",
X"ffae3883",
X"900b83e0",
X"9c0c7887",
X"32703070",
X"72078025",
X"70872b83",
X"e0bc0c51",
X"560b0b80",
X"f4c85256",
X"af833f83",
X"e00b83e0",
X"9c0c7888",
X"32703070",
X"72078025",
X"70872b83",
X"e0bc0c51",
X"560b0b80",
X"f4dc5256",
X"aedf3f86",
X"8da051f8",
X"c73f8052",
X"913d7052",
X"558bd43f",
X"83527451",
X"8bcd3f61",
X"19597880",
X"25853880",
X"59903988",
X"79258538",
X"88598739",
X"78882682",
X"ae387882",
X"2b5580f3",
X"84150804",
X"f69a3f83",
X"e0800861",
X"57557581",
X"2e098106",
X"893883e0",
X"80081055",
X"903975ff",
X"2e098106",
X"883883e0",
X"8008812c",
X"55907525",
X"85389055",
X"88397480",
X"24833881",
X"557451f5",
X"f73f81e3",
X"39f68a3f",
X"83e08008",
X"61055574",
X"80258538",
X"80558839",
X"87752583",
X"38875574",
X"51f6863f",
X"81c13960",
X"87386280",
X"2e81b838",
X"a1d80b83",
X"e0d00c83",
X"e0b40851",
X"8d9f3ffa",
X"b53f81a3",
X"39605680",
X"76259838",
X"a0f70b83",
X"e0d00c83",
X"e0941570",
X"0852558d",
X"803f7408",
X"52913975",
X"80259138",
X"83e09415",
X"0851aef0",
X"3f8052fd",
X"1951b839",
X"62802e80",
X"ea3883e0",
X"94157008",
X"83e0a008",
X"720c83e0",
X"a00cfd1a",
X"70535155",
X"988d3f83",
X"e0800856",
X"80519883",
X"3f83e080",
X"08527451",
X"94853f75",
X"52805193",
X"fe3fb439",
X"62802eaf",
X"38a1d80b",
X"83e0d00c",
X"83e0b008",
X"518c963f",
X"83e0b008",
X"51adff3f",
X"9c800a53",
X"80c08052",
X"83e08008",
X"51f8d03f",
X"81558c39",
X"6287387a",
X"802efac5",
X"38805574",
X"83e0800c",
X"943d0d04",
X"fe3d0df4",
X"f73f83e0",
X"8008802e",
X"86388051",
X"80f639f4",
X"ff3f83e0",
X"800880ea",
X"38f5a53f",
X"83e08008",
X"802eaa38",
X"8151f2f7",
X"3f839b3f",
X"800b83e0",
X"9c0cf9f4",
X"3f83e080",
X"0853ff0b",
X"83e09c0c",
X"85ee3f72",
X"bd387251",
X"f2d53fbb",
X"39f4d93f",
X"83e08008",
X"802eb038",
X"8151f2c3",
X"3f82e73f",
X"a0f70b83",
X"e0d00c83",
X"e0a00851",
X"8af33fff",
X"0b83e09c",
X"0c85b93f",
X"83e0a008",
X"52805192",
X"b23f8151",
X"f5c43f84",
X"3d0d0483",
X"e08c0802",
X"83e08c0c",
X"fa3d0d80",
X"0b83e0a0",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"f8050caf",
X"a73f83e0",
X"80088605",
X"fc0683e0",
X"8c08f405",
X"0c0283e0",
X"8c08f405",
X"08310d85",
X"3d7083e0",
X"8c08fc05",
X"08708405",
X"83e08c08",
X"fc050c0c",
X"51ac853f",
X"83e08c08",
X"f8050881",
X"0583e08c",
X"08f8050c",
X"83e08c08",
X"f8050886",
X"2e098106",
X"ffad3886",
X"88808051",
X"81aa3fff",
X"0b83e09c",
X"0c800b83",
X"e0bc0c86",
X"b8c00b83",
X"e0b80c81",
X"51f1803f",
X"8151f1a9",
X"3f8051f1",
X"a43f8151",
X"f1ce3f81",
X"51f2ab3f",
X"8251f1f5",
X"3f8e8452",
X"8051a99e",
X"3f848080",
X"52868480",
X"8051af84",
X"3f83e080",
X"0880d338",
X"94e63f80",
X"f8b851b3",
X"bc3f83e0",
X"800883e0",
X"b408540b",
X"0b80f4e4",
X"5383e080",
X"085283e0",
X"8c08f405",
X"0cae973f",
X"83e08008",
X"8438f5f6",
X"3f9c800a",
X"5480c080",
X"530b0b80",
X"f4f05283",
X"e08c08f4",
X"050851f5",
X"b83f8151",
X"f3a83f9e",
X"cd3f8151",
X"f3a03ffc",
X"cf3ffc39",
X"7183e0c4",
X"0c888080",
X"0b83e0c0",
X"0c848080",
X"0b83e0c8",
X"0c04f03d",
X"0d80f5e8",
X"08547333",
X"83e0cc34",
X"83a08056",
X"83e0c408",
X"1683e0c0",
X"08175654",
X"74337434",
X"83e0c808",
X"16548074",
X"34811656",
X"7583a0a0",
X"2e098106",
X"db3883a4",
X"805683e0",
X"c4081683",
X"e0c00817",
X"56547433",
X"743483e0",
X"c8081654",
X"80743481",
X"16567583",
X"a4a02e09",
X"8106db38",
X"83a88056",
X"83e0c408",
X"1683e0c0",
X"08175654",
X"74337434",
X"83e0c808",
X"16548074",
X"34811656",
X"7583a890",
X"2e098106",
X"db3880f5",
X"e80854ff",
X"74348056",
X"83e0c408",
X"1683e0c8",
X"08175555",
X"73337534",
X"81165675",
X"83a0802e",
X"098106e4",
X"3883b080",
X"5683e0c4",
X"081683e0",
X"c8081755",
X"55733375",
X"34811656",
X"75848080",
X"2e098106",
X"e438f2a4",
X"3f893d58",
X"a25380f3",
X"a8527751",
X"80d5e63f",
X"80578c80",
X"5683e0c8",
X"08167719",
X"55557333",
X"75348116",
X"81185856",
X"76a22e09",
X"8106e638",
X"80f68c08",
X"54867434",
X"80f69008",
X"54807434",
X"80f68808",
X"54807434",
X"80f5f808",
X"54af7434",
X"80f68408",
X"54bf7434",
X"80f68008",
X"54807434",
X"80f5fc08",
X"549f7434",
X"80f5f408",
X"54807434",
X"80f5e008",
X"54e07434",
X"80f5d808",
X"54767434",
X"80f5d408",
X"54837434",
X"80f5dc08",
X"54827434",
X"923d0d04",
X"fe3d0d80",
X"5383e0c8",
X"081383e0",
X"c4081452",
X"52703372",
X"34811353",
X"7283a080",
X"2e098106",
X"e43883b0",
X"805383e0",
X"c8081383",
X"e0c40814",
X"52527033",
X"72348113",
X"53728480",
X"802e0981",
X"06e43883",
X"a0805383",
X"e0c80813",
X"83e0c408",
X"14525270",
X"33723481",
X"13537283",
X"a0a02e09",
X"8106e438",
X"83a48053",
X"83e0c808",
X"1383e0c4",
X"08145252",
X"70337234",
X"81135372",
X"83a4a02e",
X"098106e4",
X"3883a880",
X"5383e0c8",
X"081383e0",
X"c4081452",
X"52703372",
X"34811353",
X"7283a890",
X"2e098106",
X"e43880f5",
X"e8085183",
X"e0cc3371",
X"34843d0d",
X"04fe3d0d",
X"74538073",
X"0c800b84",
X"140c800b",
X"88140c80",
X"f5ec0870",
X"337081ff",
X"0670812a",
X"81327081",
X"06515254",
X"51517080",
X"2e883881",
X"0b84140c",
X"93397181",
X"32708106",
X"51517080",
X"2e8638ff",
X"0b84140c",
X"71832a81",
X"32708106",
X"51517080",
X"2e863881",
X"730c9339",
X"71822a81",
X"32708106",
X"51517080",
X"2e8438ff",
X"730c80f5",
X"e4087033",
X"70097081",
X"06515151",
X"5170802e",
X"8638810b",
X"88140c84",
X"3d0d04fe",
X"3d0d7476",
X"54527151",
X"feeb3f72",
X"812ea238",
X"8173268d",
X"3872822e",
X"ab387283",
X"2e9f38e6",
X"397108e2",
X"38841208",
X"dd388812",
X"08d838a0",
X"39881208",
X"812e0981",
X"06cc3894",
X"39881208",
X"812e8d38",
X"71088938",
X"84120880",
X"2effb738",
X"843d0d04",
X"ffb83d0d",
X"800b80cc",
X"3d08538b",
X"3d705359",
X"5480c6fe",
X"3f80cc3d",
X"085280ca",
X"3dfdfc05",
X"5180c6ee",
X"3f893d33",
X"028405a1",
X"05330288",
X"05a20533",
X"59575573",
X"18703351",
X"5372802e",
X"be3872ae",
X"2e863881",
X"1454ec39",
X"80ca3dfe",
X"81111570",
X"33515458",
X"74732e09",
X"8106a038",
X"fe821814",
X"70335153",
X"75732e09",
X"81069038",
X"fe831814",
X"53817333",
X"54547673",
X"2e833880",
X"547383e0",
X"800c80ca",
X"3d0d04fc",
X"3d0d7670",
X"5255acaf",
X"3f83e080",
X"08548153",
X"83e08008",
X"80c13874",
X"51abf23f",
X"83e08008",
X"80f59053",
X"83e08008",
X"5253fec8",
X"3f83e080",
X"08a13880",
X"f5945272",
X"51feb93f",
X"83e08008",
X"923880f5",
X"98527251",
X"feaa3f83",
X"e0800880",
X"2e833881",
X"54735372",
X"83e0800c",
X"863d0d04",
X"fd3d0d75",
X"705254ab",
X"ce3f8153",
X"83e08008",
X"97387351",
X"ab973f80",
X"f59c5283",
X"e0800851",
X"fdf23f83",
X"e0800853",
X"7283e080",
X"0c853d0d",
X"04e03d0d",
X"a33d0870",
X"525ea1e6",
X"3f83e080",
X"0833943d",
X"56547394",
X"3880f8c8",
X"52745184",
X"d1397d52",
X"7851a4d4",
X"3f84dc39",
X"7d51a1ce",
X"3f83e080",
X"08527451",
X"a0fe3f83",
X"e0d00852",
X"933d7052",
X"5ba7b13f",
X"83e08008",
X"59800b83",
X"e0800855",
X"5c83e080",
X"087c2e94",
X"38811c74",
X"525caab2",
X"3f83e080",
X"085483e0",
X"8008ee38",
X"805aff7a",
X"437a427a",
X"415f7909",
X"709f2c7b",
X"065b547b",
X"7a248438",
X"ff1c5af6",
X"1a700970",
X"9f2c7206",
X"7bff125a",
X"5a525555",
X"80752595",
X"387651a9",
X"f13f83e0",
X"800876ff",
X"18585557",
X"738024ed",
X"38747f2e",
X"8638eaa4",
X"3f745f78",
X"ff1b7058",
X"5e58807a",
X"25953877",
X"51a9c73f",
X"83e08008",
X"76ff1858",
X"55587380",
X"24ed3880",
X"0b83e09c",
X"0c800b83",
X"e0bc0c80",
X"f5a0519e",
X"983f8180",
X"0b83e0bc",
X"0c80f5a8",
X"519e8a3f",
X"a80b83e0",
X"9c0c7680",
X"2e80e438",
X"83e09c08",
X"77793270",
X"30707207",
X"80257087",
X"2b83e0bc",
X"0c515678",
X"535656a8",
X"fe3f83e0",
X"8008802e",
X"883880f5",
X"b0519dd1",
X"3f7651a8",
X"c03f83e0",
X"80085280",
X"f4c4519d",
X"c03f7651",
X"a8c83f83",
X"e0800883",
X"e09c0855",
X"57757425",
X"8638a816",
X"56f73975",
X"83e09c0c",
X"86f07624",
X"ff983887",
X"980b83e0",
X"9c0c7780",
X"2eb13877",
X"51a7fe3f",
X"83e08008",
X"785255a8",
X"9e3f80f5",
X"b85483e0",
X"80088d38",
X"87398076",
X"34fda039",
X"80f5b454",
X"74537352",
X"80f58051",
X"9cdf3f80",
X"5480f5c0",
X"519cd63f",
X"81145473",
X"a82e0981",
X"06ef3886",
X"8da051e6",
X"b33f8052",
X"903d7052",
X"54f9c03f",
X"83527351",
X"f9b93f61",
X"802e819d",
X"387c5473",
X"ff2e9638",
X"78802e81",
X"9e387851",
X"a7a83f83",
X"e08008ff",
X"155559e7",
X"3978802e",
X"81893878",
X"51a7a43f",
X"83e08008",
X"802efc96",
X"387851a6",
X"ec3f83e0",
X"800883e0",
X"80085380",
X"f5885254",
X"80c0933f",
X"83e08008",
X"a5387a51",
X"80c1ca3f",
X"83e08008",
X"5574ff16",
X"56548074",
X"25fbfc38",
X"741b7033",
X"555673af",
X"2efecb38",
X"e8397a51",
X"80c1a63f",
X"825380f5",
X"8c5283e0",
X"80081b51",
X"80cace3f",
X"7a5180c1",
X"903f7352",
X"83e08008",
X"1b5180c0",
X"e83ffbc3",
X"397f8829",
X"6010057a",
X"0561055a",
X"fbf439a2",
X"3d0d0480",
X"3d0d81ff",
X"51800b83",
X"e0dc1234",
X"ff115170",
X"f438823d",
X"0d04ff3d",
X"0d737033",
X"53518111",
X"33713471",
X"81123483",
X"3d0d04fb",
X"3d0d7779",
X"56568070",
X"71555552",
X"717525ac",
X"38721670",
X"33701470",
X"81ff0655",
X"51515171",
X"74278938",
X"81127081",
X"ff065351",
X"71811470",
X"83ffff06",
X"55525474",
X"7324d638",
X"7183e080",
X"0c873d0d",
X"04fd3d0d",
X"755494bb",
X"3f83e080",
X"08802ef6",
X"3883e2f8",
X"08860570",
X"81ff0652",
X"5392943f",
X"8439edfc",
X"3f949c3f",
X"83e08008",
X"812ef338",
X"92f73f83",
X"e0800874",
X"3492ee3f",
X"83e08008",
X"81153492",
X"e43f83e0",
X"80088215",
X"3492da3f",
X"83e08008",
X"83153492",
X"d03f83e0",
X"80088415",
X"348439ed",
X"bb3f93db",
X"3f83e080",
X"08802ef3",
X"38733383",
X"e0dc3481",
X"143383e0",
X"dd348214",
X"3383e0de",
X"34831433",
X"83e0df34",
X"845283e0",
X"dc51fea7",
X"3f83e080",
X"0881ff06",
X"84153355",
X"5372742e",
X"0981068c",
X"3892cc3f",
X"83e08008",
X"802e9a38",
X"83e2f808",
X"a82e0981",
X"06893886",
X"0b83e2f8",
X"0c8739a8",
X"0b83e2f8",
X"0c80e451",
X"e2aa3f85",
X"3d0d04f4",
X"3d0d7e60",
X"5a55805d",
X"8075822b",
X"7183e2fc",
X"120c83e3",
X"90175c5c",
X"56757a34",
X"78762e83",
X"ce387552",
X"78519cad",
X"3f8e3dfc",
X"05549053",
X"83e2e452",
X"78519bf0",
X"3f7c5877",
X"902e0981",
X"0683ac38",
X"83e2e451",
X"fd843f83",
X"e2e651fc",
X"fd3f83e2",
X"e851fcf6",
X"3f7583e2",
X"f40c7851",
X"99bc3f80",
X"f5945283",
X"e0800851",
X"f5a23f83",
X"e0800881",
X"2e098106",
X"80e33875",
X"83e38c0c",
X"820b83e2",
X"e434ff96",
X"0b83e2e5",
X"3478519b",
X"ee3f83e0",
X"80085583",
X"e0800876",
X"25883883",
X"e080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583e2e6",
X"347483e2",
X"e734800b",
X"83e2e834",
X"ff800b83",
X"e2e93478",
X"519bc13f",
X"83e2f333",
X"83e08008",
X"0755819f",
X"3983e2e4",
X"3383e2e5",
X"3371882b",
X"07565c74",
X"83ffff2e",
X"09810680",
X"e838fe80",
X"0b83e38c",
X"0c810b83",
X"e2f40cff",
X"0b83e2e4",
X"34ff0b83",
X"e2e53478",
X"519aec3f",
X"83e08008",
X"83e3940c",
X"83e08008",
X"5583e080",
X"08802588",
X"3883e080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"e2e63474",
X"83e2e734",
X"800b83e2",
X"e834ff80",
X"0b83e2e9",
X"34810b83",
X"e2f334a4",
X"39748596",
X"2e098106",
X"81893877",
X"83e38c0c",
X"78519aa0",
X"3f83e2f3",
X"3383e080",
X"08075574",
X"83e2f334",
X"83e2f333",
X"81065574",
X"802e8a38",
X"76840770",
X"81ff0658",
X"5583e2e8",
X"3383e2e9",
X"3371882b",
X"07565674",
X"81802e09",
X"8106a138",
X"83e2e633",
X"83e2e733",
X"71882b07",
X"565cad80",
X"75278738",
X"76820755",
X"94397681",
X"07558e39",
X"7482802e",
X"0981068c",
X"38768307",
X"557481ff",
X"06578739",
X"7481ff26",
X"8a387883",
X"e2fc1c0c",
X"767a348e",
X"3d0d0480",
X"3d0d7284",
X"2983e2fc",
X"05700883",
X"e0800c51",
X"823d0d04",
X"fe3d0d80",
X"0b83e2e0",
X"0c800b83",
X"e2dc0cff",
X"0b83e0d8",
X"0ca80b83",
X"e2f80cae",
X"518cb43f",
X"800b83e2",
X"fc545280",
X"73708405",
X"550c8112",
X"5271842e",
X"098106ef",
X"38843d0d",
X"04fe3d0d",
X"74028405",
X"96052253",
X"5371802e",
X"96387270",
X"81055433",
X"518cd33f",
X"ff127083",
X"ffff0651",
X"52e73984",
X"3d0d04fe",
X"3d0d0292",
X"05225382",
X"ac51dda8",
X"3f80c351",
X"8cb03f81",
X"9651dd9c",
X"3f725283",
X"e0dc51ff",
X"b43f7252",
X"83e0dc51",
X"f8c93f83",
X"e0800881",
X"ff06518c",
X"8d3f843d",
X"0d04ffb1",
X"3d0d80d1",
X"3df80551",
X"f8f33f83",
X"e2e00881",
X"0583e2e0",
X"0c80cf3d",
X"33cf1170",
X"81ff0651",
X"56567483",
X"2688dc38",
X"758f06ff",
X"05567583",
X"e0d8082e",
X"9b387583",
X"26963875",
X"83e0d80c",
X"75842983",
X"e2fc0570",
X"08535575",
X"51fa843f",
X"80762488",
X"b8387584",
X"2983e2fc",
X"05557408",
X"802e88a9",
X"3883e0d8",
X"08842983",
X"e2fc0570",
X"08028805",
X"82b90533",
X"525b5574",
X"80d22e84",
X"a4387480",
X"d2249038",
X"74bf2e9c",
X"387480d0",
X"2e81d638",
X"87e83974",
X"80d32e80",
X"d4387480",
X"d72e81c5",
X"3887d739",
X"0282bb05",
X"3370882b",
X"81fe8006",
X"02880582",
X"ba053371",
X"05515656",
X"8b8a3f80",
X"c1518abe",
X"3ff6c03f",
X"860b83e0",
X"dc348152",
X"83e0dc51",
X"8bf93f81",
X"51fde43f",
X"74893886",
X"0b83e2f8",
X"0c8739a8",
X"0b83e2f8",
X"0c8ad93f",
X"80c1518a",
X"8d3ff68f",
X"3f900b83",
X"e2f33381",
X"06565674",
X"802e8338",
X"985683e2",
X"e83383e2",
X"e9337188",
X"2b075659",
X"7481802e",
X"0981069c",
X"3883e2e6",
X"3383e2e7",
X"3371882b",
X"075657ad",
X"8075278c",
X"38758180",
X"07568539",
X"75a00756",
X"7583e0dc",
X"34ff0b83",
X"e0dd34e0",
X"0b83e0de",
X"34800b83",
X"e0df3484",
X"5283e0dc",
X"518af03f",
X"84518690",
X"390282bb",
X"05337088",
X"2b81fe80",
X"06028805",
X"82ba0533",
X"71055156",
X"5989c93f",
X"795194dc",
X"3f83e080",
X"08802e8a",
X"3880ce51",
X"88f03f85",
X"e23980c1",
X"5188e73f",
X"89ef3f87",
X"f33f83e3",
X"8c085883",
X"75259b38",
X"83e2e833",
X"83e2e933",
X"71882b07",
X"fc177129",
X"7a058380",
X"055a5157",
X"8d397481",
X"802918ff",
X"80055881",
X"80578056",
X"76762e92",
X"3888c63f",
X"83e08008",
X"83e0dc17",
X"34811656",
X"eb3988b5",
X"3f83e080",
X"0881ff06",
X"775383e0",
X"dc5256f4",
X"b63f83e0",
X"800881ff",
X"06557575",
X"2e098106",
X"81843888",
X"b73f80c1",
X"5187eb3f",
X"88f33f77",
X"52795193",
X"843f805e",
X"80d13dfd",
X"f4055476",
X"5383e0dc",
X"52795191",
X"983f0282",
X"b9053355",
X"81587480",
X"d72e0981",
X"06bc3880",
X"d13dfdf0",
X"05547653",
X"8f3d7053",
X"7a525992",
X"9f3f8056",
X"76762ea2",
X"38751983",
X"e0dc1733",
X"71337072",
X"32703070",
X"80257030",
X"7e06811d",
X"5d5e5151",
X"51525b55",
X"db3982ac",
X"51d7ed3f",
X"77802e86",
X"3880c351",
X"843980ce",
X"5186eb3f",
X"87f33f85",
X"f73f83da",
X"390282bb",
X"05337088",
X"2b81fe80",
X"06028805",
X"82ba0533",
X"59780559",
X"5680705d",
X"5987893f",
X"80c15186",
X"bd3f83e2",
X"f408792e",
X"82db3883",
X"e3940880",
X"fc055580",
X"fd527451",
X"b5c83f83",
X"e080085b",
X"778224b2",
X"38ff1870",
X"872b83ff",
X"ff800680",
X"f7840583",
X"e0dc5957",
X"55818055",
X"75708105",
X"57337770",
X"81055934",
X"ff157081",
X"ff065155",
X"74ea3882",
X"8a397782",
X"e82e81aa",
X"387782e9",
X"2e098106",
X"81b13880",
X"f5bc518c",
X"d43f7858",
X"77873270",
X"30707207",
X"80257a8a",
X"32703070",
X"72078025",
X"73075354",
X"5a515755",
X"75802e97",
X"38787826",
X"9238a00b",
X"83e0dc1a",
X"34811970",
X"81ff065a",
X"55eb3981",
X"187081ff",
X"0659558a",
X"7827ffbc",
X"388f5883",
X"e0d71833",
X"83e0dc19",
X"34ff1870",
X"81ff0659",
X"55778426",
X"ea389058",
X"800b83e0",
X"dc193481",
X"187081ff",
X"0670982b",
X"52595574",
X"8025e938",
X"80c6557a",
X"858f2484",
X"3880c255",
X"7483e0dc",
X"3480f10b",
X"83e0df34",
X"810b83e0",
X"e0347a83",
X"e0dd347a",
X"882c5574",
X"83e0de34",
X"80c93982",
X"f0782580",
X"c2387780",
X"fd29fd97",
X"d3055279",
X"518fb63f",
X"80d13dfd",
X"ec055480",
X"fd5383e0",
X"dc527951",
X"8ef63f7b",
X"81195956",
X"7580fc24",
X"83387858",
X"77882c55",
X"7483e1d9",
X"347783e1",
X"da347583",
X"e1db3481",
X"805980ca",
X"3983e38c",
X"08578378",
X"259b3883",
X"e2e83383",
X"e2e93371",
X"882b07fc",
X"1a712979",
X"05838005",
X"5951598d",
X"39778180",
X"2917ff80",
X"05578180",
X"59765279",
X"518ec63f",
X"80d13dfd",
X"ec055478",
X"5383e0dc",
X"5279518e",
X"873f7851",
X"f6c93f84",
X"943f8298",
X"3f8b3983",
X"e2dc0881",
X"0583e2dc",
X"0c80d13d",
X"0d04f6ea",
X"3fde853f",
X"f939fc3d",
X"0d767871",
X"842983e2",
X"fc057008",
X"51535353",
X"709e3880",
X"ce723480",
X"cf0b8113",
X"3480ce0b",
X"82133480",
X"c50b8313",
X"34708413",
X"3480e739",
X"83e39013",
X"335480d2",
X"72347382",
X"2a708106",
X"515180cf",
X"53708438",
X"80d75372",
X"811334a0",
X"0b821334",
X"73830651",
X"70812e9e",
X"38708124",
X"88387080",
X"2e8f389f",
X"3970822e",
X"92387083",
X"2e923893",
X"3980d855",
X"8e3980d3",
X"55893980",
X"cd558439",
X"80c45574",
X"83133480",
X"c40b8413",
X"34800b85",
X"1334863d",
X"0d04fe3d",
X"0d80f69c",
X"08703370",
X"81ff0670",
X"842a8132",
X"81065551",
X"52537180",
X"2e8c38a8",
X"733480f6",
X"9c0851b8",
X"71347183",
X"e0800c84",
X"3d0d04fe",
X"3d0d80f6",
X"9c087033",
X"7081ff06",
X"70852a81",
X"32810655",
X"51525371",
X"802e8c38",
X"98733480",
X"f69c0851",
X"b8713471",
X"83e0800c",
X"843d0d04",
X"803d0d80",
X"f6980851",
X"93713480",
X"f6a40851",
X"ff713482",
X"3d0d04fe",
X"3d0d0293",
X"053380f6",
X"98085353",
X"8072348a",
X"51d1b53f",
X"d33f80f6",
X"a8085280",
X"f8723480",
X"f6c00852",
X"807234fa",
X"1380f6c8",
X"08535372",
X"723480f6",
X"b0085280",
X"723480f6",
X"b8085272",
X"723480f6",
X"9c085280",
X"723480f6",
X"9c0852b8",
X"7234843d",
X"0d04ff3d",
X"0d028f05",
X"3380f6a0",
X"08525271",
X"7134fe9e",
X"3f83e080",
X"08802ef6",
X"38833d0d",
X"04803d0d",
X"8439daf0",
X"3ffeb83f",
X"83e08008",
X"802ef338",
X"80f6a008",
X"70337081",
X"ff0683e0",
X"800c5151",
X"823d0d04",
X"803d0d80",
X"f6980851",
X"a3713480",
X"f6a40851",
X"ff713480",
X"f69c0851",
X"a8713480",
X"f69c0851",
X"b8713482",
X"3d0d0480",
X"3d0d80f6",
X"98087033",
X"7081c006",
X"70307080",
X"2583e080",
X"0c515151",
X"51823d0d",
X"04ff3d0d",
X"80f69c08",
X"70337081",
X"ff067083",
X"2a813270",
X"81065151",
X"51525270",
X"802ee538",
X"b0723480",
X"f69c0851",
X"b8713483",
X"3d0d0480",
X"3d0d80f6",
X"d4087008",
X"810683e0",
X"800c5182",
X"3d0d04fd",
X"3d0d7577",
X"54548073",
X"25943873",
X"70810555",
X"335280f5",
X"c451859d",
X"3fff1353",
X"e939853d",
X"0d04f63d",
X"0d7c7e60",
X"625a5d5b",
X"56805981",
X"55853974",
X"7a295574",
X"527551ad",
X"993f83e0",
X"80087a27",
X"ee387480",
X"2e80dd38",
X"74527551",
X"ad843f83",
X"e0800875",
X"53765254",
X"adab3f83",
X"e080087a",
X"53755256",
X"acec3f83",
X"e0800879",
X"30707b07",
X"9f2a7077",
X"80240751",
X"51545572",
X"873883e0",
X"8008c538",
X"768118b0",
X"16555858",
X"8974258b",
X"38b71453",
X"7a853880",
X"d7145372",
X"78348119",
X"59ff9f39",
X"8077348c",
X"3d0d04f7",
X"3d0d7b7d",
X"7f620290",
X"05bb0533",
X"5759565a",
X"5ab05872",
X"8338a058",
X"75707081",
X"05523371",
X"59545590",
X"39807425",
X"8e38ff14",
X"77708105",
X"59335454",
X"72ef3873",
X"ff155553",
X"80732589",
X"38775279",
X"51782def",
X"39753375",
X"57537280",
X"2e903872",
X"52795178",
X"2d757081",
X"05573353",
X"ed398b3d",
X"0d04ee3d",
X"0d646669",
X"69707081",
X"0552335b",
X"4a5c5e5e",
X"76802e82",
X"f93876a5",
X"2e098106",
X"82e03880",
X"70416770",
X"70810552",
X"33714a59",
X"575f76b0",
X"2e098106",
X"8c387570",
X"81055733",
X"76485781",
X"5fd01756",
X"75892680",
X"da387667",
X"5c59805c",
X"9339778a",
X"2480c338",
X"7b8a2918",
X"7b708105",
X"5d335a5c",
X"d0197081",
X"ff065858",
X"897727a4",
X"38ff9f19",
X"7081ff06",
X"ffa91b5a",
X"51568576",
X"279238ff",
X"bf197081",
X"ff065156",
X"7585268a",
X"38c91958",
X"778025ff",
X"b9387a47",
X"7b407881",
X"ff065776",
X"80e42e80",
X"e5387680",
X"e424a738",
X"7680d82e",
X"81863876",
X"80d82490",
X"3876802e",
X"81cc3876",
X"a52e81b6",
X"3881b939",
X"7680e32e",
X"818c3881",
X"af397680",
X"f52e9b38",
X"7680f524",
X"8b387680",
X"f32e8181",
X"38819939",
X"7680f82e",
X"80ca3881",
X"8f39913d",
X"70555780",
X"538a5279",
X"841b7108",
X"535b56fc",
X"813f7655",
X"ab397984",
X"1b710894",
X"3d705b5b",
X"525b5675",
X"80258c38",
X"753056ad",
X"78340280",
X"c1055776",
X"5480538a",
X"527551fb",
X"d53f7755",
X"7e54b839",
X"913d7055",
X"7780d832",
X"70307080",
X"25565158",
X"56905279",
X"841b7108",
X"535b57fb",
X"b13f7555",
X"db397984",
X"1b831233",
X"545b5698",
X"3979841b",
X"7108575b",
X"5680547f",
X"537c527d",
X"51fc9c3f",
X"87397652",
X"7d517c2d",
X"66703358",
X"810547fd",
X"8339943d",
X"0d047283",
X"e0900c71",
X"83e0940c",
X"04fb3d0d",
X"883d7070",
X"84055208",
X"57547553",
X"83e09008",
X"5283e094",
X"0851fcc6",
X"3f873d0d",
X"04ff3d0d",
X"73700853",
X"51029305",
X"33723470",
X"08810571",
X"0c833d0d",
X"04fc3d0d",
X"873d8811",
X"55785480",
X"c2b15351",
X"fc983f80",
X"52873d51",
X"d03f863d",
X"0d04803d",
X"0d725170",
X"802e8338",
X"81517083",
X"e0800c82",
X"3d0d04ff",
X"3d0d028f",
X"05337030",
X"709f2a83",
X"e0800c52",
X"52833d0d",
X"04fd3d0d",
X"75705254",
X"a4e73f83",
X"e0800814",
X"5372742e",
X"9238ff13",
X"70335353",
X"71af2e09",
X"8106ee38",
X"81135372",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"77705354",
X"54c73f83",
X"e0800873",
X"2ea13883",
X"e0800873",
X"3152ff12",
X"5271ff2e",
X"8f387270",
X"81055433",
X"74708105",
X"5634eb39",
X"ff145480",
X"7434853d",
X"0d04803d",
X"0d7251ff",
X"903f823d",
X"0d047183",
X"e0800c04",
X"803d0d72",
X"51807134",
X"810bbc12",
X"0c800b80",
X"c0120c82",
X"3d0d0480",
X"0b83e5bc",
X"08248a38",
X"a5d83fff",
X"0b83e5bc",
X"0c800b83",
X"e0800c04",
X"ff3d0d73",
X"5283e398",
X"08722e8d",
X"38d93f71",
X"5196de3f",
X"7183e398",
X"0c833d0d",
X"04f43d0d",
X"7e60625c",
X"5a558154",
X"bc150881",
X"92387451",
X"cf3f7958",
X"807a2580",
X"f73883e5",
X"ec087089",
X"2a5783ff",
X"06788480",
X"72315656",
X"57737825",
X"83387355",
X"7583e5bc",
X"082e8438",
X"ff893f83",
X"e5bc0880",
X"25a63875",
X"892b5199",
X"ca3f83e5",
X"ec088f3d",
X"fc11555c",
X"548152f8",
X"1b5197af",
X"3f761483",
X"e5ec0c75",
X"83e5bc0c",
X"74537652",
X"7851a3eb",
X"3f83e080",
X"0883e5ec",
X"081683e5",
X"ec0c7876",
X"31761b5b",
X"59567780",
X"24ff8b38",
X"617a710c",
X"547551fc",
X"f13f83e0",
X"80085473",
X"83e0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"9a3f7651",
X"feae3f86",
X"3dfc0553",
X"02a20522",
X"52775196",
X"ce3f7986",
X"3d22710c",
X"5483e080",
X"0851fcba",
X"3f863d0d",
X"04fd3d0d",
X"7683e5bc",
X"08535380",
X"72248938",
X"71732e84",
X"38fddc3f",
X"7551fdf0",
X"3f725198",
X"a23f7351",
X"fc903f85",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"e0800c51",
X"823d0d04",
X"80c40b83",
X"e0800c04",
X"fd3d0d75",
X"77715470",
X"535553a0",
X"d43f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfd803f",
X"73519485",
X"3f7383e3",
X"980c83e0",
X"800851fb",
X"b13f853d",
X"0d04fd3d",
X"0d757755",
X"53fce03f",
X"72802ea5",
X"38bc1308",
X"5273519f",
X"ea3f83e0",
X"80088f38",
X"77527251",
X"ffa63f83",
X"e0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83e0800c",
X"853d0d04",
X"ff3d0dff",
X"0b83e5bc",
X"0c7383e3",
X"9c0c7483",
X"e5b80ca0",
X"d03f83e0",
X"800881ff",
X"06527180",
X"2e883871",
X"51fadc3f",
X"903983e5",
X"d4518f82",
X"3f83e080",
X"0851fab6",
X"3f833d0d",
X"04fa3d0d",
X"787a82c4",
X"120882c4",
X"12087072",
X"24595656",
X"57577373",
X"2e098106",
X"913880c0",
X"165280c0",
X"17519de2",
X"3f83e080",
X"08557483",
X"e0800c88",
X"3d0d04f6",
X"3d0d7c5b",
X"807b715c",
X"54577a77",
X"2e8c3881",
X"1a82cc14",
X"08545a72",
X"f6388059",
X"80d9397a",
X"54815780",
X"707b7b31",
X"5a5755ff",
X"18537473",
X"2580c138",
X"82cc1408",
X"527351ff",
X"8c3f800b",
X"83e08008",
X"25a13882",
X"cc140882",
X"cc110882",
X"cc160c74",
X"82cc120c",
X"5375802e",
X"86387282",
X"cc170c72",
X"54805773",
X"82cc1508",
X"81175755",
X"56ffb839",
X"81195980",
X"0bff1b54",
X"54787325",
X"83388154",
X"76813270",
X"75065153",
X"72ff9038",
X"8c3d0d04",
X"f73d0d7b",
X"7d5a5a82",
X"d05283e5",
X"b80851a0",
X"a13f83e0",
X"800857fa",
X"8a3f7952",
X"83e5c051",
X"96c73f83",
X"e0800853",
X"805483e0",
X"8008742e",
X"09810682",
X"833883e3",
X"9c080b0b",
X"80f58853",
X"7052559d",
X"a03f0b0b",
X"80f58852",
X"80c01551",
X"9d933f74",
X"bc160c72",
X"82c0160c",
X"810b82c4",
X"160c810b",
X"82c8160c",
X"ff177357",
X"57819739",
X"83e3a833",
X"70822a70",
X"81065154",
X"54728186",
X"3873812a",
X"81065877",
X"80fc3876",
X"802e8190",
X"3882d015",
X"ff187584",
X"2a810682",
X"c4130c83",
X"e3a83381",
X"0682c813",
X"0c7b5471",
X"5358569c",
X"b43f7551",
X"9ccb3f83",
X"e0800816",
X"53af7370",
X"81055534",
X"72bc170c",
X"83e3a952",
X"72519c95",
X"3f83e3a0",
X"0882c017",
X"0c83e3b6",
X"52839015",
X"519c823f",
X"7782cc17",
X"0c78802e",
X"8d387551",
X"782d83e0",
X"8008802e",
X"8d387480",
X"2e863875",
X"82cc160c",
X"755583e3",
X"a05283e5",
X"c05195e7",
X"3f83e080",
X"088a3883",
X"e3a93353",
X"72fed138",
X"800b82cc",
X"170c7880",
X"2e893883",
X"e39c0851",
X"fcb93f83",
X"e39c0854",
X"7383e080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb63f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f6b9",
X"3f83e080",
X"08745387",
X"3d705355",
X"55f6d93f",
X"f7b93f73",
X"51d33f63",
X"53745283",
X"e0800851",
X"fac03f92",
X"3d0d0471",
X"83e0800c",
X"0480c012",
X"83e0800c",
X"04803d0d",
X"7282c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"e0800c51",
X"823d0d04",
X"f63d0d7c",
X"83e09808",
X"59598179",
X"2782a938",
X"78881908",
X"2782a138",
X"77335675",
X"822e819b",
X"38758224",
X"89387581",
X"2e8d3882",
X"8b397583",
X"2e81b738",
X"82823978",
X"83ffff06",
X"70812a11",
X"7083ffff",
X"067083ff",
X"0671892a",
X"903d5f52",
X"5a515155",
X"7683ff2e",
X"8e388254",
X"76538c18",
X"08155279",
X"51a93975",
X"5476538c",
X"18081552",
X"79519abe",
X"3f83e080",
X"0881bd38",
X"755483e0",
X"8008538c",
X"18081581",
X"05528c3d",
X"fd05519a",
X"a13f83e0",
X"800881a0",
X"3802a905",
X"338c3d33",
X"71882b07",
X"7a810671",
X"842a5357",
X"58567486",
X"38769fff",
X"06567555",
X"81803975",
X"54781083",
X"fe065378",
X"882a8c19",
X"0805528c",
X"3dfc0551",
X"99e03f83",
X"e0800880",
X"df3802a9",
X"05338c3d",
X"3371882b",
X"07565780",
X"d1398454",
X"78822b83",
X"fc065378",
X"872a8c19",
X"0805528c",
X"3dfc0551",
X"99b03f83",
X"e08008b0",
X"3802ab05",
X"33028405",
X"aa053371",
X"982b7190",
X"2b07028c",
X"05a90533",
X"70882b72",
X"07903d33",
X"7180ffff",
X"fe800607",
X"51525357",
X"58568339",
X"81557483",
X"e0800c8c",
X"3d0d04fb",
X"3d0d83e0",
X"9808fe19",
X"881208fe",
X"05555654",
X"80567473",
X"278d3882",
X"14337571",
X"29941608",
X"05575375",
X"83e0800c",
X"873d0d04",
X"fc3d0d76",
X"83e09808",
X"55558075",
X"23881508",
X"5372812e",
X"88388814",
X"08732685",
X"388152b2",
X"39729038",
X"73335271",
X"832e0981",
X"06853890",
X"14085372",
X"8c160c72",
X"802e8d38",
X"7251ff93",
X"3f83e080",
X"08528539",
X"90140852",
X"7190160c",
X"80527183",
X"e0800c86",
X"3d0d04fa",
X"3d0d7883",
X"e0980871",
X"22810570",
X"83ffff06",
X"57545755",
X"73802e88",
X"38901508",
X"53728638",
X"835280e7",
X"39738f06",
X"527180da",
X"38811390",
X"160c8c15",
X"08537290",
X"38830b84",
X"17225752",
X"73762780",
X"c638bf39",
X"821633ff",
X"0574842a",
X"065271b2",
X"387251fb",
X"db3f8152",
X"7183e080",
X"0827a838",
X"835283e0",
X"80088817",
X"08279c38",
X"83e08008",
X"8c160c83",
X"e0800851",
X"fdf93f83",
X"e0800890",
X"160c7375",
X"23805271",
X"83e0800c",
X"883d0d04",
X"f23d0d60",
X"6264585d",
X"5b753355",
X"74a02e09",
X"81068838",
X"81167044",
X"56ef3962",
X"70335656",
X"74af2e09",
X"81068438",
X"81164380",
X"0b881c0c",
X"62703351",
X"5574a026",
X"91387a51",
X"fdd23f83",
X"e0800856",
X"807c3483",
X"a839933d",
X"841c0870",
X"585a5f8a",
X"55a07670",
X"81055834",
X"ff155574",
X"ff2e0981",
X"06ef3880",
X"70595d88",
X"7f085f5a",
X"7c811e70",
X"81ff0660",
X"13703370",
X"af327030",
X"a0732771",
X"80250751",
X"51525b53",
X"5f575574",
X"80d83876",
X"ae2e0981",
X"06833881",
X"55777a27",
X"75075574",
X"802e9f38",
X"79883270",
X"3078ae32",
X"70307073",
X"079f2a53",
X"51575156",
X"75ac3888",
X"588b5aff",
X"ab39ff9f",
X"17557499",
X"268938e0",
X"177081ff",
X"06585577",
X"81197081",
X"ff06721c",
X"535a5755",
X"767534ff",
X"87397c1e",
X"7f0c8055",
X"76a02683",
X"38815574",
X"8b1a347a",
X"51fc913f",
X"83e08008",
X"80f538a0",
X"547a2270",
X"852b83e0",
X"06545590",
X"1b08527b",
X"5194b73f",
X"83e08008",
X"5783e080",
X"08818238",
X"7b335574",
X"802e80f5",
X"388b1c33",
X"70832a70",
X"81065156",
X"5674b438",
X"8b7c841d",
X"0883e080",
X"08595b5b",
X"58ff1858",
X"77ff2e9a",
X"38797081",
X"055b3379",
X"7081055b",
X"33717131",
X"52565675",
X"802ee238",
X"86397580",
X"2ebc387a",
X"51fbf43f",
X"ff863983",
X"e0800856",
X"83e08008",
X"802ea938",
X"83e08008",
X"832e0981",
X"0680de38",
X"841b088b",
X"11335155",
X"7480d238",
X"845680cd",
X"398356ec",
X"39815680",
X"c4397656",
X"841b088b",
X"11335155",
X"74b7388b",
X"1c337084",
X"2a708106",
X"51565774",
X"802ed538",
X"951c3394",
X"1d337198",
X"2b71902b",
X"079b1f33",
X"7f9a0533",
X"71882b07",
X"72077f88",
X"050c5a58",
X"5658fcda",
X"397583e0",
X"800c903d",
X"0d04f83d",
X"0d7a7c59",
X"57825483",
X"fe537752",
X"765192c6",
X"3f835683",
X"e0800880",
X"ec388117",
X"33773371",
X"882b0756",
X"56825674",
X"82d4d52e",
X"09810680",
X"d4387554",
X"b6537752",
X"7651929a",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"ac388254",
X"80d25377",
X"52765191",
X"f13f83e0",
X"80089838",
X"81173377",
X"3371882b",
X"0783e080",
X"08525656",
X"748182c6",
X"2e833881",
X"567583e0",
X"800c8a3d",
X"0d04ec3d",
X"0d665980",
X"0b83e098",
X"0c785678",
X"802e83e8",
X"38919e3f",
X"83e08008",
X"81065582",
X"567483d8",
X"38747553",
X"8e3d7053",
X"5858fec2",
X"3f83e080",
X"0881ff06",
X"5675812e",
X"09810680",
X"d4389054",
X"83be5374",
X"52765190",
X"fd3f83e0",
X"800880c9",
X"388e3d33",
X"5574802e",
X"80c93802",
X"bb053302",
X"8405ba05",
X"3371982b",
X"71902b07",
X"028c05b9",
X"05337088",
X"2b720794",
X"3d337107",
X"70587c57",
X"54525d57",
X"5956fde6",
X"3f83e080",
X"0881ff06",
X"5675832e",
X"09810686",
X"38815682",
X"db397580",
X"2e863887",
X"5682d139",
X"a4548d53",
X"77527651",
X"90943f81",
X"5683e080",
X"0882bd38",
X"02ba0533",
X"028405b9",
X"05337188",
X"2b07585c",
X"76ab3802",
X"80ca0533",
X"02840580",
X"c9053371",
X"982b7190",
X"2b07963d",
X"3370882b",
X"72070294",
X"0580c705",
X"33710754",
X"525d5758",
X"5602b305",
X"33777129",
X"028805b2",
X"0533028c",
X"05b10533",
X"71882b07",
X"701c708c",
X"1f0c5e59",
X"57585c8d",
X"3d33821a",
X"3402b505",
X"338f3d33",
X"71882b07",
X"595b7784",
X"1a2302b7",
X"05330284",
X"05b60533",
X"71882b07",
X"565b74ab",
X"380280c6",
X"05330284",
X"0580c505",
X"3371982b",
X"71902b07",
X"953d3370",
X"882b7207",
X"02940580",
X"c3053371",
X"07515253",
X"575d5b74",
X"76317731",
X"78842a8f",
X"3d335471",
X"71315356",
X"5690833f",
X"83e08008",
X"82057088",
X"1b0c709f",
X"f6268105",
X"575583ff",
X"f6752783",
X"38835675",
X"79347583",
X"2e098106",
X"af380280",
X"d2053302",
X"840580d1",
X"05337198",
X"2b71902b",
X"07983d33",
X"70882b72",
X"07029405",
X"80cf0533",
X"7107901f",
X"0c525d57",
X"59568639",
X"761a901a",
X"0c841922",
X"8c1a0818",
X"71842a05",
X"941b0c5c",
X"800b811a",
X"347883e0",
X"980c8056",
X"7583e080",
X"0c963d0d",
X"04e93d0d",
X"83e09808",
X"56865475",
X"802e81a6",
X"38800b81",
X"1734993d",
X"e011466a",
X"54c01153",
X"ec0551f6",
X"cf3f83e0",
X"80085483",
X"e0800881",
X"8538893d",
X"33547380",
X"2e933802",
X"ab053370",
X"842a7081",
X"06515555",
X"73802e86",
X"38835480",
X"e53902b5",
X"05338f3d",
X"3371982b",
X"71902b07",
X"028c05bb",
X"05330290",
X"05ba0533",
X"71882b07",
X"7207a01b",
X"0c029005",
X"bf053302",
X"9405be05",
X"3371982b",
X"71902b07",
X"029c05bd",
X"05337088",
X"2b720799",
X"3d337107",
X"7f9c050c",
X"5283e080",
X"08981f0c",
X"565a5252",
X"53575957",
X"810b8117",
X"3483e080",
X"08547383",
X"e0800c99",
X"3d0d04f5",
X"3d0d7d60",
X"028805ba",
X"05227283",
X"e098085b",
X"5d5a5c5c",
X"807b2386",
X"5676802e",
X"81e03881",
X"17338106",
X"55855674",
X"802e81d2",
X"389c1708",
X"98180831",
X"55747827",
X"87387483",
X"ffff0658",
X"77802e81",
X"ae389817",
X"087083ff",
X"06565674",
X"80ca3882",
X"1733ff05",
X"76892a06",
X"7081ff06",
X"5a5578a0",
X"38758738",
X"a0170855",
X"8d39a417",
X"0851efe0",
X"3f83e080",
X"08558175",
X"2780f838",
X"74a4180c",
X"a4170851",
X"f28d3f83",
X"e0800880",
X"2e80e438",
X"83e08008",
X"19a8180c",
X"98170883",
X"ff068480",
X"71317083",
X"ffff0658",
X"51557776",
X"27833877",
X"56755498",
X"170883ff",
X"0653a817",
X"08527955",
X"7b83387b",
X"5574518a",
X"b93f83e0",
X"8008a438",
X"98170816",
X"98180c75",
X"1a787731",
X"7083ffff",
X"067d2279",
X"05525a56",
X"5a747b23",
X"fece3980",
X"56883980",
X"0b811834",
X"81567583",
X"e0800c8d",
X"3d0d04fa",
X"3d0d7883",
X"e0980855",
X"56865573",
X"802e81dc",
X"38811433",
X"81065385",
X"5572802e",
X"81ce389c",
X"14085372",
X"76278338",
X"72569814",
X"0857800b",
X"98150c75",
X"802e81a9",
X"38821433",
X"70892b56",
X"5376802e",
X"b5387452",
X"ff16518a",
X"f13f83e0",
X"8008ff18",
X"76547053",
X"58538ae2",
X"3f83e080",
X"08732696",
X"38743070",
X"78067098",
X"170c7771",
X"31a41708",
X"52585153",
X"8939a014",
X"0870a416",
X"0c537476",
X"27b43872",
X"51edc13f",
X"83e08008",
X"53810b83",
X"e0800827",
X"80cb3883",
X"e0800888",
X"15082780",
X"c03883e0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c9399814",
X"08167098",
X"160c7352",
X"56efc83f",
X"83e08008",
X"802e9638",
X"821433ff",
X"0576892a",
X"0683e080",
X"0805a815",
X"0c805588",
X"39800b81",
X"15348155",
X"7483e080",
X"0c883d0d",
X"04ee3d0d",
X"64568655",
X"83e09808",
X"802e80f6",
X"38943df4",
X"1184180c",
X"6654d405",
X"527551f1",
X"973f83e0",
X"80085583",
X"e0800880",
X"cf38893d",
X"33547380",
X"2ebc3802",
X"ab053370",
X"842a7081",
X"06515555",
X"84557380",
X"2ebc3802",
X"b505338f",
X"3d337198",
X"2b71902b",
X"07028c05",
X"bb053302",
X"9005ba05",
X"3371882b",
X"07720788",
X"1b0c5357",
X"59577551",
X"eed23f83",
X"e0800855",
X"74832e09",
X"81068338",
X"84557483",
X"e0800c94",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405d",
X"865683e0",
X"9808802e",
X"849b389e",
X"3df40584",
X"1e0c7e98",
X"387c51ee",
X"973f83e0",
X"80085684",
X"84398141",
X"82803983",
X"4181fb39",
X"933d7f96",
X"05415980",
X"7f829505",
X"5f567560",
X"81ff0534",
X"8341901d",
X"08762e81",
X"dd38a054",
X"7c227085",
X"2b83e006",
X"5458901d",
X"08527851",
X"86943f83",
X"e0800841",
X"83e08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"e8387b81",
X"bf065574",
X"8f2480dd",
X"389a1933",
X"557480d5",
X"389c1933",
X"5574802e",
X"80cb38f3",
X"1e70585e",
X"8156758b",
X"2e098106",
X"85388e56",
X"8b39759a",
X"2e098106",
X"83389c56",
X"75197070",
X"81055233",
X"7133811a",
X"821a5f5b",
X"525b5574",
X"86387977",
X"34853980",
X"df773477",
X"7b57577a",
X"a02e0981",
X"06c03881",
X"567b81e5",
X"32703070",
X"9f2a5151",
X"557bae2e",
X"93387480",
X"2e8e3861",
X"832a7081",
X"06515574",
X"802e9738",
X"7c51ecf7",
X"3f83e080",
X"084183e0",
X"80088738",
X"901d08fe",
X"a5388060",
X"3475802e",
X"88387d52",
X"7f5183b1",
X"3f60802e",
X"8638800b",
X"901e0c60",
X"5660832e",
X"09810688",
X"38800b90",
X"1e0c8539",
X"6081d238",
X"891f5790",
X"1d08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347c51ea",
X"fe3f83e0",
X"80085683",
X"e0800883",
X"2e098106",
X"8838800b",
X"901e0c80",
X"56961f33",
X"55748a38",
X"891f5296",
X"1f5181b1",
X"3f7583e0",
X"800c9e3d",
X"0d04fd3d",
X"0d757753",
X"54733351",
X"70893871",
X"33517080",
X"2ea13873",
X"33723352",
X"53727127",
X"8538ff51",
X"94397073",
X"27853881",
X"518b3981",
X"14811353",
X"54d33980",
X"517083e0",
X"800c853d",
X"0d04fd3d",
X"0d757754",
X"54723370",
X"81ff0652",
X"5270802e",
X"a3387181",
X"ff068114",
X"ffbf1253",
X"54527099",
X"268938a0",
X"127081ff",
X"06535171",
X"74708105",
X"5634d239",
X"80743485",
X"3d0d04ff",
X"bd3d0d80",
X"c63d0852",
X"a53d7052",
X"54ffb33f",
X"80c73d08",
X"52853d70",
X"5253ffa6",
X"3f725273",
X"51fedf3f",
X"80c53d0d",
X"04fe3d0d",
X"74765353",
X"71708105",
X"53335170",
X"73708105",
X"553470f0",
X"38843d0d",
X"04fe3d0d",
X"74528072",
X"33525370",
X"732e8d38",
X"81128114",
X"71335354",
X"5270f538",
X"7283e080",
X"0c843d0d",
X"04fd3d0d",
X"75547383",
X"e684082e",
X"a83880f6",
X"e4087481",
X"800a0771",
X"0c80f6f4",
X"08535371",
X"08517080",
X"2ef93880",
X"730c7108",
X"5170fb38",
X"7383e684",
X"0c853d0d",
X"04ff0b83",
X"e6840c81",
X"80800b83",
X"e6800c80",
X"0b83e080",
X"0c04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"9c3f7280",
X"2ea33883",
X"e6800814",
X"52713375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552da",
X"39800b83",
X"e0800c86",
X"3d0d04f7",
X"3d0d7b7d",
X"7f115855",
X"59805573",
X"762eb138",
X"83e68008",
X"8b3d5957",
X"74197033",
X"75fc0619",
X"70085d76",
X"83067b07",
X"53545451",
X"72713479",
X"720c8114",
X"81165654",
X"73762e09",
X"8106d938",
X"800b83e0",
X"800c8b3d",
X"0d04fe3d",
X"0d80f6e4",
X"0883e684",
X"0880c00a",
X"07710c80",
X"f6f40853",
X"53710851",
X"70802ef9",
X"3880730c",
X"71085170",
X"fb38843d",
X"0d0483e0",
X"8c080283",
X"e08c0cfd",
X"3d0d8053",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"83d43f83",
X"e0800870",
X"83e0800c",
X"54853d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cfd3d",
X"0d815383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"05085183",
X"a13f83e0",
X"80087083",
X"e0800c54",
X"853d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cf93d0d",
X"800b83e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"8025b938",
X"83e08c08",
X"88050830",
X"83e08c08",
X"88050c80",
X"0b83e08c",
X"08f4050c",
X"83e08c08",
X"fc05088a",
X"38810b83",
X"e08c08f4",
X"050c83e0",
X"8c08f405",
X"0883e08c",
X"08fc050c",
X"83e08c08",
X"8c050880",
X"25b93883",
X"e08c088c",
X"05083083",
X"e08c088c",
X"050c800b",
X"83e08c08",
X"f0050c83",
X"e08c08fc",
X"05088a38",
X"810b83e0",
X"8c08f005",
X"0c83e08c",
X"08f00508",
X"83e08c08",
X"fc050c80",
X"5383e08c",
X"088c0508",
X"5283e08c",
X"08880508",
X"5181df3f",
X"83e08008",
X"7083e08c",
X"08f8050c",
X"5483e08c",
X"08fc0508",
X"802e9038",
X"83e08c08",
X"f8050830",
X"83e08c08",
X"f8050c83",
X"e08c08f8",
X"05087083",
X"e0800c54",
X"893d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"800b83e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"80259938",
X"83e08c08",
X"88050830",
X"83e08c08",
X"88050c81",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"8c050880",
X"25903883",
X"e08c088c",
X"05083083",
X"e08c088c",
X"050c8153",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"bd3f83e0",
X"80087083",
X"e08c08f8",
X"050c5483",
X"e08c08fc",
X"0508802e",
X"903883e0",
X"8c08f805",
X"083083e0",
X"8c08f805",
X"0c83e08c",
X"08f80508",
X"7083e080",
X"0c54873d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cfd",
X"3d0d810b",
X"83e08c08",
X"fc050c80",
X"0b83e08c",
X"08f8050c",
X"83e08c08",
X"8c050883",
X"e08c0888",
X"050827b9",
X"3883e08c",
X"08fc0508",
X"802eae38",
X"800b83e0",
X"8c088c05",
X"0824a238",
X"83e08c08",
X"8c050810",
X"83e08c08",
X"8c050c83",
X"e08c08fc",
X"05081083",
X"e08c08fc",
X"050cffb8",
X"3983e08c",
X"08fc0508",
X"802e80e1",
X"3883e08c",
X"088c0508",
X"83e08c08",
X"88050826",
X"ad3883e0",
X"8c088805",
X"0883e08c",
X"088c0508",
X"3183e08c",
X"0888050c",
X"83e08c08",
X"f8050883",
X"e08c08fc",
X"05080783",
X"e08c08f8",
X"050c83e0",
X"8c08fc05",
X"08812a83",
X"e08c08fc",
X"050c83e0",
X"8c088c05",
X"08812a83",
X"e08c088c",
X"050cff95",
X"3983e08c",
X"08900508",
X"802e9338",
X"83e08c08",
X"88050870",
X"83e08c08",
X"f4050c51",
X"913983e0",
X"8c08f805",
X"087083e0",
X"8c08f405",
X"0c5183e0",
X"8c08f405",
X"0883e080",
X"0c853d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cff3d",
X"0d800b83",
X"e08c08fc",
X"050c83e0",
X"8c088805",
X"088106ff",
X"11700970",
X"83e08c08",
X"8c050806",
X"83e08c08",
X"fc050811",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"0508812a",
X"83e08c08",
X"88050c83",
X"e08c088c",
X"05081083",
X"e08c088c",
X"050c5151",
X"515183e0",
X"8c088805",
X"08802e84",
X"38ffab39",
X"83e08c08",
X"fc050870",
X"83e0800c",
X"51833d0d",
X"83e08c0c",
X"04fc3d0d",
X"7670797b",
X"55555555",
X"8f72278c",
X"38727507",
X"83065170",
X"802ea938",
X"ff125271",
X"ff2e9838",
X"72708105",
X"54337470",
X"81055634",
X"ff125271",
X"ff2e0981",
X"06ea3874",
X"83e0800c",
X"863d0d04",
X"74517270",
X"84055408",
X"71708405",
X"530c7270",
X"84055408",
X"71708405",
X"530c7270",
X"84055408",
X"71708405",
X"530c7270",
X"84055408",
X"71708405",
X"530cf012",
X"52718f26",
X"c9388372",
X"27953872",
X"70840554",
X"08717084",
X"05530cfc",
X"12527183",
X"26ed3870",
X"54ff8139",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"00000809",
X"00000811",
X"00000819",
X"00000821",
X"00000829",
X"00000831",
X"00000839",
X"00000841",
X"000009f0",
X"00000a31",
X"00000a53",
X"00000a71",
X"00000a71",
X"00000a71",
X"00000a71",
X"00000ae0",
X"00000b10",
X"70704740",
X"9c704268",
X"9c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"43617274",
X"72696467",
X"6520386b",
X"2073696d",
X"706c6500",
X"45786974",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"25732025",
X"73000000",
X"2e2e0000",
X"2f000000",
X"41545200",
X"58464400",
X"58455800",
X"524f4d00",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"6e616d65",
X"20000000",
X"25303278",
X"00000000",
X"00000000",
X"00000000",
X"0001d20f",
X"0001d400",
X"0001d401",
X"0001d409",
X"0001d010",
X"0001d301",
X"0001d300",
X"0001d20a",
X"0001d01b",
X"0001d016",
X"0001d019",
X"0001d018",
X"0001d017",
X"0001d01a",
X"0001d403",
X"0001d402",
X"0001d40e",
X"0004007c",
X"00040078",
X"00040074",
X"00040068",
X"00040060",
X"0004005c",
X"00040058",
X"00040054",
X"00040050",
X"0004004c",
X"00040048",
X"00040044",
X"00040040",
X"00040034",
X"00040030",
X"0004002c",
X"00040028",
X"00040024",
X"00040020",
X"0004001c",
X"00040018",
X"00040014",
X"00040010",
X"0004000c",
X"00040008",
X"00040004",
X"00040000",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
