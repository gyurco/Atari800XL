
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f6",
X"e0738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80fa",
X"980c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f2",
X"a82d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580f0bc",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80da9704",
X"f93d0d80",
X"0b83e080",
X"0c893d0d",
X"04fc3d0d",
X"76705255",
X"b3c93f83",
X"e0800815",
X"ff055473",
X"752e8e38",
X"73335372",
X"ae2e8638",
X"ff1454ef",
X"39775281",
X"1451b2e1",
X"3f83e080",
X"08307083",
X"e0800807",
X"802583e0",
X"800c5386",
X"3d0d04fc",
X"3d0d7670",
X"52559a82",
X"3f83e080",
X"08548153",
X"83e08008",
X"80c73874",
X"5199c53f",
X"83e08008",
X"0b0b80f8",
X"a05383e0",
X"80085253",
X"ff8f3f83",
X"e08008a5",
X"380b0b80",
X"f8a45272",
X"51fefe3f",
X"83e08008",
X"94380b0b",
X"80f8a852",
X"7251feed",
X"3f83e080",
X"08802e83",
X"38815473",
X"537283e0",
X"800c863d",
X"0d04fd3d",
X"0d757052",
X"54999b3f",
X"815383e0",
X"80089838",
X"735198e4",
X"3f83e0a0",
X"085283e0",
X"800851fe",
X"b43f83e0",
X"80085372",
X"83e0800c",
X"853d0d04",
X"e03d0da3",
X"3d087052",
X"5e8f893f",
X"83e08008",
X"33943d56",
X"54739438",
X"80fecc52",
X"745184c7",
X"397d5278",
X"51928c3f",
X"84d1397d",
X"518ef13f",
X"83e08008",
X"5274518e",
X"a13f83e0",
X"a8085293",
X"3d70525d",
X"94fc3f83",
X"e0800859",
X"800b83e0",
X"8008555b",
X"83e08008",
X"7b2e9438",
X"811b7452",
X"5b97fe3f",
X"83e08008",
X"5483e080",
X"08ee3880",
X"5aff7a43",
X"7a427a41",
X"5f790970",
X"9f2c7b06",
X"5b547a7a",
X"248438ff",
X"1b5af61a",
X"7009709f",
X"2c72067b",
X"ff125a5a",
X"52555580",
X"75259538",
X"765197bd",
X"3f83e080",
X"0876ff18",
X"58555773",
X"8024ed38",
X"747f2e87",
X"3880c3a1",
X"3f745f78",
X"ff1b7058",
X"5d58807a",
X"25953877",
X"5197923f",
X"83e08008",
X"76ff1858",
X"55587380",
X"24ed3880",
X"0b83e7bc",
X"0c800b83",
X"e7dc0c0b",
X"0b80f8ac",
X"518be43f",
X"81800b83",
X"e7dc0c0b",
X"0b80f8b4",
X"518bd43f",
X"a80b83e7",
X"bc0c7680",
X"2e80e838",
X"83e7bc08",
X"77793270",
X"30707207",
X"80257087",
X"2b83e7dc",
X"0c515678",
X"53565696",
X"c53f83e0",
X"8008802e",
X"8a380b0b",
X"80f8bc51",
X"8b993f76",
X"5196853f",
X"83e08008",
X"520b0b80",
X"f9c8518b",
X"863f7651",
X"968b3f83",
X"e0800883",
X"e7bc0855",
X"57757425",
X"8638a816",
X"56f73975",
X"83e7bc0c",
X"86f07624",
X"ff943887",
X"980b83e7",
X"bc0c7780",
X"2eb73877",
X"5195c13f",
X"83e08008",
X"78525595",
X"e13f0b0b",
X"80f8c454",
X"83e08008",
X"8f388739",
X"807634fd",
X"95390b0b",
X"80f8c054",
X"74537352",
X"0b0b80f8",
X"94518a9f",
X"3f80540b",
X"0b80fa94",
X"518a943f",
X"81145473",
X"a82e0981",
X"06ed3886",
X"8da051bf",
X"a03f8052",
X"903d7052",
X"5480e085",
X"3f835273",
X"5180dffd",
X"3f61802e",
X"80ff387b",
X"5473ff2e",
X"96387880",
X"2e818038",
X"785194e1",
X"3f83e080",
X"08ff1555",
X"59e73978",
X"802e80eb",
X"38785194",
X"dd3f83e0",
X"8008802e",
X"fc833878",
X"5194a53f",
X"83e08008",
X"520b0b80",
X"f89c51ac",
X"833f83e0",
X"8008a438",
X"7c51adbb",
X"3f83e080",
X"085574ff",
X"16565480",
X"7425fbee",
X"38741d70",
X"33555673",
X"af2efec8",
X"38e83978",
X"5193e33f",
X"83e08008",
X"527c51ac",
X"f23ffbce",
X"397f8829",
X"6010057a",
X"0561055a",
X"fbff39a2",
X"3d0d04fe",
X"3d0d80fd",
X"d4087033",
X"7081ff06",
X"70842a81",
X"32810655",
X"51525371",
X"802e8c38",
X"a8733480",
X"fdd40851",
X"b8713471",
X"83e0800c",
X"843d0d04",
X"fe3d0d80",
X"fdd40870",
X"337081ff",
X"0670852a",
X"81328106",
X"55515253",
X"71802e8c",
X"38987334",
X"80fdd408",
X"51b87134",
X"7183e080",
X"0c843d0d",
X"04803d0d",
X"80fdd008",
X"51937134",
X"80fddc08",
X"51ff7134",
X"823d0d04",
X"fe3d0d02",
X"93053380",
X"fdd00853",
X"53807234",
X"8a51bce9",
X"3fd33f80",
X"fde00852",
X"80f87234",
X"80fdf808",
X"52807234",
X"fa1380fe",
X"80085353",
X"72723480",
X"fde80852",
X"80723480",
X"fdf00852",
X"72723480",
X"fdd40852",
X"80723480",
X"fdd40852",
X"b8723484",
X"3d0d04ff",
X"3d0d028f",
X"053380fd",
X"d8085252",
X"717134fe",
X"9e3f83e0",
X"8008802e",
X"f638833d",
X"0d04803d",
X"0d853980",
X"c6933ffe",
X"b73f83e0",
X"8008802e",
X"f23880fd",
X"d8087033",
X"7081ff06",
X"83e0800c",
X"5151823d",
X"0d04803d",
X"0d80fdd0",
X"0851a371",
X"3480fddc",
X"0851ff71",
X"3480fdd4",
X"0851a871",
X"3480fdd4",
X"0851b871",
X"34823d0d",
X"04803d0d",
X"80fdd008",
X"70337081",
X"c0067030",
X"70802583",
X"e0800c51",
X"51515182",
X"3d0d04ff",
X"3d0d80fd",
X"d4087033",
X"7081ff06",
X"70832a81",
X"32708106",
X"51515152",
X"5270802e",
X"e538b072",
X"3480fdd4",
X"0851b871",
X"34833d0d",
X"04803d0d",
X"80fe8c08",
X"70088106",
X"83e0800c",
X"51823d0d",
X"04fd3d0d",
X"75775454",
X"80732594",
X"38737081",
X"05553352",
X"80f8c851",
X"85a13fff",
X"1353e939",
X"853d0d04",
X"f63d0d7c",
X"7e60625a",
X"5d5b5680",
X"59815585",
X"39747a29",
X"55745275",
X"5180dbde",
X"3f83e080",
X"087a27ed",
X"3874802e",
X"80e03874",
X"52755180",
X"dbc83f83",
X"e0800875",
X"53765254",
X"80dbee3f",
X"83e08008",
X"7a537552",
X"5680dbae",
X"3f83e080",
X"08793070",
X"7b079f2a",
X"70778024",
X"07515154",
X"55728738",
X"83e08008",
X"c2387681",
X"18b01655",
X"58588974",
X"258b38b7",
X"14537a85",
X"3880d714",
X"53727834",
X"811959ff",
X"9c398077",
X"348c3d0d",
X"04f73d0d",
X"7b7d7f62",
X"029005bb",
X"05335759",
X"565a5ab0",
X"58728338",
X"a0587570",
X"70810552",
X"33715954",
X"55903980",
X"74258e38",
X"ff147770",
X"81055933",
X"545472ef",
X"3873ff15",
X"55538073",
X"25893877",
X"52795178",
X"2def3975",
X"33755753",
X"72802e90",
X"38725279",
X"51782d75",
X"70810557",
X"3353ed39",
X"8b3d0d04",
X"ee3d0d64",
X"66696970",
X"70810552",
X"335b4a5c",
X"5e5e7680",
X"2e82f938",
X"76a52e09",
X"810682e0",
X"38807041",
X"67707081",
X"05523371",
X"4a59575f",
X"76b02e09",
X"81068c38",
X"75708105",
X"57337648",
X"57815fd0",
X"17567589",
X"2680da38",
X"76675c59",
X"805c9339",
X"778a2480",
X"c3387b8a",
X"29187b70",
X"81055d33",
X"5a5cd019",
X"7081ff06",
X"58588977",
X"27a438ff",
X"9f197081",
X"ff06ffa9",
X"1b5a5156",
X"85762792",
X"38ffbf19",
X"7081ff06",
X"51567585",
X"268a38c9",
X"19587780",
X"25ffb938",
X"7a477b40",
X"7881ff06",
X"577680e4",
X"2e80e538",
X"7680e424",
X"a7387680",
X"d82e8186",
X"387680d8",
X"24903876",
X"802e81cc",
X"3876a52e",
X"81b63881",
X"b9397680",
X"e32e818c",
X"3881af39",
X"7680f52e",
X"9b387680",
X"f5248b38",
X"7680f32e",
X"81813881",
X"99397680",
X"f82e80ca",
X"38818f39",
X"913d7055",
X"5780538a",
X"5279841b",
X"7108535b",
X"56fbfd3f",
X"7655ab39",
X"79841b71",
X"08943d70",
X"5b5b525b",
X"56758025",
X"8c387530",
X"56ad7834",
X"0280c105",
X"57765480",
X"538a5275",
X"51fbd13f",
X"77557e54",
X"b839913d",
X"70557780",
X"d8327030",
X"70802556",
X"51585690",
X"5279841b",
X"7108535b",
X"57fbad3f",
X"7555db39",
X"79841b83",
X"1233545b",
X"56983979",
X"841b7108",
X"575b5680",
X"547f537c",
X"527d51fc",
X"9c3f8739",
X"76527d51",
X"7c2d6670",
X"33588105",
X"47fd8339",
X"943d0d04",
X"7283e090",
X"0c7183e0",
X"940c04fb",
X"3d0d883d",
X"70708405",
X"52085754",
X"755383e0",
X"90085283",
X"e0940851",
X"fcc63f87",
X"3d0d04ff",
X"3d0d7370",
X"08535102",
X"93053372",
X"34700881",
X"05710c83",
X"3d0d04fc",
X"3d0d873d",
X"88115578",
X"54999353",
X"51fc993f",
X"8052873d",
X"51d13f86",
X"3d0d04fd",
X"3d0d7570",
X"5254a3c3",
X"3f83e080",
X"08145372",
X"742e9238",
X"ff137033",
X"535371af",
X"2e098106",
X"ee388113",
X"537283e0",
X"800c853d",
X"0d04fd3d",
X"0d757770",
X"535454c7",
X"3f83e080",
X"08732ea1",
X"3883e080",
X"08733152",
X"ff125271",
X"ff2e8f38",
X"72708105",
X"54337470",
X"81055634",
X"eb39ff14",
X"54807434",
X"853d0d04",
X"803d0d72",
X"51ff903f",
X"823d0d04",
X"7183e080",
X"0c04803d",
X"0d725180",
X"7134810b",
X"bc120c80",
X"0b80c012",
X"0c823d0d",
X"04800b83",
X"e2d40824",
X"8a38a4ad",
X"3fff0b83",
X"e2d40c80",
X"0b83e080",
X"0c04ff3d",
X"0d735283",
X"e0b00872",
X"2e8d38d9",
X"3f715196",
X"983f7183",
X"e0b00c83",
X"3d0d04f4",
X"3d0d7e60",
X"625c5a55",
X"8154bc15",
X"08819138",
X"7451cf3f",
X"7958807a",
X"2580f738",
X"83e38408",
X"70892a57",
X"83ff0678",
X"84807231",
X"56565773",
X"78258338",
X"73557583",
X"e2d4082e",
X"8438ff89",
X"3f83e2d4",
X"088025a6",
X"3875892b",
X"5198db3f",
X"83e38408",
X"8f3dfc11",
X"555c5481",
X"52f81b51",
X"96c53f76",
X"1483e384",
X"0c7583e2",
X"d40c7453",
X"76527851",
X"a2de3f83",
X"e0800883",
X"e3840816",
X"83e3840c",
X"78763176",
X"1b5b5956",
X"778024ff",
X"8b38617a",
X"710c5475",
X"5475802e",
X"83388154",
X"7383e080",
X"0c8e3d0d",
X"04fc3d0d",
X"fe9b3f76",
X"51feaf3f",
X"863dfc05",
X"53785277",
X"5195e83f",
X"7975710c",
X"5483e080",
X"085483e0",
X"8008802e",
X"83388154",
X"7383e080",
X"0c863d0d",
X"04fe3d0d",
X"7583e2d4",
X"08535380",
X"72248938",
X"71732e84",
X"38fdd63f",
X"7451fdea",
X"3f725197",
X"ad3f83e0",
X"80085283",
X"e0800880",
X"2e833881",
X"527183e0",
X"800c843d",
X"0d04803d",
X"0d7280c0",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d72bc",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"c40b83e0",
X"800c04fd",
X"3d0d7577",
X"71547053",
X"55539f9b",
X"3f82c813",
X"08bc150c",
X"82c01308",
X"80c0150c",
X"fceb3f73",
X"5193aa3f",
X"7383e0b0",
X"0c83e080",
X"085383e0",
X"8008802e",
X"83388153",
X"7283e080",
X"0c853d0d",
X"04fd3d0d",
X"75775553",
X"fcbf3f72",
X"802ea538",
X"bc130852",
X"73519ea5",
X"3f83e080",
X"088f3877",
X"527251ff",
X"9a3f83e0",
X"8008538a",
X"3982cc13",
X"0853d839",
X"81537283",
X"e0800c85",
X"3d0d04fe",
X"3d0dff0b",
X"83e2d40c",
X"7483e0b4",
X"0c7583e2",
X"d00c9f92",
X"3f83e080",
X"0881ff06",
X"52815371",
X"993883e2",
X"ec518e94",
X"3f83e080",
X"085283e0",
X"8008802e",
X"83387252",
X"71537283",
X"e0800c84",
X"3d0d04fa",
X"3d0d787a",
X"82c41208",
X"82c41208",
X"70722459",
X"56565757",
X"73732e09",
X"81069138",
X"80c01652",
X"80c01751",
X"9c963f83",
X"e0800855",
X"7483e080",
X"0c883d0d",
X"04f63d0d",
X"7c5b807b",
X"715c5457",
X"7a772e8c",
X"38811a82",
X"cc140854",
X"5a72f638",
X"805980d9",
X"397a5481",
X"5780707b",
X"7b315a57",
X"55ff1853",
X"74732580",
X"c13882cc",
X"14085273",
X"51ff8c3f",
X"800b83e0",
X"800825a1",
X"3882cc14",
X"0882cc11",
X"0882cc16",
X"0c7482cc",
X"120c5375",
X"802e8638",
X"7282cc17",
X"0c725480",
X"577382cc",
X"15088117",
X"575556ff",
X"b8398119",
X"59800bff",
X"1b545478",
X"73258338",
X"81547681",
X"32707506",
X"515372ff",
X"90388c3d",
X"0d04f73d",
X"0d7b7d5a",
X"5a82d052",
X"83e2d008",
X"5180cee6",
X"3f83e080",
X"0857f9e1",
X"3f795283",
X"e2d85195",
X"b43f83e0",
X"80085480",
X"5383e080",
X"08732e09",
X"81068283",
X"3883e0b4",
X"080b0b80",
X"f89c5370",
X"52569bd3",
X"3f0b0b80",
X"f89c5280",
X"c016519b",
X"c63f75bc",
X"170c7382",
X"c0170c81",
X"0b82c417",
X"0c810b82",
X"c8170c73",
X"82cc170c",
X"ff1782d0",
X"17555781",
X"913983e0",
X"c0337082",
X"2a708106",
X"51545572",
X"81803874",
X"812a8106",
X"587780f6",
X"3874842a",
X"810682c4",
X"150c83e0",
X"c0338106",
X"82c8150c",
X"79527351",
X"9aed3f73",
X"519b843f",
X"83e08008",
X"1453af73",
X"70810555",
X"3472bc15",
X"0c83e0c1",
X"5272519a",
X"ce3f83e0",
X"b80882c0",
X"150c83e0",
X"ce5280c0",
X"14519abb",
X"3f78802e",
X"8d387351",
X"782d83e0",
X"8008802e",
X"99387782",
X"cc150c75",
X"802e8638",
X"7382cc17",
X"0c7382d0",
X"15ff1959",
X"55567680",
X"2e9b3883",
X"e0b85283",
X"e2d85194",
X"aa3f83e0",
X"80088a38",
X"83e0c133",
X"5372fed2",
X"3878802e",
X"893883e0",
X"b40851fc",
X"b83f83e0",
X"b4085372",
X"83e0800c",
X"8b3d0d04",
X"ff3d0d80",
X"527351fd",
X"b53f833d",
X"0d04f03d",
X"0d627052",
X"54f6903f",
X"83e08008",
X"7453873d",
X"70535555",
X"f6b03ff7",
X"903f7351",
X"d33f6353",
X"745283e0",
X"800851fa",
X"b83f923d",
X"0d047183",
X"e0800c04",
X"80c01283",
X"e0800c04",
X"803d0d72",
X"82c01108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"7282cc11",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282c4",
X"110883e0",
X"800c5182",
X"3d0d04f9",
X"3d0d7983",
X"e0980857",
X"57817727",
X"81963876",
X"88170827",
X"818e3875",
X"33557482",
X"2e893874",
X"832eb338",
X"80fe3974",
X"54761083",
X"fe065376",
X"882a8c17",
X"08055289",
X"3dfc0551",
X"99c03f83",
X"e0800880",
X"df38029d",
X"0533893d",
X"3371882b",
X"07565680",
X"d1398454",
X"76822b83",
X"fc065376",
X"872a8c17",
X"08055289",
X"3dfc0551",
X"99903f83",
X"e08008b0",
X"38029f05",
X"33028405",
X"9e053371",
X"982b7190",
X"2b07028c",
X"059d0533",
X"70882b72",
X"078d3d33",
X"7180ffff",
X"fe800607",
X"51525357",
X"58568339",
X"81557483",
X"e0800c89",
X"3d0d04fb",
X"3d0d83e0",
X"9808fe19",
X"881208fe",
X"05555654",
X"80567473",
X"278d3882",
X"14337571",
X"29941608",
X"05575375",
X"83e0800c",
X"873d0d04",
X"fc3d0d76",
X"52800b83",
X"e0980870",
X"33515253",
X"70832e09",
X"81069138",
X"95123394",
X"13337198",
X"2b71902b",
X"07555551",
X"9b12339a",
X"13337188",
X"2b077407",
X"83e0800c",
X"55863d0d",
X"04fc3d0d",
X"7683e098",
X"08555580",
X"75238815",
X"08537281",
X"2e883888",
X"14087326",
X"85388152",
X"b2397290",
X"38733352",
X"71832e09",
X"81068538",
X"90140853",
X"728c160c",
X"72802e8d",
X"387251fe",
X"d63f83e0",
X"80085285",
X"39901408",
X"52719016",
X"0c805271",
X"83e0800c",
X"863d0d04",
X"fa3d0d78",
X"83e09808",
X"71228105",
X"7083ffff",
X"06575457",
X"5573802e",
X"88389015",
X"08537286",
X"38835280",
X"e739738f",
X"06527180",
X"da388113",
X"90160c8c",
X"15085372",
X"9038830b",
X"84172257",
X"52737627",
X"80c638bf",
X"39821633",
X"ff057484",
X"2a065271",
X"b2387251",
X"fcb13f81",
X"527183e0",
X"800827a8",
X"38835283",
X"e0800888",
X"1708279c",
X"3883e080",
X"088c160c",
X"83e08008",
X"51fdbc3f",
X"83e08008",
X"90160c73",
X"75238052",
X"7183e080",
X"0c883d0d",
X"04f23d0d",
X"60626458",
X"5e5b7533",
X"5574a02e",
X"09810688",
X"38811670",
X"4456ef39",
X"62703356",
X"5674af2e",
X"09810684",
X"38811643",
X"800b881c",
X"0c627033",
X"5155749f",
X"2691387a",
X"51fdd23f",
X"83e08008",
X"56807d34",
X"83813993",
X"3d841c08",
X"7058595f",
X"8a55a076",
X"70810558",
X"34ff1555",
X"74ff2e09",
X"8106ef38",
X"80705a5c",
X"887f085f",
X"5a7b811d",
X"7081ff06",
X"60137033",
X"70af3270",
X"30a07327",
X"71802507",
X"5151525b",
X"535e5755",
X"7480e738",
X"76ae2e09",
X"81068338",
X"8155787a",
X"27750755",
X"74802e9f",
X"38798832",
X"703078ae",
X"32703070",
X"73079f2a",
X"53515751",
X"5675bb38",
X"88598b5a",
X"ffab3976",
X"982b5574",
X"80258738",
X"80f5f017",
X"3357ff9f",
X"17557499",
X"268938e0",
X"177081ff",
X"06585578",
X"811a7081",
X"ff06721b",
X"535b5755",
X"767534fe",
X"f8397b1e",
X"7f0c8055",
X"76a02683",
X"38815574",
X"8b19347a",
X"51fc823f",
X"83e08008",
X"80f538a0",
X"547a2270",
X"852b83e0",
X"06545590",
X"1b08527c",
X"5193cb3f",
X"83e08008",
X"5783e080",
X"08818138",
X"7c335574",
X"802e80f4",
X"388b1d33",
X"70832a70",
X"81065156",
X"5674b438",
X"8b7d841d",
X"0883e080",
X"08595b5b",
X"58ff1858",
X"77ff2e9a",
X"38797081",
X"055b3379",
X"7081055b",
X"33717131",
X"52565675",
X"802ee238",
X"86397580",
X"2e96387a",
X"51fbe53f",
X"ff863983",
X"e0800856",
X"83e08008",
X"b6388339",
X"7656841b",
X"088b1133",
X"515574a7",
X"388b1d33",
X"70842a70",
X"81065156",
X"56748938",
X"83569439",
X"81569039",
X"7c51fa94",
X"3f83e080",
X"08881c0c",
X"fd813975",
X"83e0800c",
X"903d0d04",
X"f83d0d7a",
X"7c595782",
X"5483fe53",
X"77527651",
X"92903f83",
X"5683e080",
X"0880ec38",
X"81173377",
X"3371882b",
X"07565682",
X"567482d4",
X"d52e0981",
X"0680d438",
X"7554b653",
X"77527651",
X"91e43f83",
X"e0800898",
X"38811733",
X"77337188",
X"2b0783e0",
X"80085256",
X"56748182",
X"c62eac38",
X"825480d2",
X"53775276",
X"5191bb3f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62e83",
X"38815675",
X"83e0800c",
X"8a3d0d04",
X"eb3d0d67",
X"5a800b83",
X"e0980c90",
X"dd3f83e0",
X"80088106",
X"55825674",
X"83ee3874",
X"75538f3d",
X"70535759",
X"feca3f83",
X"e0800881",
X"ff065776",
X"812e0981",
X"0680d438",
X"905483be",
X"53745275",
X"5190cf3f",
X"83e08008",
X"80c9388f",
X"3d335574",
X"802e80c9",
X"3802bf05",
X"33028405",
X"be053371",
X"982b7190",
X"2b07028c",
X"05bd0533",
X"70882b72",
X"07953d33",
X"71077058",
X"7b575e52",
X"5e575957",
X"fdee3f83",
X"e0800881",
X"ff065776",
X"832e0981",
X"06863881",
X"5682f139",
X"76802e86",
X"38865682",
X"e739a454",
X"8d537852",
X"75518fe6",
X"3f815683",
X"e0800882",
X"d33802be",
X"05330284",
X"05bd0533",
X"71882b07",
X"595d77ab",
X"380280ce",
X"05330284",
X"0580cd05",
X"3371982b",
X"71902b07",
X"973d3370",
X"882b7207",
X"02940580",
X"cb053371",
X"0754525e",
X"57595602",
X"b7053378",
X"71290288",
X"05b60533",
X"028c05b5",
X"05337188",
X"2b07701d",
X"707f8c05",
X"0c5f5957",
X"595d8e3d",
X"33821b34",
X"02b90533",
X"903d3371",
X"882b075a",
X"5c78841b",
X"2302bb05",
X"33028405",
X"ba053371",
X"882b0756",
X"5c74ab38",
X"0280ca05",
X"33028405",
X"80c90533",
X"71982b71",
X"902b0796",
X"3d337088",
X"2b720702",
X"940580c7",
X"05337107",
X"51525357",
X"5e5c7476",
X"31783179",
X"842a903d",
X"33547171",
X"31535656",
X"bfcc3f83",
X"e0800882",
X"0570881c",
X"0c83e080",
X"08e08a05",
X"56567483",
X"dffe2683",
X"38825783",
X"fff67627",
X"85388357",
X"89398656",
X"76802e80",
X"db38767a",
X"3476832e",
X"098106b0",
X"380280d6",
X"05330284",
X"0580d505",
X"3371982b",
X"71902b07",
X"993d3370",
X"882b7207",
X"02940580",
X"d3053371",
X"077f9005",
X"0c525e57",
X"58568639",
X"771b901b",
X"0c841a22",
X"8c1b0819",
X"71842a05",
X"941c0c5d",
X"800b811b",
X"347983e0",
X"980c8056",
X"7583e080",
X"0c973d0d",
X"04e93d0d",
X"83e09808",
X"56855475",
X"802e8182",
X"38800b81",
X"1734993d",
X"e011466a",
X"548a3d70",
X"5458ec05",
X"51f6e63f",
X"83e08008",
X"5483e080",
X"0880df38",
X"893d3354",
X"73802e91",
X"3802ab05",
X"3370842a",
X"81065155",
X"74802e86",
X"38835480",
X"c1397651",
X"f48a3f83",
X"e08008a0",
X"170c02bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"3371079c",
X"1c0c5278",
X"981b0c53",
X"56595781",
X"0b811734",
X"74547383",
X"e0800c99",
X"3d0d04f5",
X"3d0d7d7f",
X"617283e0",
X"98085a5d",
X"5d595c80",
X"7b0c8557",
X"75802e81",
X"e0388116",
X"33810655",
X"84577480",
X"2e81d238",
X"91397481",
X"17348639",
X"800b8117",
X"34815781",
X"c0399c16",
X"08981708",
X"31557478",
X"27833874",
X"5877802e",
X"81a93898",
X"16087083",
X"ff065657",
X"7480cf38",
X"821633ff",
X"0577892a",
X"067081ff",
X"065a5578",
X"a0387687",
X"38a01608",
X"558d39a4",
X"160851f0",
X"ea3f83e0",
X"80085581",
X"7527ffa8",
X"3874a417",
X"0ca41608",
X"51f2843f",
X"83e08008",
X"5583e080",
X"08802eff",
X"893883e0",
X"800819a8",
X"170c9816",
X"0883ff06",
X"84807131",
X"51557775",
X"27833877",
X"557483ff",
X"ff065498",
X"160883ff",
X"0653a816",
X"08527957",
X"7b83387b",
X"5776518a",
X"8d3f83e0",
X"8008fed0",
X"38981608",
X"1598170c",
X"741a7876",
X"317c0817",
X"7d0c595a",
X"fed33980",
X"577683e0",
X"800c8d3d",
X"0d04fa3d",
X"0d7883e0",
X"98085556",
X"85557380",
X"2e81e138",
X"81143381",
X"06538455",
X"72802e81",
X"d3389c14",
X"08537276",
X"27833872",
X"56981408",
X"57800b98",
X"150c7580",
X"2e81b738",
X"82143370",
X"892b5653",
X"76802eb5",
X"387452ff",
X"1651bace",
X"3f83e080",
X"08ff1876",
X"54705358",
X"53babf3f",
X"83e08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed93f83",
X"e0800853",
X"810b83e0",
X"8008278b",
X"38881408",
X"83e08008",
X"26883880",
X"0b811534",
X"b03983e0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc83f",
X"83e08008",
X"8c3883e0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683e0",
X"800805a8",
X"150c8055",
X"7483e080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83e09808",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1d23f",
X"83e08008",
X"5583e080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef8",
X"3f83e080",
X"0888170c",
X"7551efa9",
X"3f83e080",
X"08557483",
X"e0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683e0",
X"9808802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f83f83e0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"86983f83",
X"e0800841",
X"83e08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"ede23f83",
X"e0800841",
X"83e08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"83a53f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f33f83e0",
X"80088332",
X"70307072",
X"079f2c83",
X"e0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"81b13f75",
X"83e0800c",
X"9e3d0d04",
X"fd3d0d75",
X"77535473",
X"33517089",
X"38713351",
X"70802ea1",
X"38733372",
X"33525372",
X"71278538",
X"ff519439",
X"70732785",
X"3881518b",
X"39811481",
X"135354d3",
X"39805170",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"77545472",
X"337081ff",
X"06525270",
X"802ea338",
X"7181ff06",
X"8114ffbf",
X"12535452",
X"70992689",
X"38a01270",
X"81ff0653",
X"51717470",
X"81055634",
X"d2398074",
X"34853d0d",
X"04ffbd3d",
X"0d80c63d",
X"0852a53d",
X"705254ff",
X"b33f80c7",
X"3d085285",
X"3d705253",
X"ffa63f72",
X"527351fe",
X"df3f80c5",
X"3d0d04fe",
X"3d0d7476",
X"53537170",
X"81055333",
X"51707370",
X"81055534",
X"70f03884",
X"3d0d04fe",
X"3d0d7452",
X"80723352",
X"5370732e",
X"8d388112",
X"81147133",
X"53545270",
X"f5387283",
X"e0800c84",
X"3d0d04fc",
X"3d0d7655",
X"7483e398",
X"082eaf38",
X"80537451",
X"87cb3f83",
X"e0800881",
X"ff06ff14",
X"7081ff06",
X"7230709f",
X"2a515255",
X"53547280",
X"2e843871",
X"dd3873fe",
X"387483e3",
X"980c863d",
X"0d04ff3d",
X"0dff0b83",
X"e3980c84",
X"af3f8151",
X"878f3f83",
X"e0800881",
X"ff065271",
X"ee3881d6",
X"3f7183e0",
X"800c833d",
X"0d04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"823f7280",
X"2ea03883",
X"e3ac1433",
X"75708105",
X"57348114",
X"7083ffff",
X"06ff1570",
X"83ffff06",
X"56525552",
X"dd39800b",
X"83e0800c",
X"863d0d04",
X"fc3d0d76",
X"787a1156",
X"53558053",
X"71742e93",
X"38721551",
X"703383e3",
X"ac133481",
X"12811454",
X"52ea3980",
X"0b83e080",
X"0c863d0d",
X"04fd3d0d",
X"905483e3",
X"98085186",
X"fe3f83e0",
X"800881ff",
X"06ff1571",
X"30713070",
X"73079f2a",
X"729f2a06",
X"52555255",
X"5372db38",
X"853d0d04",
X"ff3d0d83",
X"e3a40810",
X"83e39c08",
X"0780fe90",
X"0852710c",
X"833d0d04",
X"800b83e3",
X"a40ce13f",
X"04810b83",
X"e3a40cd8",
X"3f04ed3f",
X"047183e3",
X"a00c0480",
X"3d0d8051",
X"f43f810b",
X"83e3a40c",
X"810b83e3",
X"9c0cffb8",
X"3f823d0d",
X"04803d0d",
X"72307074",
X"07802583",
X"e39c0c51",
X"ffa23f82",
X"3d0d04fe",
X"3d0d0293",
X"053380fe",
X"94085473",
X"0c80fe90",
X"08527108",
X"70810651",
X"5170f738",
X"72087081",
X"ff0683e0",
X"800c5184",
X"3d0d0480",
X"3d0d81ff",
X"51cd3f83",
X"e0800881",
X"ff0683e0",
X"800c823d",
X"0d04ff3d",
X"0d74902b",
X"740780fe",
X"84085271",
X"0c833d0d",
X"0404fb3d",
X"0d780284",
X"059f0533",
X"70982b55",
X"57557280",
X"259b3875",
X"80ff0656",
X"805280f7",
X"51e03f83",
X"e0800881",
X"ff065473",
X"812680ff",
X"388051fe",
X"e03fff9f",
X"3f8151fe",
X"d83fff97",
X"3f7551fe",
X"e63f7498",
X"2a51fedf",
X"3f74902a",
X"7081ff06",
X"5253fed3",
X"3f74882a",
X"7081ff06",
X"5253fec7",
X"3f7481ff",
X"0651febf",
X"3f815575",
X"80c02e09",
X"81068638",
X"8195558d",
X"397580c8",
X"2e098106",
X"84388187",
X"557451fe",
X"9e3f8a55",
X"fec53f83",
X"e0800881",
X"ff067098",
X"2b545472",
X"80258c38",
X"ff157081",
X"ff065653",
X"74e23873",
X"83e0800c",
X"873d0d04",
X"fa3d0dfd",
X"be3f8051",
X"fdd33f8a",
X"54fe903f",
X"ff147081",
X"ff065553",
X"73f33873",
X"74535580",
X"c051fea6",
X"3f83e080",
X"0881ff06",
X"5473812e",
X"09810682",
X"9f3883aa",
X"5280c851",
X"fe8c3f83",
X"e0800881",
X"ff065372",
X"812e0981",
X"0681a838",
X"7454873d",
X"74115456",
X"fdc53f83",
X"e0800873",
X"34811470",
X"81ff0655",
X"53837427",
X"e538029a",
X"05335372",
X"812e0981",
X"0681d938",
X"029b0533",
X"5380ce90",
X"547281aa",
X"2e8d3881",
X"c73980e4",
X"518ace3f",
X"ff145473",
X"802e81b8",
X"38820a52",
X"81e951fd",
X"a53f83e0",
X"800881ff",
X"065372de",
X"38725280",
X"fa51fd92",
X"3f83e080",
X"0881ff06",
X"53728190",
X"38725473",
X"1653fcd3",
X"3f83e080",
X"08733481",
X"147081ff",
X"06555383",
X"7427e838",
X"873d3370",
X"862a7081",
X"06515454",
X"8c557280",
X"e3388455",
X"80de3974",
X"5281e951",
X"fccc3f83",
X"e0800881",
X"ff065382",
X"5581e956",
X"81732786",
X"38735580",
X"c15680ce",
X"90548a39",
X"80e45189",
X"c03fff14",
X"5473802e",
X"a9388052",
X"7551fc9a",
X"3f83e080",
X"0881ff06",
X"5372e138",
X"84805280",
X"d051fc86",
X"3f83e080",
X"0881ff06",
X"5372802e",
X"83388055",
X"7483e3a8",
X"348051fb",
X"803ffbbf",
X"3f883d0d",
X"04fb3d0d",
X"7754800b",
X"83e3a833",
X"70832a70",
X"81065155",
X"57557275",
X"2e098106",
X"85387389",
X"2b547352",
X"80d151fb",
X"bd3f83e0",
X"800881ff",
X"065372bd",
X"3882b8c0",
X"54fb803f",
X"83e08008",
X"81ff0653",
X"7281ff2e",
X"09810689",
X"38ff1454",
X"73e7389f",
X"397281fe",
X"2e098106",
X"963883e7",
X"ac5283e3",
X"ac51faea",
X"3ffad03f",
X"facd3f83",
X"39815580",
X"51fa823f",
X"fac13f74",
X"81ff0683",
X"e0800c87",
X"3d0d04fb",
X"3d0d7783",
X"e3ac5654",
X"8151f9e5",
X"3f83e3a8",
X"3370832a",
X"70810651",
X"54567285",
X"3873892b",
X"54735280",
X"d851fab6",
X"3f83e080",
X"0881ff06",
X"537280e4",
X"3881ff51",
X"f9cd3f81",
X"fe51f9c7",
X"3f848053",
X"74708105",
X"563351f9",
X"ba3fff13",
X"7083ffff",
X"06515372",
X"eb387251",
X"f9a93f72",
X"51f9a43f",
X"f9cd3f83",
X"e080089f",
X"0653a788",
X"5472852e",
X"8c389939",
X"80e45186",
X"f83fff14",
X"54f9b03f",
X"83e08008",
X"81ff2e84",
X"3873e938",
X"8051f8dd",
X"3ff99c3f",
X"800b83e0",
X"800c873d",
X"0d047183",
X"e7b00c88",
X"80800b83",
X"e7ac0c84",
X"80800b83",
X"e7b40c04",
X"fd3d0d77",
X"70175577",
X"05ff1a53",
X"5371ff2e",
X"94387370",
X"81055533",
X"51707370",
X"81055534",
X"ff1252e9",
X"39853d0d",
X"04fc3d0d",
X"80fda008",
X"55743383",
X"e7b834a0",
X"5483a080",
X"5383e7b0",
X"085283e7",
X"ac0851ff",
X"b73fa054",
X"83a48053",
X"83e7b008",
X"5283e7ac",
X"0851ffa4",
X"3f905483",
X"a8805383",
X"e7b00852",
X"83e7ac08",
X"51ff913f",
X"a0538052",
X"83e7b408",
X"83a08005",
X"5185d23f",
X"a0538052",
X"83e7b408",
X"83a48005",
X"5185c23f",
X"90538052",
X"83e7b408",
X"83a88005",
X"5185b23f",
X"80fda008",
X"55ff7534",
X"83a08054",
X"805383e7",
X"b0085283",
X"e7b40851",
X"fec63f80",
X"d0805483",
X"b0805383",
X"e7b00852",
X"83e7b408",
X"51feb13f",
X"86d33fa2",
X"54805383",
X"e7b4088c",
X"80055280",
X"fb9451fe",
X"9b3f80fd",
X"c4085586",
X"753480fd",
X"c8085580",
X"753480fd",
X"c0085580",
X"753480fd",
X"b00855af",
X"753480fd",
X"bc0855bf",
X"753480fd",
X"b8085580",
X"753480fd",
X"b408559f",
X"753480fd",
X"ac085580",
X"753480fd",
X"980855e0",
X"753480fd",
X"900855a2",
X"753480fd",
X"8c085583",
X"753480fd",
X"94085582",
X"7534863d",
X"0d04fc3d",
X"0d83a080",
X"54805383",
X"e7b40852",
X"83e7b008",
X"51fda13f",
X"80d08054",
X"83b08053",
X"83e7b408",
X"5283e7b0",
X"0851fd8c",
X"3fa05483",
X"a0805383",
X"e7b40852",
X"83e7b008",
X"51fcf93f",
X"a05483a4",
X"805383e7",
X"b4085283",
X"e7b00851",
X"fce63f90",
X"5483a880",
X"5383e7b4",
X"085283e7",
X"b00851fc",
X"d33f80fd",
X"a0085583",
X"e7b83375",
X"34863d0d",
X"04803d0d",
X"80fea808",
X"70088106",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"80fea808",
X"700870fe",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d80fe",
X"a8087008",
X"70812c81",
X"0683e080",
X"0c515182",
X"3d0d04ff",
X"3d0d80fe",
X"a8087008",
X"70fd0676",
X"1007720c",
X"5252833d",
X"0d04803d",
X"0d80fea8",
X"08700870",
X"822cbf06",
X"83e0800c",
X"5151823d",
X"0d04ff3d",
X"0d80fea8",
X"08700870",
X"fe830676",
X"822b0772",
X"0c525283",
X"3d0d0480",
X"3d0d80fe",
X"a8087008",
X"70882c87",
X"0683e080",
X"0c515182",
X"3d0d04ff",
X"3d0d80fe",
X"a8087008",
X"70f1ff06",
X"76882b07",
X"720c5252",
X"833d0d04",
X"803d0d80",
X"fea80870",
X"08708b2c",
X"bf0683e0",
X"800c5151",
X"823d0d04",
X"ff3d0d80",
X"fea80870",
X"0870f88f",
X"ff06768b",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d80fea8",
X"08700870",
X"912cbf06",
X"83e0800c",
X"5151823d",
X"0d04ff3d",
X"0d80fea8",
X"08700870",
X"fc87ffff",
X"0676912b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"80feb808",
X"70087088",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04803d0d",
X"80feb808",
X"70087089",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04803d0d",
X"80feb808",
X"7008708a",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04803d0d",
X"80feb808",
X"7008708b",
X"2c810683",
X"e0800c51",
X"51823d0d",
X"04fd3d0d",
X"7581e629",
X"872a80fe",
X"98085473",
X"0c853d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727081",
X"055434ff",
X"1151f039",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708405",
X"540cff11",
X"51f03984",
X"3d0d04fe",
X"3d0d8480",
X"80538052",
X"88800a51",
X"ffb33f81",
X"80805380",
X"5282800a",
X"51c63f84",
X"3d0d0480",
X"3d0d8151",
X"fc9b3f72",
X"802e8338",
X"d23f8151",
X"fcbd3f80",
X"51fcb83f",
X"8051fc85",
X"3f823d0d",
X"04fd3d0d",
X"75528054",
X"80ff7225",
X"8838810b",
X"ff801353",
X"54ffbf12",
X"51709926",
X"8638e012",
X"529e39ff",
X"9f125199",
X"71279538",
X"d012e013",
X"70545451",
X"89712788",
X"388f7327",
X"83388052",
X"73802e85",
X"38818012",
X"527181ff",
X"0683e080",
X"0c853d0d",
X"04803d0d",
X"84d8c051",
X"80717081",
X"05533470",
X"84e0c02e",
X"098106f0",
X"38823d0d",
X"04fe3d0d",
X"02970533",
X"51ff863f",
X"83e08008",
X"81ff0683",
X"e7bc0854",
X"52807324",
X"9b3883e7",
X"d8081372",
X"83e7dc08",
X"07535371",
X"733483e7",
X"bc088105",
X"83e7bc0c",
X"843d0d04",
X"fa3d0d82",
X"800a1b55",
X"8057883d",
X"fc055479",
X"53745278",
X"51cbd23f",
X"883d0d04",
X"fe3d0d83",
X"e7d00852",
X"7451d2b6",
X"3f83e080",
X"088c3876",
X"53755283",
X"e7d00851",
X"c73f843d",
X"0d04fe3d",
X"0d83e7d0",
X"08537552",
X"7451ccf5",
X"3f83e080",
X"088d3877",
X"53765283",
X"e7d00851",
X"ffa23f84",
X"3d0d04fe",
X"3d0d83e7",
X"d40851cb",
X"e93f83e0",
X"80088180",
X"802e0981",
X"068738b1",
X"8080539a",
X"3983e7d4",
X"0851cbce",
X"3f83e080",
X"0880d080",
X"2e098106",
X"9238b1b0",
X"805383e0",
X"80085283",
X"e7d40851",
X"feda3f84",
X"3d0d0480",
X"3d0dfa9b",
X"3f83e080",
X"08842980",
X"fbb80570",
X"0883e080",
X"0c51823d",
X"0d04ee3d",
X"0d804380",
X"42804180",
X"705a5bfd",
X"d43f800b",
X"83e7bc0c",
X"800b83e7",
X"dc0c80f9",
X"9451c6bb",
X"3f81800b",
X"83e7dc0c",
X"80f99851",
X"c6ad3f80",
X"d00b83e7",
X"bc0c7830",
X"707a0780",
X"2570872b",
X"83e7dc0c",
X"5155f98a",
X"3f83e080",
X"085280f9",
X"a051c687",
X"3f80f80b",
X"83e7bc0c",
X"78813270",
X"30707207",
X"80257087",
X"2b83e7dc",
X"0c515656",
X"fef13f83",
X"e0800852",
X"80f9ac51",
X"c5dd3f81",
X"a00b83e7",
X"bc0c7882",
X"32703070",
X"72078025",
X"70872b83",
X"e7dc0c51",
X"5683e7d4",
X"085256c6",
X"f73f83e0",
X"80085280",
X"f9b451c5",
X"ae3f81f0",
X"0b83e7bc",
X"0c810b83",
X"e7c05b58",
X"83e7bc08",
X"82197a32",
X"70307072",
X"07802570",
X"872b83e7",
X"dc0c5157",
X"8e3d7055",
X"ff1b5457",
X"57579992",
X"3f797084",
X"055b0851",
X"c6ae3f74",
X"5483e080",
X"08537752",
X"80f9bc51",
X"c4e13fa8",
X"1783e7bc",
X"0c811858",
X"77852e09",
X"8106ffb0",
X"3883900b",
X"83e7bc0c",
X"78873270",
X"30707207",
X"80257087",
X"2b83e7dc",
X"0c515656",
X"f8bc3f80",
X"f9cc5583",
X"e0800880",
X"2e8e3883",
X"e7d00851",
X"c5da3f83",
X"e0800855",
X"745280f9",
X"d451c48f",
X"3f83e00b",
X"83e7bc0c",
X"78883270",
X"30707207",
X"80257087",
X"2b83e7dc",
X"0c515780",
X"f9e05255",
X"c3ed3f86",
X"8da051f9",
X"843f8052",
X"913d7052",
X"5599ea3f",
X"83527451",
X"99e33f61",
X"19597880",
X"25853880",
X"59903988",
X"79258538",
X"88598739",
X"78882682",
X"db387882",
X"2b5580f7",
X"f0150804",
X"f6a43f83",
X"e0800861",
X"57557581",
X"2e098106",
X"893883e0",
X"80081055",
X"903975ff",
X"2e098106",
X"883883e0",
X"8008812c",
X"55907525",
X"85389055",
X"88397480",
X"24833881",
X"557451f6",
X"813f8290",
X"39f6943f",
X"83e08008",
X"61055574",
X"80258538",
X"80558839",
X"87752583",
X"38875574",
X"51f6903f",
X"81ee3960",
X"87386280",
X"2e81e538",
X"83e0a408",
X"83e0a00c",
X"8aea0b83",
X"e0a80c83",
X"e7d40851",
X"ffb4d53f",
X"fae93f81",
X"c7396056",
X"80762599",
X"388a830b",
X"83e0a80c",
X"83e7b415",
X"70085255",
X"ffb4b53f",
X"74085291",
X"39758025",
X"913883e7",
X"b4150851",
X"c3c83f80",
X"52fd1951",
X"b8396280",
X"2e818d38",
X"83e7b415",
X"700883e7",
X"c008720c",
X"83e7c00c",
X"fd1a7053",
X"51558b82",
X"3f83e080",
X"08568051",
X"8af83f83",
X"e0800852",
X"74518790",
X"3f755280",
X"5187893f",
X"80d63960",
X"55807525",
X"b83883e0",
X"ac0883e0",
X"a00c8aea",
X"0b83e0a8",
X"0c83e7d0",
X"0851ffb3",
X"bf3f83e7",
X"d00851ff",
X"b1ce3f83",
X"e0800881",
X"ff067052",
X"55f5a33f",
X"74802e9c",
X"388155a0",
X"39748025",
X"933883e7",
X"d00851c2",
X"b93f8051",
X"f5883f84",
X"39628738",
X"7a802efa",
X"8a388055",
X"7483e080",
X"0c943d0d",
X"04fe3d0d",
X"f5873f83",
X"e0800880",
X"2e863880",
X"5180f739",
X"f58f3f83",
X"e0800880",
X"eb38f5b5",
X"3f83e080",
X"08802eaa",
X"388151f2",
X"d43fefa9",
X"3f800b83",
X"e7bc0cf9",
X"b93f83e0",
X"800853ff",
X"0b83e7bc",
X"0cf1b33f",
X"72be3872",
X"51f2b23f",
X"bc39f4e9",
X"3f83e080",
X"08802eb1",
X"388151f2",
X"a03feef5",
X"3f8a830b",
X"83e0a80c",
X"83e7c008",
X"51ffb284",
X"3fff0b83",
X"e7bc0cf0",
X"fd3f83e7",
X"c0085280",
X"5185993f",
X"8151f5d3",
X"3f843d0d",
X"04fc3d0d",
X"84808052",
X"84a48080",
X"51c58c3f",
X"83e08008",
X"80c33888",
X"ea3f80fe",
X"bc51c9cc",
X"3f83e080",
X"0883e7d4",
X"085480f9",
X"e85383e0",
X"80085255",
X"c4a73f83",
X"e0800884",
X"38f7c03f",
X"b0808054",
X"80c08053",
X"80f9f452",
X"7451f78a",
X"3f8151f4",
X"fa3f92f6",
X"3f8151f4",
X"f23ffe91",
X"3ffc3983",
X"e08c0802",
X"83e08c0c",
X"fb3d0d02",
X"80fa840b",
X"83e0a40c",
X"80fa880b",
X"83e09c0c",
X"80fa8c0b",
X"83e0ac0c",
X"83e08c08",
X"fc050c80",
X"0b83e7c0",
X"0b83e08c",
X"08f8050c",
X"83e08c08",
X"f4050cc2",
X"ee3f83e0",
X"80088605",
X"fc0683e0",
X"8c08f005",
X"0c0283e0",
X"8c08f005",
X"08310d83",
X"3d7083e0",
X"8c08f805",
X"08708405",
X"83e08c08",
X"f8050c0c",
X"51ffbfb6",
X"3f83e08c",
X"08f40508",
X"810583e0",
X"8c08f405",
X"0c83e08c",
X"08f40508",
X"862e0981",
X"06ffac38",
X"84a88080",
X"51ec8b3f",
X"ff0b83e7",
X"bc0c800b",
X"83e7dc0c",
X"84d8c00b",
X"83e7d80c",
X"8151efd9",
X"3f8151f0",
X"823f8051",
X"effd3f81",
X"51f0a73f",
X"8151f184",
X"3f8251f0",
X"ce3f8051",
X"f1ac3f80",
X"d0955280",
X"51ffbcf4",
X"3ffdbe3f",
X"83e08c08",
X"fc05080d",
X"800b83e0",
X"800c873d",
X"0d83e08c",
X"0c04803d",
X"0d81ff51",
X"800b83e7",
X"e81234ff",
X"115170f4",
X"38823d0d",
X"04ff3d0d",
X"73703353",
X"51811133",
X"71347181",
X"1234833d",
X"0d04fb3d",
X"0d777956",
X"56807071",
X"55555271",
X"7525ac38",
X"72167033",
X"70147081",
X"ff065551",
X"51517174",
X"27893881",
X"127081ff",
X"06535171",
X"81147083",
X"ffff0655",
X"52547473",
X"24d63871",
X"83e0800c",
X"873d0d04",
X"fc3d0d76",
X"55ffb69d",
X"3f83e080",
X"08802ef5",
X"3883ea84",
X"08860570",
X"81ff0652",
X"53ffb3f4",
X"3f8439fb",
X"803fffb5",
X"fc3f83e0",
X"8008812e",
X"f2388054",
X"731553ff",
X"b4d03f83",
X"e0800873",
X"34811454",
X"73852e09",
X"8106e938",
X"8439fad5",
X"3fffb5d1",
X"3f83e080",
X"08802ef2",
X"38743383",
X"e7e83481",
X"153383e7",
X"e9348215",
X"3383e7ea",
X"34831533",
X"83e7eb34",
X"845283e7",
X"e851feba",
X"3f83e080",
X"0881ff06",
X"84163356",
X"5372752e",
X"0981068d",
X"38ffb4c1",
X"3f83e080",
X"08802e9a",
X"3883ea84",
X"08a82e09",
X"81068938",
X"860b83ea",
X"840c8739",
X"a80b83ea",
X"840c80e4",
X"51efd23f",
X"863d0d04",
X"f43d0d7e",
X"60595580",
X"5d807582",
X"2b7183ea",
X"88120c83",
X"ea9c175b",
X"5b577679",
X"3477772e",
X"83b83876",
X"527751ff",
X"bdff3f8e",
X"3dfc0554",
X"905383e9",
X"f0527751",
X"ffbdba3f",
X"7c567590",
X"2e098106",
X"83943883",
X"e9f051fd",
X"943f83e9",
X"f251fd8d",
X"3f83e9f4",
X"51fd863f",
X"7683ea80",
X"0c7751ff",
X"bb863f80",
X"f8a45283",
X"e0800851",
X"ffaa8a3f",
X"83e08008",
X"812e0981",
X"0680d438",
X"7683ea98",
X"0c820b83",
X"e9f034ff",
X"960b83e9",
X"f1347751",
X"ffbdcb3f",
X"83e08008",
X"5583e080",
X"08772588",
X"3883e080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"e9f23474",
X"83e9f334",
X"7683e9f4",
X"34ff800b",
X"83e9f534",
X"81903983",
X"e9f03383",
X"e9f13371",
X"882b0756",
X"5b7483ff",
X"ff2e0981",
X"0680e838",
X"fe800b83",
X"ea980c81",
X"0b83ea80",
X"0cff0b83",
X"e9f034ff",
X"0b83e9f1",
X"347751ff",
X"bcd83f83",
X"e0800883",
X"eaa00c83",
X"e0800855",
X"83e08008",
X"80258838",
X"83e08008",
X"8f055574",
X"842c7083",
X"ffff0670",
X"882a5851",
X"557583e9",
X"f2347483",
X"e9f33476",
X"83e9f434",
X"ff800b83",
X"e9f53481",
X"0b83e9ff",
X"34a53974",
X"85962e09",
X"810680fe",
X"387583ea",
X"980c7751",
X"ffbc8c3f",
X"83e9ff33",
X"83e08008",
X"07557483",
X"e9ff3483",
X"e9ff3381",
X"06557480",
X"2e833884",
X"5783e9f4",
X"3383e9f5",
X"3371882b",
X"07565c74",
X"81802e09",
X"8106a138",
X"83e9f233",
X"83e9f333",
X"71882b07",
X"565bad80",
X"75278738",
X"76820757",
X"9c397681",
X"07579639",
X"7482802e",
X"09810687",
X"38768307",
X"57873974",
X"81ff268a",
X"387783ea",
X"881b0c76",
X"79348e3d",
X"0d04803d",
X"0d728429",
X"83ea8805",
X"700883e0",
X"800c5182",
X"3d0d04fe",
X"3d0d800b",
X"83e9ec0c",
X"800b83e9",
X"e80cff0b",
X"83e7e40c",
X"a80b83ea",
X"840cae51",
X"ffaebd3f",
X"800b83ea",
X"88545280",
X"73708405",
X"550c8112",
X"5271842e",
X"098106ef",
X"38843d0d",
X"04fe3d0d",
X"74028405",
X"96052253",
X"5371802e",
X"97387270",
X"81055433",
X"51ffaedb",
X"3fff1270",
X"83ffff06",
X"5152e639",
X"843d0d04",
X"fe3d0d02",
X"92052253",
X"82ac51ea",
X"e43f80c3",
X"51ffaeb7",
X"3f819651",
X"ead73f72",
X"5283e7e8",
X"51ffb23f",
X"725283e7",
X"e851f8ee",
X"3f83e080",
X"0881ff06",
X"51ffae93",
X"3f843d0d",
X"04ffb13d",
X"0d80d13d",
X"f80551f9",
X"973f83e9",
X"ec088105",
X"83e9ec0c",
X"80cf3d33",
X"cf117081",
X"ff065156",
X"56748326",
X"88ed3875",
X"8f06ff05",
X"567583e7",
X"e4082e9b",
X"38758326",
X"96387583",
X"e7e40c75",
X"842983ea",
X"88057008",
X"53557551",
X"fa963f80",
X"762488c9",
X"38758429",
X"83ea8805",
X"55740880",
X"2e88ba38",
X"83e7e408",
X"842983ea",
X"88057008",
X"02880582",
X"b9053352",
X"5b557480",
X"d22e84b1",
X"387480d2",
X"24903874",
X"bf2e9c38",
X"7480d02e",
X"81d73887",
X"f8397480",
X"d32e80d2",
X"387480d7",
X"2e81c638",
X"87e73902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"5656ffad",
X"953f80c1",
X"51ffacc7",
X"3ff6e73f",
X"860b83e7",
X"e8348152",
X"83e7e851",
X"ffae823f",
X"8151fde4",
X"3f748938",
X"860b83ea",
X"840c8739",
X"a80b83ea",
X"840cffac",
X"e13f80c1",
X"51ffac93",
X"3ff6b33f",
X"900b83e9",
X"ff338106",
X"56567480",
X"2e833898",
X"5683e9f4",
X"3383e9f5",
X"3371882b",
X"07565974",
X"81802e09",
X"81069c38",
X"83e9f233",
X"83e9f333",
X"71882b07",
X"5657ad80",
X"75278c38",
X"75818007",
X"56853975",
X"a0075675",
X"83e7e834",
X"ff0b83e7",
X"e934e00b",
X"83e7ea34",
X"800b83e7",
X"eb348452",
X"83e7e851",
X"ffacf63f",
X"8451869e",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055659",
X"ffabd33f",
X"7951ffb6",
X"d23f83e0",
X"8008802e",
X"8b3880ce",
X"51ffaaf7",
X"3f85f239",
X"80c151ff",
X"aaed3fff",
X"abf53fff",
X"a9f73f83",
X"ea980858",
X"8375259b",
X"3883e9f4",
X"3383e9f5",
X"3371882b",
X"07fc1771",
X"297a0583",
X"80055a51",
X"578d3974",
X"81802918",
X"ff800558",
X"81805780",
X"5676762e",
X"9338ffaa",
X"c93f83e0",
X"800883e7",
X"e8173481",
X"1656ea39",
X"ffaab73f",
X"83e08008",
X"81ff0677",
X"5383e7e8",
X"5256f4d6",
X"3f83e080",
X"0881ff06",
X"5575752e",
X"09810681",
X"8a38ffaa",
X"b93f80c1",
X"51ffa9eb",
X"3fffaaf3",
X"3f775279",
X"51ffb4e1",
X"3f805e80",
X"d13dfdf4",
X"05547653",
X"83e7e852",
X"7951ffb2",
X"ee3f0282",
X"b9053355",
X"81587480",
X"d72e0981",
X"06bd3880",
X"d13dfdf0",
X"05547653",
X"8f3d7053",
X"7a5259ff",
X"b3f33f80",
X"5676762e",
X"a2387519",
X"83e7e817",
X"33713370",
X"72327030",
X"70802570",
X"307e0681",
X"1d5d5e51",
X"5151525b",
X"55db3982",
X"ac51e59d",
X"3f77802e",
X"863880c3",
X"51843980",
X"ce51ffa8",
X"e63fffa9",
X"ee3fffa7",
X"f03f83dd",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055955",
X"80705d59",
X"ffa9873f",
X"80c151ff",
X"a8b93f83",
X"ea800879",
X"2e82de38",
X"83eaa008",
X"80fc0555",
X"80fd5274",
X"51868b3f",
X"83e08008",
X"5b778224",
X"b238ff18",
X"70872b83",
X"ffff8006",
X"80fbd805",
X"83e7e859",
X"57558180",
X"55757081",
X"05573377",
X"70810559",
X"34ff1570",
X"81ff0651",
X"5574ea38",
X"828d3977",
X"82e82e81",
X"ab387782",
X"e92e0981",
X"0681b238",
X"80fa9051",
X"ffaed43f",
X"78587787",
X"32703070",
X"72078025",
X"7a8a3270",
X"30707207",
X"80257307",
X"53545a51",
X"57557580",
X"2e973878",
X"78269238",
X"a00b83e7",
X"e81a3481",
X"197081ff",
X"065a55eb",
X"39811870",
X"81ff0659",
X"558a7827",
X"ffbc388f",
X"5883e7e3",
X"183383e7",
X"e81934ff",
X"187081ff",
X"06595577",
X"8426ea38",
X"9058800b",
X"83e7e819",
X"34811870",
X"81ff0670",
X"982b5259",
X"55748025",
X"e93880c6",
X"557a858f",
X"24843880",
X"c2557483",
X"e7e83480",
X"f10b83e7",
X"eb34810b",
X"83e7ec34",
X"7a83e7e9",
X"347a882c",
X"557483e7",
X"ea3480cb",
X"3982f078",
X"2580c438",
X"7780fd29",
X"fd97d305",
X"527951ff",
X"b18f3f80",
X"d13dfdec",
X"055480fd",
X"5383e7e8",
X"527951ff",
X"b0c73f7b",
X"81195956",
X"7580fc24",
X"83387858",
X"77882c55",
X"7483e8e5",
X"347783e8",
X"e6347583",
X"e8e73481",
X"805980cc",
X"3983ea98",
X"08578378",
X"259b3883",
X"e9f43383",
X"e9f53371",
X"882b07fc",
X"1a712979",
X"05838005",
X"5951598d",
X"39778180",
X"2917ff80",
X"05578180",
X"59765279",
X"51ffb09d",
X"3f80d13d",
X"fdec0554",
X"785383e7",
X"e8527951",
X"ffafd63f",
X"7851f6b8",
X"3fffa68b",
X"3fffa48d",
X"3f8b3983",
X"e9e80881",
X"0583e9e8",
X"0c80d13d",
X"0d04f6d9",
X"3feb9e3f",
X"f939fc3d",
X"0d767871",
X"842983ea",
X"88057008",
X"51535353",
X"709e3880",
X"ce723480",
X"cf0b8113",
X"3480ce0b",
X"82133480",
X"c50b8313",
X"34708413",
X"3480e739",
X"83ea9c13",
X"335480d2",
X"72347382",
X"2a708106",
X"515180cf",
X"53708438",
X"80d75372",
X"811334a0",
X"0b821334",
X"73830651",
X"70812e9e",
X"38708124",
X"88387080",
X"2e8f389f",
X"3970822e",
X"92387083",
X"2e923893",
X"3980d855",
X"8e3980d3",
X"55893980",
X"cd558439",
X"80c45574",
X"83133480",
X"c40b8413",
X"34800b85",
X"1334863d",
X"0d04fd3d",
X"0d755480",
X"740c800b",
X"84150c80",
X"0b88150c",
X"80fda408",
X"70337081",
X"ff067081",
X"2a813271",
X"81327181",
X"06718106",
X"31841a0c",
X"56567083",
X"2a813271",
X"822a8132",
X"71810671",
X"81063179",
X"0c525551",
X"515180fd",
X"9c087033",
X"70098106",
X"88170c51",
X"51853d0d",
X"04fe3d0d",
X"74765452",
X"7151ff9a",
X"3f72812e",
X"a2388173",
X"268d3872",
X"822eab38",
X"72832e9f",
X"38e63971",
X"08e23884",
X"1208dd38",
X"881208d8",
X"38a03988",
X"1208812e",
X"098106cc",
X"38943988",
X"1208812e",
X"8d387108",
X"89388412",
X"08802eff",
X"b738843d",
X"0d0483e0",
X"8c080283",
X"e08c0cfd",
X"3d0d8053",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"83d43f83",
X"e0800870",
X"83e0800c",
X"54853d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cfd3d",
X"0d815383",
X"e08c088c",
X"05085283",
X"e08c0888",
X"05085183",
X"a13f83e0",
X"80087083",
X"e0800c54",
X"853d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cf93d0d",
X"800b83e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"8025b938",
X"83e08c08",
X"88050830",
X"83e08c08",
X"88050c80",
X"0b83e08c",
X"08f4050c",
X"83e08c08",
X"fc05088a",
X"38810b83",
X"e08c08f4",
X"050c83e0",
X"8c08f405",
X"0883e08c",
X"08fc050c",
X"83e08c08",
X"8c050880",
X"25b93883",
X"e08c088c",
X"05083083",
X"e08c088c",
X"050c800b",
X"83e08c08",
X"f0050c83",
X"e08c08fc",
X"05088a38",
X"810b83e0",
X"8c08f005",
X"0c83e08c",
X"08f00508",
X"83e08c08",
X"fc050c80",
X"5383e08c",
X"088c0508",
X"5283e08c",
X"08880508",
X"5181df3f",
X"83e08008",
X"7083e08c",
X"08f8050c",
X"5483e08c",
X"08fc0508",
X"802e9038",
X"83e08c08",
X"f8050830",
X"83e08c08",
X"f8050c83",
X"e08c08f8",
X"05087083",
X"e0800c54",
X"893d0d83",
X"e08c0c04",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"800b83e0",
X"8c08fc05",
X"0c83e08c",
X"08880508",
X"80259938",
X"83e08c08",
X"88050830",
X"83e08c08",
X"88050c81",
X"0b83e08c",
X"08fc050c",
X"83e08c08",
X"8c050880",
X"25903883",
X"e08c088c",
X"05083083",
X"e08c088c",
X"050c8153",
X"83e08c08",
X"8c050852",
X"83e08c08",
X"88050851",
X"bd3f83e0",
X"80087083",
X"e08c08f8",
X"050c5483",
X"e08c08fc",
X"0508802e",
X"903883e0",
X"8c08f805",
X"083083e0",
X"8c08f805",
X"0c83e08c",
X"08f80508",
X"7083e080",
X"0c54873d",
X"0d83e08c",
X"0c0483e0",
X"8c080283",
X"e08c0cfd",
X"3d0d810b",
X"83e08c08",
X"fc050c80",
X"0b83e08c",
X"08f8050c",
X"83e08c08",
X"8c050883",
X"e08c0888",
X"050827b9",
X"3883e08c",
X"08fc0508",
X"802eae38",
X"800b83e0",
X"8c088c05",
X"0824a238",
X"83e08c08",
X"8c050810",
X"83e08c08",
X"8c050c83",
X"e08c08fc",
X"05081083",
X"e08c08fc",
X"050cffb8",
X"3983e08c",
X"08fc0508",
X"802e80e1",
X"3883e08c",
X"088c0508",
X"83e08c08",
X"88050826",
X"ad3883e0",
X"8c088805",
X"0883e08c",
X"088c0508",
X"3183e08c",
X"0888050c",
X"83e08c08",
X"f8050883",
X"e08c08fc",
X"05080783",
X"e08c08f8",
X"050c83e0",
X"8c08fc05",
X"08812a83",
X"e08c08fc",
X"050c83e0",
X"8c088c05",
X"08812a83",
X"e08c088c",
X"050cff95",
X"3983e08c",
X"08900508",
X"802e9338",
X"83e08c08",
X"88050870",
X"83e08c08",
X"f4050c51",
X"913983e0",
X"8c08f805",
X"087083e0",
X"8c08f405",
X"0c5183e0",
X"8c08f405",
X"0883e080",
X"0c853d0d",
X"83e08c0c",
X"0483e08c",
X"080283e0",
X"8c0cff3d",
X"0d800b83",
X"e08c08fc",
X"050c83e0",
X"8c088805",
X"088106ff",
X"11700970",
X"83e08c08",
X"8c050806",
X"83e08c08",
X"fc050811",
X"83e08c08",
X"fc050c83",
X"e08c0888",
X"0508812a",
X"83e08c08",
X"88050c83",
X"e08c088c",
X"05081083",
X"e08c088c",
X"050c5151",
X"515183e0",
X"8c088805",
X"08802e84",
X"38ffab39",
X"83e08c08",
X"fc050870",
X"83e0800c",
X"51833d0d",
X"83e08c0c",
X"04000000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002ac4",
X"00002b05",
X"00002b27",
X"00002b4e",
X"00002b4e",
X"00002b4e",
X"00002b4e",
X"00002bbf",
X"00002c11",
X"25732025",
X"73000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"524f4d00",
X"42494e00",
X"43415200",
X"6e616d65",
X"20000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00003c50",
X"00003c54",
X"00003c5c",
X"00003c68",
X"00003c74",
X"00003c80",
X"00003c8c",
X"00003c90",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"0001d20f",
X"0001d400",
X"0001d401",
X"0001d409",
X"0001d010",
X"0001d301",
X"0001d300",
X"0001d20a",
X"0001d01b",
X"0001d016",
X"0001d019",
X"0001d018",
X"0001d017",
X"0001d01a",
X"0001d403",
X"0001d402",
X"0001d40e",
X"0004007c",
X"00040078",
X"00040074",
X"00040068",
X"00040060",
X"0004005c",
X"00040058",
X"00040054",
X"00040050",
X"0004004c",
X"00040048",
X"00040044",
X"00040040",
X"00040034",
X"00040030",
X"0004002c",
X"00040028",
X"00040024",
X"00040020",
X"0004001c",
X"00040018",
X"00040014",
X"00040010",
X"0004000c",
X"00040008",
X"00040004",
X"00040000",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
