
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b81d3",
X"b4738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b81da",
X"c80c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83c08008",
X"83c08408",
X"83c08808",
X"757580f1",
X"942d5050",
X"83c08008",
X"5683c088",
X"0c83c084",
X"0c83c080",
X"0c510483",
X"c0800883",
X"c0840883",
X"c0880875",
X"7580f0d3",
X"2d505083",
X"c0800856",
X"83c0880c",
X"83c0840c",
X"83c0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80dbef04",
X"fd3d0d75",
X"705254ae",
X"a63f83c0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"c0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83c0",
X"8008732e",
X"a13883c0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183c0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83c2d008",
X"248a38b4",
X"f73fff0b",
X"83c2d00c",
X"800b83c0",
X"800c04ff",
X"3d0d7352",
X"83c0ac08",
X"722e8d38",
X"d93f7151",
X"96993f71",
X"83c0ac0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"558154bc",
X"15088191",
X"387451cf",
X"3f795880",
X"7a2580f7",
X"3883c380",
X"0870892a",
X"5783ff06",
X"78848072",
X"31565657",
X"73782583",
X"38735575",
X"83c2d008",
X"2e8438ff",
X"893f83c2",
X"d0088025",
X"a6387589",
X"2b5198dc",
X"3f83c380",
X"088f3dfc",
X"11555c54",
X"8152f81b",
X"5196c63f",
X"761483c3",
X"800c7583",
X"c2d00c74",
X"53765278",
X"51b3a83f",
X"83c08008",
X"83c38008",
X"1683c380",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8b3861",
X"7a710c54",
X"75547580",
X"2e833881",
X"547383c0",
X"800c8e3d",
X"0d04fc3d",
X"0dfe9b3f",
X"7651feaf",
X"3f863dfc",
X"05537852",
X"775195e9",
X"3f797571",
X"0c5483c0",
X"80085483",
X"c0800880",
X"2e833881",
X"547383c0",
X"800c863d",
X"0d04fe3d",
X"0d7583c2",
X"d0085353",
X"80722489",
X"3871732e",
X"8438fdd6",
X"3f7451fd",
X"ea3f7251",
X"97ae3f83",
X"c0800852",
X"83c08008",
X"802e8338",
X"81527183",
X"c0800c84",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"c0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"c0800c51",
X"823d0d04",
X"80c40b83",
X"c0800c04",
X"fd3d0d75",
X"77715470",
X"535553a9",
X"fe3f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfceb3f",
X"735193ab",
X"3f7383c0",
X"ac0c83c0",
X"80085383",
X"c0800880",
X"2e833881",
X"537283c0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcbf3f",
X"72802ea5",
X"38bc1308",
X"527351a9",
X"883f83c0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"c0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83c0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83c2d0",
X"0c7483c0",
X"b00c7583",
X"c2cc0caf",
X"dc3f83c0",
X"800881ff",
X"06528153",
X"71993883",
X"c2e8518e",
X"943f83c0",
X"80085283",
X"c0800880",
X"2e833872",
X"52715372",
X"83c0800c",
X"843d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"51a6f93f",
X"83c08008",
X"557483c0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"c0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283c2cc",
X"085180df",
X"d63f83c0",
X"800857f9",
X"e13f7952",
X"83c2d451",
X"95b73f83",
X"c0800854",
X"805383c0",
X"8008732e",
X"09810682",
X"833883c0",
X"b0080b0b",
X"81d8bc53",
X"705256a6",
X"b63f0b0b",
X"81d8bc52",
X"80c01651",
X"a6a93f75",
X"bc170c73",
X"82c0170c",
X"810b82c4",
X"170c810b",
X"82c8170c",
X"7382cc17",
X"0cff1782",
X"d0175557",
X"81913983",
X"c0bc3370",
X"822a7081",
X"06515455",
X"72818038",
X"74812a81",
X"06587780",
X"f6387484",
X"2a810682",
X"c4150c83",
X"c0bc3381",
X"0682c815",
X"0c795273",
X"51a5d03f",
X"7351a5e7",
X"3f83c080",
X"081453af",
X"73708105",
X"553472bc",
X"150c83c0",
X"bd527251",
X"a5b13f83",
X"c0b40882",
X"c0150c83",
X"c0ca5280",
X"c01451a5",
X"9e3f7880",
X"2e8d3873",
X"51782d83",
X"c0800880",
X"2e993877",
X"82cc150c",
X"75802e86",
X"387382cc",
X"170c7382",
X"d015ff19",
X"59555676",
X"802e9b38",
X"83c0b452",
X"83c2d451",
X"94ad3f83",
X"c080088a",
X"3883c0bd",
X"335372fe",
X"d2387880",
X"2e893883",
X"c0b00851",
X"fcb83f83",
X"c0b00853",
X"7283c080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb53f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f690",
X"3f83c080",
X"08745387",
X"3d705355",
X"55f6b03f",
X"f7903f73",
X"51d33f63",
X"53745283",
X"c0800851",
X"fab83f92",
X"3d0d0471",
X"83c0800c",
X"0480c012",
X"83c0800c",
X"04803d0d",
X"7282c011",
X"0883c080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883c0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"c0800c51",
X"823d0d04",
X"f93d0d79",
X"83c09008",
X"57578177",
X"27819638",
X"76881708",
X"27818e38",
X"75335574",
X"822e8938",
X"74832eb3",
X"3880fe39",
X"74547610",
X"83fe0653",
X"76882a8c",
X"17080552",
X"893dfc05",
X"51aa8a3f",
X"83c08008",
X"80df3802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d13984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"51a9da3f",
X"83c08008",
X"b038029f",
X"05330284",
X"059e0533",
X"71982b71",
X"902b0702",
X"8c059d05",
X"3370882b",
X"72078d3d",
X"337180ff",
X"fffe8006",
X"07515253",
X"57585683",
X"39815574",
X"83c0800c",
X"893d0d04",
X"fb3d0d83",
X"c09008fe",
X"19881208",
X"fe055556",
X"54805674",
X"73278d38",
X"82143375",
X"71299416",
X"08055753",
X"7583c080",
X"0c873d0d",
X"04fc3d0d",
X"7652800b",
X"83c09008",
X"70335152",
X"5370832e",
X"09810691",
X"38951233",
X"94133371",
X"982b7190",
X"2b075555",
X"519b1233",
X"9a133371",
X"882b0774",
X"0783c080",
X"0c55863d",
X"0d04fc3d",
X"0d7683c0",
X"90085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"fed63f83",
X"c0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183c080",
X"0c863d0d",
X"04fa3d0d",
X"7883c090",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fcb13f",
X"81527183",
X"c0800827",
X"a8388352",
X"83c08008",
X"88170827",
X"9c3883c0",
X"80088c16",
X"0c83c080",
X"0851fdbc",
X"3f83c080",
X"0890160c",
X"73752380",
X"527183c0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585e5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"9f269138",
X"7a51fdd2",
X"3f83c080",
X"0856807d",
X"34838139",
X"933d841c",
X"08705859",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"3880705a",
X"5c887f08",
X"5f5a7b81",
X"1d7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535e57",
X"557480e7",
X"3876ae2e",
X"09810683",
X"38815578",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675bb",
X"3888598b",
X"5affab39",
X"76982b55",
X"74802587",
X"3881d2c4",
X"173357ff",
X"9f175574",
X"99268938",
X"e0177081",
X"ff065855",
X"78811a70",
X"81ff0672",
X"1b535b57",
X"55767534",
X"fef8397b",
X"1e7f0c80",
X"5576a026",
X"83388155",
X"748b1934",
X"7a51fc82",
X"3f83c080",
X"0880f538",
X"a0547a22",
X"70852b83",
X"e0065455",
X"901b0852",
X"7c51a495",
X"3f83c080",
X"085783c0",
X"80088181",
X"387c3355",
X"74802e80",
X"f4388b1d",
X"3370832a",
X"70810651",
X"565674b4",
X"388b7d84",
X"1d0883c0",
X"8008595b",
X"5b58ff18",
X"5877ff2e",
X"9a387970",
X"81055b33",
X"79708105",
X"5b337171",
X"31525656",
X"75802ee2",
X"38863975",
X"802e9638",
X"7a51fbe5",
X"3fff8639",
X"83c08008",
X"5683c080",
X"08b63883",
X"39765684",
X"1b088b11",
X"33515574",
X"a7388b1d",
X"3370842a",
X"70810651",
X"56567489",
X"38835694",
X"39815690",
X"397c51fa",
X"943f83c0",
X"8008881c",
X"0cfd8139",
X"7583c080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"51a2da3f",
X"835683c0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"51a2ae3f",
X"83c08008",
X"98388117",
X"33773371",
X"882b0783",
X"c0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"7651a285",
X"3f83c080",
X"08983881",
X"17337733",
X"71882b07",
X"83c08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583c080",
X"0c8a3d0d",
X"04eb3d0d",
X"675a800b",
X"83c0900c",
X"a1a73f83",
X"c0800881",
X"06558256",
X"7483ef38",
X"7475538f",
X"3d705357",
X"59feca3f",
X"83c08008",
X"81ff0657",
X"76812e09",
X"810680d4",
X"38905483",
X"be537452",
X"7551a199",
X"3f83c080",
X"0880c938",
X"8f3d3355",
X"74802e80",
X"c93802bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"33710770",
X"587b575e",
X"525e5759",
X"57fdee3f",
X"83c08008",
X"81ff0657",
X"76832e09",
X"81068638",
X"815682f2",
X"3976802e",
X"86388656",
X"82e839a4",
X"548d5378",
X"527551a0",
X"b03f8156",
X"83c08008",
X"82d43802",
X"be053302",
X"8405bd05",
X"3371882b",
X"07595d77",
X"ab380280",
X"ce053302",
X"840580cd",
X"05337198",
X"2b71902b",
X"07973d33",
X"70882b72",
X"07029405",
X"80cb0533",
X"71075452",
X"5e575956",
X"02b70533",
X"78712902",
X"8805b605",
X"33028c05",
X"b5053371",
X"882b0770",
X"1d707f8c",
X"050c5f59",
X"57595d8e",
X"3d33821b",
X"3402b905",
X"33903d33",
X"71882b07",
X"5a5c7884",
X"1b2302bb",
X"05330284",
X"05ba0533",
X"71882b07",
X"565c74ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"07515253",
X"575e5c74",
X"76317831",
X"79842a90",
X"3d335471",
X"71315356",
X"5680d0bb",
X"3f83c080",
X"08820570",
X"881c0c83",
X"c08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83c0900c",
X"80567583",
X"c0800c97",
X"3d0d04e9",
X"3d0d83c0",
X"90085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e53f83c0",
X"80085483",
X"c0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f489",
X"3f83c080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383c080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83c09008",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0e93f",
X"83c08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"833f83c0",
X"80085583",
X"c0800880",
X"2eff8938",
X"83c08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"519ad63f",
X"83c08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83c0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83c09008",
X"55568555",
X"73802e81",
X"e3388114",
X"33810653",
X"84557280",
X"2e81d538",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b9388214",
X"3370892b",
X"56537680",
X"2eb73874",
X"52ff1651",
X"80cbbc3f",
X"83c08008",
X"ff187654",
X"70535853",
X"80cbac3f",
X"83c08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed63f83",
X"c0800853",
X"810b83c0",
X"8008278b",
X"38881408",
X"83c08008",
X"26883880",
X"0b811534",
X"b03983c0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc53f",
X"83c08008",
X"8c3883c0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683c0",
X"800805a8",
X"150c8055",
X"7483c080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83c09008",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1cf3f",
X"83c08008",
X"5583c080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef5",
X"3f83c080",
X"0888170c",
X"7551efa6",
X"3f83c080",
X"08557483",
X"c0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683c0",
X"9008802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f53f83c0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"96df3f83",
X"c0800841",
X"83c08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"eddf3f83",
X"c0800841",
X"83c08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"8e853f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f03f83c0",
X"80088332",
X"70307072",
X"079f2c83",
X"c0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"8c913f75",
X"83c0800c",
X"9e3d0d04",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"7751e0d2",
X"3f83c080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3381dad0",
X"0b81dad0",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"527751e0",
X"813f83c0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583c0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"558b983f",
X"83c08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"8114518a",
X"b03f83c0",
X"80083070",
X"83c08008",
X"07802583",
X"c0800c53",
X"863d0d04",
X"fc3d0d76",
X"705255e6",
X"ee3f83c0",
X"80085481",
X"5383c080",
X"0880c138",
X"7451e6b1",
X"3f83c080",
X"0881d8cc",
X"5383c080",
X"085253ff",
X"913f83c0",
X"8008a138",
X"81d8d052",
X"7251ff82",
X"3f83c080",
X"08923881",
X"d8d45272",
X"51fef33f",
X"83c08008",
X"802e8338",
X"81547353",
X"7283c080",
X"0c863d0d",
X"04fd3d0d",
X"75705254",
X"e68d3f81",
X"5383c080",
X"08983873",
X"51e5d63f",
X"83c39808",
X"5283c080",
X"0851feba",
X"3f83c080",
X"08537283",
X"c0800c85",
X"3d0d04df",
X"3d0da43d",
X"0870525e",
X"dbfb3f83",
X"c0800833",
X"953d5654",
X"73963881",
X"dde05274",
X"5189903f",
X"9a397d52",
X"7851defc",
X"3f84cf39",
X"7d51dbe1",
X"3f83c080",
X"08527451",
X"db913f80",
X"43804280",
X"41804083",
X"c3a00852",
X"943d7052",
X"5de1e43f",
X"83c08008",
X"59800b83",
X"c0800855",
X"5b83c080",
X"087b2e94",
X"38811b74",
X"525be4e6",
X"3f83c080",
X"085483c0",
X"8008ee38",
X"805aff5f",
X"7909709f",
X"2c7b065b",
X"547a7a24",
X"8438ff1b",
X"5af61a70",
X"09709f2c",
X"72067bff",
X"125a5a52",
X"55558075",
X"25953876",
X"51e4ab3f",
X"83c08008",
X"76ff1858",
X"55577380",
X"24ed3874",
X"7f2e8638",
X"a0d83f74",
X"5f78ff1b",
X"70585d58",
X"807a2595",
X"387751e4",
X"813f83c0",
X"800876ff",
X"18585558",
X"738024ed",
X"38800b83",
X"c7d00c80",
X"0b83c894",
X"0c81d8d8",
X"518d8f3f",
X"81800b83",
X"c8940c81",
X"d8e0518d",
X"813fa80b",
X"83c7d00c",
X"76802e80",
X"e43883c7",
X"d0087779",
X"32703070",
X"72078025",
X"70872b83",
X"c8940c51",
X"56785356",
X"56e3b83f",
X"83c08008",
X"802e8838",
X"81d8e851",
X"8cc83f76",
X"51e2fa3f",
X"83c08008",
X"5281d9f4",
X"518cb73f",
X"7651e382",
X"3f83c080",
X"0883c7d0",
X"08555775",
X"74258638",
X"a81656f7",
X"397583c7",
X"d00c86f0",
X"7624ff98",
X"3887980b",
X"83c7d00c",
X"77802eb1",
X"387751e2",
X"b83f83c0",
X"80087852",
X"55e2d83f",
X"81d8f054",
X"83c08008",
X"8d388739",
X"80763481",
X"d03981d8",
X"ec547453",
X"735281d8",
X"c0518bd6",
X"3f805481",
X"d8c8518b",
X"cd3f8114",
X"5473a82e",
X"098106ef",
X"38868da0",
X"519cdd3f",
X"8052903d",
X"70525780",
X"c19e3f83",
X"52765180",
X"c1963f62",
X"818f3861",
X"802e80fb",
X"387b5473",
X"ff2e9638",
X"78802e81",
X"89387851",
X"e1dc3f83",
X"c08008ff",
X"155559e7",
X"3978802e",
X"80f43878",
X"51e1d83f",
X"83c08008",
X"802efc8e",
X"387851e1",
X"a03f83c0",
X"80085281",
X"d8bc5183",
X"e33f83c0",
X"8008a338",
X"7c51859b",
X"3f83c080",
X"085574ff",
X"16565480",
X"7425ae38",
X"741d7033",
X"555673af",
X"2efecd38",
X"e9397851",
X"e0e13f83",
X"c0800852",
X"7c5184d3",
X"3f8f397f",
X"88296010",
X"057a0561",
X"055afc90",
X"3962802e",
X"fbd13880",
X"527651bf",
X"f73fa33d",
X"0d04803d",
X"0d9088b8",
X"337081ff",
X"0670842a",
X"81327081",
X"06515151",
X"5170802e",
X"8d38a80b",
X"9088b834",
X"b80b9088",
X"b8347083",
X"c0800c82",
X"3d0d0480",
X"3d0d9088",
X"b8337081",
X"ff067085",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d3898",
X"0b9088b8",
X"34b80b90",
X"88b83470",
X"83c0800c",
X"823d0d04",
X"930b9088",
X"bc34ff0b",
X"9088a834",
X"04ff3d0d",
X"028f0533",
X"52800b90",
X"88bc348a",
X"519aa53f",
X"df3f80f8",
X"0b9088a0",
X"34800b90",
X"888834fa",
X"12527190",
X"88803480",
X"0b908898",
X"34719088",
X"90349088",
X"b8528072",
X"34b87234",
X"833d0d04",
X"803d0d02",
X"8b053351",
X"709088b4",
X"34febf3f",
X"83c08008",
X"802ef638",
X"823d0d04",
X"803d0d84",
X"39a3fe3f",
X"fed93f83",
X"c0800880",
X"2ef33890",
X"88b43370",
X"81ff0683",
X"c0800c51",
X"823d0d04",
X"803d0da3",
X"0b9088bc",
X"34ff0b90",
X"88a83490",
X"88b851a8",
X"7134b871",
X"34823d0d",
X"04803d0d",
X"9088bc33",
X"7081c006",
X"70307080",
X"2583c080",
X"0c515151",
X"823d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"832a8132",
X"70810651",
X"51515170",
X"802ee838",
X"b00b9088",
X"b834b80b",
X"9088b834",
X"823d0d04",
X"803d0d90",
X"80ac0881",
X"0683c080",
X"0c823d0d",
X"04fd3d0d",
X"75775454",
X"80732594",
X"38737081",
X"05553352",
X"81d8f451",
X"87843fff",
X"1353e939",
X"853d0d04",
X"fd3d0d75",
X"77535473",
X"33517089",
X"38713351",
X"70802ea1",
X"38733372",
X"33525372",
X"71278538",
X"ff519439",
X"70732785",
X"3881518b",
X"39811481",
X"135354d3",
X"39805170",
X"83c0800c",
X"853d0d04",
X"fd3d0d75",
X"77545472",
X"337081ff",
X"06525270",
X"802ea338",
X"7181ff06",
X"8114ffbf",
X"12535452",
X"70992689",
X"38a01270",
X"81ff0653",
X"51717470",
X"81055634",
X"d2398074",
X"34853d0d",
X"04ffbd3d",
X"0d80c63d",
X"0852a53d",
X"705254ff",
X"b33f80c7",
X"3d085285",
X"3d705253",
X"ffa63f72",
X"527351fe",
X"df3f80c5",
X"3d0d04fe",
X"3d0d7476",
X"53537170",
X"81055333",
X"51707370",
X"81055534",
X"70f03884",
X"3d0d04fe",
X"3d0d7452",
X"80723352",
X"5370732e",
X"8d388112",
X"81147133",
X"53545270",
X"f5387283",
X"c0800c84",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"b8913f83",
X"c080087a",
X"27ee3874",
X"802e80dd",
X"38745275",
X"51b7fc3f",
X"83c08008",
X"75537652",
X"54b8803f",
X"83c08008",
X"7a537552",
X"56b7e43f",
X"83c08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"c08008c5",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9f",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fc813f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd53f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbb13f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83c0940c",
X"7183c098",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383c094",
X"085283c0",
X"980851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"bdba5351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fc3d",
X"0d765574",
X"83c3a808",
X"2eaf3880",
X"53745187",
X"c13f83c0",
X"800881ff",
X"06ff1470",
X"81ff0672",
X"30709f2a",
X"51525553",
X"5472802e",
X"843871dd",
X"3873fe38",
X"7483c3a8",
X"0c863d0d",
X"04ff3d0d",
X"ff0b83c3",
X"a80c84a5",
X"3f815187",
X"853f83c0",
X"800881ff",
X"065271ee",
X"3881d33f",
X"7183c080",
X"0c833d0d",
X"04fc3d0d",
X"76028405",
X"a2052202",
X"8805a605",
X"227a5455",
X"5555ff82",
X"3f72802e",
X"a03883c3",
X"bc143375",
X"70810557",
X"34811470",
X"83ffff06",
X"ff157083",
X"ffff0656",
X"525552dd",
X"39800b83",
X"c0800c86",
X"3d0d04fc",
X"3d0d7678",
X"7a115653",
X"55805371",
X"742e9338",
X"72155170",
X"3383c3bc",
X"13348112",
X"81145452",
X"ea39800b",
X"83c0800c",
X"863d0d04",
X"fd3d0d90",
X"5483c3a8",
X"085186f4",
X"3f83c080",
X"0881ff06",
X"ff157130",
X"71307073",
X"079f2a72",
X"9f2a0652",
X"55525553",
X"72db3885",
X"3d0d0480",
X"3d0d83c3",
X"b4081083",
X"c3ac0807",
X"9080a80c",
X"823d0d04",
X"800b83c3",
X"b40ce43f",
X"04810b83",
X"c3b40cdb",
X"3f04ed3f",
X"047183c3",
X"b00c0480",
X"3d0d8051",
X"f43f810b",
X"83c3b40c",
X"810b83c3",
X"ac0cffbb",
X"3f823d0d",
X"04803d0d",
X"72307074",
X"07802583",
X"c3ac0c51",
X"ffa53f82",
X"3d0d0480",
X"3d0d028b",
X"05339080",
X"a40c9080",
X"a8087081",
X"06515170",
X"f5389080",
X"a4087081",
X"ff0683c0",
X"800c5182",
X"3d0d0480",
X"3d0d81ff",
X"51d13f83",
X"c0800881",
X"ff0683c0",
X"800c823d",
X"0d04803d",
X"0d73902b",
X"73079080",
X"b40c823d",
X"0d0404fb",
X"3d0d7802",
X"84059f05",
X"3370982b",
X"55575572",
X"80259b38",
X"7580ff06",
X"56805280",
X"f751e03f",
X"83c08008",
X"81ff0654",
X"73812680",
X"ff388051",
X"fee73fff",
X"a23f8151",
X"fedf3fff",
X"9a3f7551",
X"feed3f74",
X"982a51fe",
X"e63f7490",
X"2a7081ff",
X"065253fe",
X"da3f7488",
X"2a7081ff",
X"065253fe",
X"ce3f7481",
X"ff0651fe",
X"c63f8155",
X"7580c02e",
X"09810686",
X"38819555",
X"8d397580",
X"c82e0981",
X"06843881",
X"87557451",
X"fea53f8a",
X"55fec83f",
X"83c08008",
X"81ff0670",
X"982b5454",
X"7280258c",
X"38ff1570",
X"81ff0656",
X"5374e238",
X"7383c080",
X"0c873d0d",
X"04fa3d0d",
X"fdc53f80",
X"51fdda3f",
X"8a54fe93",
X"3fff1470",
X"81ff0655",
X"5373f338",
X"73745355",
X"80c051fe",
X"a63f83c0",
X"800881ff",
X"06547381",
X"2e098106",
X"829f3883",
X"aa5280c8",
X"51fe8c3f",
X"83c08008",
X"81ff0653",
X"72812e09",
X"810681a8",
X"38745487",
X"3d741154",
X"56fdc83f",
X"83c08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e53802",
X"9a053353",
X"72812e09",
X"810681d9",
X"38029b05",
X"335380ce",
X"90547281",
X"aa2e8d38",
X"81c73980",
X"e4518acc",
X"3fff1454",
X"73802e81",
X"b838820a",
X"5281e951",
X"fda53f83",
X"c0800881",
X"ff065372",
X"de387252",
X"80fa51fd",
X"923f83c0",
X"800881ff",
X"06537281",
X"90387254",
X"731653fc",
X"d63f83c0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e8",
X"38873d33",
X"70862a70",
X"81065154",
X"548c5572",
X"80e33884",
X"5580de39",
X"745281e9",
X"51fccc3f",
X"83c08008",
X"81ff0653",
X"825581e9",
X"56817327",
X"86387355",
X"80c15680",
X"ce90548a",
X"3980e451",
X"89be3fff",
X"14547380",
X"2ea93880",
X"527551fc",
X"9a3f83c0",
X"800881ff",
X"065372e1",
X"38848052",
X"80d051fc",
X"863f83c0",
X"800881ff",
X"06537280",
X"2e833880",
X"557483c3",
X"b8348051",
X"fb873ffb",
X"c23f883d",
X"0d04fb3d",
X"0d775480",
X"0b83c3b8",
X"3370832a",
X"70810651",
X"55575572",
X"752e0981",
X"06853873",
X"892b5473",
X"5280d151",
X"fbbd3f83",
X"c0800881",
X"ff065372",
X"bd3882b8",
X"c054fb83",
X"3f83c080",
X"0881ff06",
X"537281ff",
X"2e098106",
X"8938ff14",
X"5473e738",
X"9f397281",
X"fe2e0981",
X"06963883",
X"c7bc5283",
X"c3bc51fa",
X"ed3ffad3",
X"3ffad03f",
X"83398155",
X"8051fa89",
X"3ffac43f",
X"7481ff06",
X"83c0800c",
X"873d0d04",
X"fb3d0d77",
X"83c3bc56",
X"548151f9",
X"ec3f83c3",
X"b8337083",
X"2a708106",
X"51545672",
X"85387389",
X"2b547352",
X"80d851fa",
X"b63f83c0",
X"800881ff",
X"06537280",
X"e43881ff",
X"51f9d43f",
X"81fe51f9",
X"ce3f8480",
X"53747081",
X"05563351",
X"f9c13fff",
X"137083ff",
X"ff065153",
X"72eb3872",
X"51f9b03f",
X"7251f9ab",
X"3ff9d03f",
X"83c08008",
X"9f0653a7",
X"88547285",
X"2e8c3899",
X"3980e451",
X"86f63fff",
X"1454f9b3",
X"3f83c080",
X"0881ff2e",
X"843873e9",
X"388051f8",
X"e43ff99f",
X"3f800b83",
X"c0800c87",
X"3d0d0471",
X"83c7c00c",
X"8880800b",
X"83c7bc0c",
X"8480800b",
X"83c7c40c",
X"04fd3d0d",
X"77701755",
X"7705ff1a",
X"535371ff",
X"2e943873",
X"70810555",
X"33517073",
X"70810555",
X"34ff1252",
X"e939853d",
X"0d04fc3d",
X"0d87a681",
X"55743383",
X"c7c834a0",
X"5483a080",
X"5383c7c0",
X"085283c7",
X"bc0851ff",
X"b83fa054",
X"83a48053",
X"83c7c008",
X"5283c7bc",
X"0851ffa5",
X"3f905483",
X"a8805383",
X"c7c00852",
X"83c7bc08",
X"51ff923f",
X"a0538052",
X"83c7c408",
X"83a08005",
X"5185ce3f",
X"a0538052",
X"83c7c408",
X"83a48005",
X"5185be3f",
X"90538052",
X"83c7c408",
X"83a88005",
X"5185ae3f",
X"ff753483",
X"a0805480",
X"5383c7c0",
X"085283c7",
X"c40851fe",
X"cc3f80d0",
X"805483b0",
X"805383c7",
X"c0085283",
X"c7c40851",
X"feb73f86",
X"e13fa254",
X"805383c7",
X"c4088c80",
X"055281db",
X"c451fea1",
X"3f860b87",
X"a8833480",
X"0b87a882",
X"34800b87",
X"a09a34af",
X"0b87a096",
X"34bf0b87",
X"a0973480",
X"0b87a098",
X"349f0b87",
X"a0993480",
X"0b87a09b",
X"34e00b87",
X"a88934a2",
X"0b87a880",
X"34830b87",
X"a48f3482",
X"0b87a881",
X"34863d0d",
X"04fd3d0d",
X"83a08054",
X"805383c7",
X"c4085283",
X"c7c00851",
X"fdbf3f80",
X"d0805483",
X"b0805383",
X"c7c40852",
X"83c7c008",
X"51fdaa3f",
X"a05483a0",
X"805383c7",
X"c4085283",
X"c7c00851",
X"fd973fa0",
X"5483a480",
X"5383c7c4",
X"085283c7",
X"c00851fd",
X"843f9054",
X"83a88053",
X"83c7c408",
X"5283c7c0",
X"0851fcf1",
X"3f83c7c8",
X"3387a681",
X"34853d0d",
X"04803d0d",
X"90809008",
X"810683c0",
X"800c823d",
X"0d04ff3d",
X"0d908090",
X"700870fe",
X"06760772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087081",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fd0676",
X"1007720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870822c",
X"bf0683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe830676",
X"822b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087088",
X"2c870683",
X"c0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70f1ff06",
X"76882b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"8b2cbf06",
X"83c0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f88f",
X"ff06768b",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870912c",
X"bf0683c0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fc87ffff",
X"0676912b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70992c81",
X"0683c080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870ff",
X"bf0a0676",
X"992b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"80087088",
X"2c810683",
X"c0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"892c8106",
X"83c0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708a2c81",
X"0683c080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708b2c",
X"810683c0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708c",
X"2cbf0683",
X"c0800c51",
X"823d0d04",
X"fe3d0d74",
X"81e62987",
X"2a9080a0",
X"0c843d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727081",
X"055434ff",
X"1151f039",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708405",
X"540cff11",
X"51f03984",
X"3d0d04fe",
X"3d0d8480",
X"80538052",
X"88800a51",
X"ffb33f81",
X"80805380",
X"5282800a",
X"51c63f84",
X"3d0d0480",
X"3d0d8151",
X"fbfc3f72",
X"802e9038",
X"8051fdfe",
X"3fcd3f83",
X"c7cc3351",
X"fdf43f81",
X"51fc8d3f",
X"8051fc88",
X"3f8051fb",
X"d93f823d",
X"0d04fd3d",
X"0d755280",
X"5480ff72",
X"25883881",
X"0bff8013",
X"5354ffbf",
X"12517099",
X"268638e0",
X"12529e39",
X"ff9f1251",
X"99712795",
X"38d012e0",
X"13705454",
X"51897127",
X"88388f73",
X"27833880",
X"5273802e",
X"85388180",
X"12527181",
X"ff0683c0",
X"800c853d",
X"0d04803d",
X"0d84d8c0",
X"51807170",
X"81055334",
X"7084e0c0",
X"2e098106",
X"f038823d",
X"0d04fe3d",
X"0d029705",
X"3351ff86",
X"3f83c080",
X"0881ff06",
X"83c7d008",
X"54528073",
X"249b3883",
X"c8900813",
X"7283c894",
X"08075353",
X"71733483",
X"c7d00881",
X"0583c7d0",
X"0c843d0d",
X"04fa3d0d",
X"82800a1b",
X"55805788",
X"3dfc0554",
X"79537452",
X"7851ffbb",
X"893f883d",
X"0d04fe3d",
X"0d83c7e8",
X"08527451",
X"c1ed3f83",
X"c080088c",
X"38765375",
X"5283c7e8",
X"0851c63f",
X"843d0d04",
X"fe3d0d83",
X"c7e80853",
X"75527451",
X"ffbcab3f",
X"83c08008",
X"8d387753",
X"765283c7",
X"e80851ff",
X"a03f843d",
X"0d04fe3d",
X"0d83c7e8",
X"0851ffbb",
X"9e3f83c0",
X"80088180",
X"802e0981",
X"06883883",
X"c1808053",
X"9c3983c7",
X"e80851ff",
X"bb813f83",
X"c0800880",
X"d0802e09",
X"81069338",
X"83c1b080",
X"5383c080",
X"085283c7",
X"e80851fe",
X"d43f843d",
X"0d04803d",
X"0df9e03f",
X"83c08008",
X"842981db",
X"e8057008",
X"83c0800c",
X"51823d0d",
X"04ed3d0d",
X"80448043",
X"80428041",
X"80705a5b",
X"fdcc3f80",
X"0b83c7d0",
X"0c800b83",
X"c8940c81",
X"d9c051ea",
X"a53f8180",
X"0b83c894",
X"0c81d9c4",
X"51ea973f",
X"80d00b83",
X"c7d00c78",
X"30707a07",
X"80257087",
X"2b83c894",
X"0c5155f8",
X"d13f83c0",
X"80085281",
X"d9cc51e9",
X"f13f80f8",
X"0b83c7d0",
X"0c788132",
X"70307072",
X"07802570",
X"872b83c8",
X"940c5156",
X"56feef3f",
X"83c08008",
X"5281d9d8",
X"51e9c73f",
X"81a00b83",
X"c7d00c78",
X"82327030",
X"70720780",
X"2570872b",
X"83c8940c",
X"515683c7",
X"e8085256",
X"ffb6a63f",
X"83c08008",
X"5281d9e0",
X"51e9973f",
X"81f00b83",
X"c7d00c81",
X"0b83c7d4",
X"5b5883c7",
X"d0088219",
X"7a327030",
X"70720780",
X"2570872b",
X"83c8940c",
X"51578e3d",
X"7055ff1b",
X"54575757",
X"9a8f3f79",
X"7084055b",
X"0851ffb5",
X"dc3f7454",
X"83c08008",
X"53775281",
X"d9e851e8",
X"c93fa817",
X"83c7d00c",
X"81185877",
X"852e0981",
X"06ffaf38",
X"83900b83",
X"c7d00c78",
X"87327030",
X"70720780",
X"2570872b",
X"83c8940c",
X"515656f7",
X"f53f81d9",
X"f85583c0",
X"8008802e",
X"8f3883c7",
X"e40851ff",
X"b5873f83",
X"c0800855",
X"745281da",
X"8051e7f6",
X"3f83e00b",
X"83c7d00c",
X"78883270",
X"30707207",
X"80257087",
X"2b83c894",
X"0c515781",
X"da8c5255",
X"e7d43f86",
X"8da051f8",
X"ef3f8052",
X"913d7052",
X"559db13f",
X"83527451",
X"9daa3f63",
X"557482fa",
X"38611959",
X"78802585",
X"38745990",
X"39887925",
X"85388859",
X"87397888",
X"2682d938",
X"78822b55",
X"81d4c415",
X"0804f5e2",
X"3f83c080",
X"08615755",
X"75812e09",
X"81068938",
X"83c08008",
X"10559039",
X"75ff2e09",
X"81068838",
X"83c08008",
X"812c5590",
X"75258538",
X"90558839",
X"74802483",
X"38815574",
X"51f5bc3f",
X"828e39f5",
X"ce3f83c0",
X"80086105",
X"55748025",
X"85388055",
X"88398775",
X"25833887",
X"557451f5",
X"c73f81ec",
X"39608738",
X"62802e81",
X"e33883c3",
X"9c0883c3",
X"980cade5",
X"0b83c3a0",
X"0c83c7e8",
X"0851d78b",
X"3ffadb3f",
X"81c63960",
X"56807625",
X"9838ad84",
X"0b83c3a0",
X"0c83c7c8",
X"15700852",
X"55d6ec3f",
X"74085292",
X"39758025",
X"923883c7",
X"c8150851",
X"ffb2f03f",
X"8052fd19",
X"51b83962",
X"802e818c",
X"3883c7c8",
X"15700883",
X"c7d40872",
X"0c83c7d4",
X"0cfd1a70",
X"5351558c",
X"953f83c0",
X"80085680",
X"518c8b3f",
X"83c08008",
X"52745188",
X"a23f7552",
X"8051889b",
X"3f80d539",
X"60558075",
X"25b63883",
X"c3a40883",
X"c3980cad",
X"e50b83c3",
X"a00c83c7",
X"e40851d5",
X"f63f83c7",
X"e40851d3",
X"973f83c0",
X"800881ff",
X"06705255",
X"f4d53f74",
X"802e9d38",
X"8155a139",
X"74802594",
X"3883c7e4",
X"0851ffb1",
X"e23f8051",
X"f4b93f84",
X"39628738",
X"7a802efa",
X"83388055",
X"7483c080",
X"0c953d0d",
X"04fe3d0d",
X"83c88051",
X"80f3d03f",
X"83c7f051",
X"80f3c83f",
X"f4d53f83",
X"c0800880",
X"2e863880",
X"51818a39",
X"f4da3f83",
X"c0800880",
X"fe38f4fa",
X"3f83c080",
X"08802eb9",
X"388151f2",
X"893f8051",
X"f4903fee",
X"fd3f800b",
X"83c7d00c",
X"f99b3f83",
X"c0800853",
X"ff0b83c7",
X"d00cf0e9",
X"3f7280cb",
X"3883c7cc",
X"3351f3ea",
X"3f7251f1",
X"d93f80c0",
X"39f4a23f",
X"83c08008",
X"802eb538",
X"8151f1c6",
X"3f8051f3",
X"cd3feeba",
X"3fad840b",
X"83c3a00c",
X"83c7d408",
X"51d4983f",
X"ff0b83c7",
X"d00cf0a5",
X"3f83c7d4",
X"08528051",
X"86893f81",
X"51f5943f",
X"843d0d04",
X"fb3d0d80",
X"5283c880",
X"5180e2d7",
X"3f815283",
X"c7f05180",
X"e2cd3f80",
X"0b83c7cc",
X"34908080",
X"52868480",
X"8051ffb3",
X"f73f83c0",
X"80088197",
X"3889c03f",
X"81ddc851",
X"ffb8b63f",
X"83c08008",
X"559c800a",
X"5480c080",
X"5381da94",
X"5283c080",
X"0851f6d4",
X"3f83c7e8",
X"085381da",
X"a4527451",
X"ffb2ff3f",
X"83c08008",
X"8438f6e2",
X"3f83c7ec",
X"085381da",
X"b0527451",
X"ffb2e73f",
X"83c08008",
X"b638873d",
X"fc055484",
X"80805386",
X"a8808052",
X"83c7ec08",
X"51ffb0f2",
X"3f83c080",
X"08933875",
X"8480802e",
X"09810689",
X"38810b83",
X"c7cc3487",
X"39800b83",
X"c7cc3483",
X"c7cc3351",
X"f1e03f81",
X"51f3cc3f",
X"92de3f81",
X"51f3c43f",
X"8151fcfd",
X"3ffa3983",
X"c08c0802",
X"83c08c0c",
X"fb3d0d02",
X"81dabc0b",
X"83c39c0c",
X"81dac00b",
X"83c3940c",
X"81dac40b",
X"83c3a40c",
X"83c08c08",
X"fc050c80",
X"0b83c7d4",
X"0b83c08c",
X"08f8050c",
X"83c08c08",
X"f4050cff",
X"b1823f83",
X"c0800886",
X"05fc0683",
X"c08c08f0",
X"050c0283",
X"c08c08f0",
X"0508310d",
X"833d7083",
X"c08c08f8",
X"05087084",
X"0583c08c",
X"08f8050c",
X"0c51ffad",
X"ca3f83c0",
X"8c08f405",
X"08810583",
X"c08c08f4",
X"050c83c0",
X"8c08f405",
X"08872e09",
X"8106ffab",
X"38869480",
X"8051eadf",
X"3fff0b83",
X"c7d00c80",
X"0b83c894",
X"0c84d8c0",
X"0b83c890",
X"0c8151ee",
X"893f8151",
X"eeae3f80",
X"51eea93f",
X"8151eecf",
X"3f8151ef",
X"a43f8251",
X"eef23f80",
X"51efc83f",
X"8051eff2",
X"3f80d0ca",
X"528051df",
X"be3ffcc8",
X"3f83c08c",
X"08fc0508",
X"0d800b83",
X"c0800c87",
X"3d0d83c0",
X"8c0c0480",
X"3d0d81ff",
X"51800b83",
X"c8a01234",
X"ff115170",
X"f438823d",
X"0d04ff3d",
X"0d737033",
X"53518111",
X"33713471",
X"81123483",
X"3d0d04fb",
X"3d0d7779",
X"56568070",
X"71555552",
X"717525ac",
X"38721670",
X"33701470",
X"81ff0655",
X"51515171",
X"74278938",
X"81127081",
X"ff065351",
X"71811470",
X"83ffff06",
X"55525474",
X"7324d638",
X"7183c080",
X"0c873d0d",
X"04fb3d0d",
X"7756d788",
X"3f83c080",
X"08802ef6",
X"3883cabc",
X"08860570",
X"81ff0652",
X"53d58a3f",
X"810b9088",
X"d4349088",
X"d4337081",
X"ff065153",
X"728638f9",
X"d83fef39",
X"80557416",
X"75822b54",
X"549088c0",
X"13337434",
X"81155574",
X"852e0981",
X"06e83881",
X"0b9088d4",
X"34753383",
X"c8a03481",
X"163383c8",
X"a1348216",
X"3383c8a2",
X"34831633",
X"83c8a334",
X"845283c8",
X"a051febf",
X"3f83c080",
X"0881ff06",
X"84173357",
X"5372762e",
X"0981068c",
X"38d5b63f",
X"83c08008",
X"802e9a38",
X"83cabc08",
X"a82e0981",
X"06893886",
X"0b83cabc",
X"0c8739a8",
X"0b83cabc",
X"0c80e451",
X"eea63f87",
X"3d0d04f4",
X"3d0d7e60",
X"5955805d",
X"8075822b",
X"7183cac0",
X"120c83ca",
X"d4175b5b",
X"57767934",
X"77772e83",
X"b9387652",
X"7751ffac",
X"953f8e3d",
X"fc055490",
X"5383caa8",
X"527751ff",
X"abd03f7c",
X"5675902e",
X"09810683",
X"953883ca",
X"a851fd9a",
X"3f83caaa",
X"51fd933f",
X"83caac51",
X"fd8c3f76",
X"83cab80c",
X"7751ffa9",
X"9c3f0b0b",
X"81d8d052",
X"83c08008",
X"51cbb33f",
X"83c08008",
X"812e0981",
X"0680d438",
X"7683cad0",
X"0c820b83",
X"caa834ff",
X"960b83ca",
X"a9347751",
X"ffabe03f",
X"83c08008",
X"5583c080",
X"08772588",
X"3883c080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"caaa3474",
X"83caab34",
X"7683caac",
X"34ff800b",
X"83caad34",
X"81903983",
X"caa83383",
X"caa93371",
X"882b0756",
X"5b7483ff",
X"ff2e0981",
X"0680e838",
X"fe800b83",
X"cad00c81",
X"0b83cab8",
X"0cff0b83",
X"caa834ff",
X"0b83caa9",
X"347751ff",
X"aaed3f83",
X"c0800883",
X"cad80c83",
X"c0800855",
X"83c08008",
X"80258838",
X"83c08008",
X"8f055574",
X"842c7083",
X"ffff0670",
X"882a5851",
X"557583ca",
X"aa347483",
X"caab3476",
X"83caac34",
X"ff800b83",
X"caad3481",
X"0b83cab7",
X"34a53974",
X"85962e09",
X"810680fe",
X"387583ca",
X"d00c7751",
X"ffaaa13f",
X"83cab733",
X"83c08008",
X"07557483",
X"cab73483",
X"cab73381",
X"06557480",
X"2e833884",
X"5783caac",
X"3383caad",
X"3371882b",
X"07565c74",
X"81802e09",
X"8106a138",
X"83caaa33",
X"83caab33",
X"71882b07",
X"565bad80",
X"75278738",
X"76820757",
X"9c397681",
X"07579639",
X"7482802e",
X"09810687",
X"38768307",
X"57873974",
X"81ff268a",
X"387783ca",
X"c01b0c76",
X"79348e3d",
X"0d04803d",
X"0d728429",
X"83cac005",
X"700883c0",
X"800c5182",
X"3d0d04fe",
X"3d0d800b",
X"83caa40c",
X"800b83ca",
X"a00cff0b",
X"83c89c0c",
X"a80b83ca",
X"bc0cae51",
X"cfd73f80",
X"0b83cac0",
X"54528073",
X"70840555",
X"0c811252",
X"71842e09",
X"8106ef38",
X"843d0d04",
X"fe3d0d74",
X"02840596",
X"05225353",
X"71802e96",
X"38727081",
X"05543351",
X"cfe23fff",
X"127083ff",
X"ff065152",
X"e739843d",
X"0d04fe3d",
X"0d029205",
X"225382ac",
X"51e9b93f",
X"80c351cf",
X"bf3f8196",
X"51e9ad3f",
X"725283c8",
X"a051ffb4",
X"3f725283",
X"c8a051f8",
X"f63f83c0",
X"800881ff",
X"0651cf9c",
X"3f843d0d",
X"04ffb13d",
X"0d80d13d",
X"f80551f9",
X"a03f83ca",
X"a4088105",
X"83caa40c",
X"80cf3d33",
X"cf117081",
X"ff065156",
X"56748326",
X"88d73875",
X"8f06ff05",
X"567583c8",
X"9c082e9b",
X"38758326",
X"96387583",
X"c89c0c75",
X"842983ca",
X"c0057008",
X"53557551",
X"fa993f80",
X"762488b3",
X"38758429",
X"83cac005",
X"55740880",
X"2e88a438",
X"83c89c08",
X"842983ca",
X"c0057008",
X"02880582",
X"b9053352",
X"5b557480",
X"d22e84a7",
X"387480d2",
X"24903874",
X"bf2e9c38",
X"7480d02e",
X"81d13887",
X"e3397480",
X"d32e80cf",
X"387480d7",
X"2e81c038",
X"87d23902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"5656ce98",
X"3f80c151",
X"cdd23ff6",
X"f23f860b",
X"83c8a034",
X"815283c8",
X"a051cef5",
X"3f8151fd",
X"e93f7489",
X"38860b83",
X"cabc0c87",
X"39a80b83",
X"cabc0ccd",
X"e73f80c1",
X"51cda13f",
X"f6c13f90",
X"0b83cab7",
X"33810656",
X"5674802e",
X"83389856",
X"83caac33",
X"83caad33",
X"71882b07",
X"56597481",
X"802e0981",
X"069c3883",
X"caaa3383",
X"caab3371",
X"882b0756",
X"57ad8075",
X"278c3875",
X"81800756",
X"853975a0",
X"07567583",
X"c8a034ff",
X"0b83c8a1",
X"34e00b83",
X"c8a23480",
X"0b83c8a3",
X"34845283",
X"c8a051cd",
X"ec3f8451",
X"86903902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"5659ccdc",
X"3f7951ff",
X"a4f23f83",
X"c0800880",
X"2e8a3880",
X"ce51cc88",
X"3f85e639",
X"80c151cb",
X"ff3fccf4",
X"3fcba93f",
X"83cad008",
X"58837525",
X"9b3883ca",
X"ac3383ca",
X"ad337188",
X"2b07fc17",
X"71297a05",
X"8380055a",
X"51578d39",
X"74818029",
X"18ff8005",
X"58818057",
X"80567676",
X"2e9238cb",
X"db3f83c0",
X"800883c8",
X"a0173481",
X"1656eb39",
X"cbca3f83",
X"c0800881",
X"ff067753",
X"83c8a052",
X"56f4ec3f",
X"83c08008",
X"81ff0655",
X"75752e09",
X"81068190",
X"38cbc93f",
X"80c151cb",
X"833fcbf8",
X"3f775279",
X"51ffa38a",
X"3f805e80",
X"d13dfdf4",
X"05547653",
X"83c8a052",
X"7951ffa1",
X"973f0282",
X"b9053355",
X"81597480",
X"d72e0981",
X"0680c538",
X"77527951",
X"ffa2db3f",
X"80d13dfd",
X"f0055476",
X"538f3d70",
X"537a5258",
X"ffa2933f",
X"80567676",
X"2ea23875",
X"1883c8a0",
X"17337133",
X"70723270",
X"30708025",
X"70307f06",
X"811d5d5f",
X"51515152",
X"5b55db39",
X"82ac51e3",
X"fb3f7880",
X"2e863880",
X"c3518439",
X"80ce51c9",
X"f73fcaec",
X"3fc9a13f",
X"83d23902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"59558070",
X"5d59ca94",
X"3f80c151",
X"c9ce3f83",
X"cab80879",
X"2e82d638",
X"83cad808",
X"80fc0555",
X"80fd5274",
X"5185a03f",
X"83c08008",
X"5b778224",
X"b238ff18",
X"70872b83",
X"ffff8006",
X"81dc8805",
X"83c8a059",
X"57558180",
X"55757081",
X"05573377",
X"70810559",
X"34ff1570",
X"81ff0651",
X"5574ea38",
X"82853977",
X"82e82e81",
X"a3387782",
X"e92e0981",
X"0681aa38",
X"78587787",
X"32703070",
X"72078025",
X"7a8a3270",
X"30707207",
X"80257307",
X"53545a51",
X"57557580",
X"2e973878",
X"78269238",
X"a00b83c8",
X"a01a3481",
X"197081ff",
X"065a55eb",
X"39811870",
X"81ff0659",
X"558a7827",
X"ffbc388f",
X"5883c89b",
X"183383c8",
X"a01934ff",
X"187081ff",
X"06595577",
X"8426ea38",
X"9058800b",
X"83c8a019",
X"34811870",
X"81ff0670",
X"982b5259",
X"55748025",
X"e93880c6",
X"557a858f",
X"24843880",
X"c2557483",
X"c8a03480",
X"f10b83c8",
X"a334810b",
X"83c8a434",
X"7a83c8a1",
X"347a882c",
X"557483c8",
X"a23480cb",
X"3982f078",
X"2580c438",
X"7780fd29",
X"fd97d305",
X"527951ff",
X"9fbc3f80",
X"d13dfdec",
X"055480fd",
X"5383c8a0",
X"527951ff",
X"9ef43f7b",
X"81195956",
X"7580fc24",
X"83387858",
X"77882c55",
X"7483c99d",
X"347783c9",
X"9e347583",
X"c99f3481",
X"805980cc",
X"3983cad0",
X"08578378",
X"259b3883",
X"caac3383",
X"caad3371",
X"882b07fc",
X"1a712979",
X"05838005",
X"5951598d",
X"39778180",
X"2917ff80",
X"05578180",
X"59765279",
X"51ff9eca",
X"3f80d13d",
X"fdec0554",
X"785383c8",
X"a0527951",
X"ff9e833f",
X"7851f6ce",
X"3fc7953f",
X"c5ca3f8b",
X"3983caa0",
X"08810583",
X"caa00c80",
X"d13d0d04",
X"f6ef3ffc",
X"39fc3d0d",
X"76787184",
X"2983cac0",
X"05700851",
X"53535370",
X"9e3880ce",
X"723480cf",
X"0b811334",
X"80ce0b82",
X"133480c5",
X"0b831334",
X"70841334",
X"80e73983",
X"cad41333",
X"5480d272",
X"3473822a",
X"70810651",
X"5180cf53",
X"70843880",
X"d7537281",
X"1334a00b",
X"82133473",
X"83065170",
X"812e9e38",
X"70812488",
X"3870802e",
X"8f389f39",
X"70822e92",
X"3870832e",
X"92389339",
X"80d8558e",
X"3980d355",
X"893980cd",
X"55843980",
X"c4557483",
X"133480c4",
X"0b841334",
X"800b8513",
X"34863d0d",
X"04fc3d0d",
X"76785354",
X"81538055",
X"87397110",
X"73105452",
X"73722651",
X"72802ea7",
X"3870802e",
X"86387180",
X"25e83872",
X"802e9838",
X"71742689",
X"38737231",
X"75740756",
X"5472812a",
X"72812a53",
X"53e53973",
X"51788338",
X"74517083",
X"c0800c86",
X"3d0d04fe",
X"3d0d8053",
X"75527451",
X"ffa33f84",
X"3d0d04fe",
X"3d0d8153",
X"75527451",
X"ff933f84",
X"3d0d04fb",
X"3d0d7779",
X"55558056",
X"74762586",
X"38743055",
X"81567380",
X"25883873",
X"30768132",
X"57548053",
X"73527451",
X"fee73f83",
X"c0800854",
X"75802e87",
X"3883c080",
X"08305473",
X"83c0800c",
X"873d0d04",
X"fa3d0d78",
X"7a575580",
X"57747725",
X"86387430",
X"55815775",
X"9f2c5481",
X"53757432",
X"74315274",
X"51feaa3f",
X"83c08008",
X"5476802e",
X"873883c0",
X"80083054",
X"7383c080",
X"0c883d0d",
X"04fc3d0d",
X"76558075",
X"0c800b84",
X"160c800b",
X"88160c80",
X"0b8c160c",
X"83c88051",
X"80dad43f",
X"83c7f051",
X"80dacc3f",
X"87a68033",
X"7081ff06",
X"5152dca3",
X"3f71812a",
X"81327281",
X"32718106",
X"71810631",
X"84180c54",
X"5471832a",
X"81327282",
X"2a813271",
X"81067181",
X"0631770c",
X"535387a0",
X"90337009",
X"81068817",
X"0c5283c0",
X"8008802e",
X"80c23883",
X"c0800881",
X"2a708106",
X"83c08008",
X"81063184",
X"170c5283",
X"c0800883",
X"2a83c080",
X"08822a71",
X"81067181",
X"0631770c",
X"535383c0",
X"8008842a",
X"81068816",
X"0c83c080",
X"08852a81",
X"068c160c",
X"863d0d04",
X"fe3d0d74",
X"76545271",
X"51febe3f",
X"72812ea2",
X"38817326",
X"8d387282",
X"2ea83872",
X"832e9c38",
X"e6397108",
X"e2388412",
X"08dd3888",
X"1208d838",
X"a5398812",
X"08812e9e",
X"38913988",
X"1208812e",
X"95387108",
X"91388412",
X"088c388c",
X"1208812e",
X"098106ff",
X"b238843d",
X"0d04fb3d",
X"0d780284",
X"059f0533",
X"5556800b",
X"81d6d456",
X"5381732b",
X"74065271",
X"802e8338",
X"81527470",
X"82055622",
X"7073902b",
X"0790809c",
X"0c518113",
X"5372882e",
X"098106d9",
X"38805383",
X"cae01333",
X"517081ff",
X"2eb23870",
X"1081d4f4",
X"05702255",
X"51807317",
X"70337010",
X"81d4f405",
X"70225151",
X"51525273",
X"712e9138",
X"81125271",
X"862e0981",
X"06f13873",
X"90809c0c",
X"81135372",
X"862e0981",
X"06ffb838",
X"80537216",
X"70335151",
X"7081ff2e",
X"94387010",
X"81d4f405",
X"70227084",
X"80800790",
X"809c0c51",
X"51811353",
X"72862e09",
X"8106d738",
X"80537216",
X"51703383",
X"cae01434",
X"81135372",
X"862e0981",
X"06ec3887",
X"3d0d0404",
X"ff3d0d74",
X"0284058f",
X"05335252",
X"70883871",
X"9080940c",
X"8e397081",
X"2e098106",
X"86387190",
X"80980c83",
X"3d0d04fb",
X"3d0d029f",
X"05337998",
X"2b70982c",
X"7c982b70",
X"982c83ca",
X"fc157033",
X"70982b70",
X"982c5158",
X"5c5a5155",
X"51545470",
X"732e0981",
X"06943883",
X"cadc1433",
X"70982b70",
X"982c5152",
X"5670722e",
X"b1387275",
X"347183ca",
X"dc153483",
X"cadd3383",
X"cafd3371",
X"982b7190",
X"2b0783ca",
X"dc337088",
X"2b720783",
X"cafc3371",
X"079080b8",
X"0c525953",
X"5452873d",
X"0d04fe3d",
X"0d748111",
X"33713371",
X"882b0783",
X"c0800c53",
X"51843d0d",
X"0483cae8",
X"3383c080",
X"0c04f53d",
X"0d02bb05",
X"33028405",
X"bf053302",
X"880580c3",
X"0533028c",
X"0580c605",
X"22665c5a",
X"5e5c567a",
X"557b5489",
X"53a1527d",
X"5180d0c0",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8d3d0d04",
X"83c08c08",
X"0283c08c",
X"0cf53d0d",
X"83c08c08",
X"88050883",
X"c08c088f",
X"053383c0",
X"8c089205",
X"22028c05",
X"73900583",
X"c08c08e8",
X"050c83c0",
X"8c08f805",
X"0c83c08c",
X"08f0050c",
X"83c08c08",
X"ec050c83",
X"c08c08f4",
X"050c800b",
X"83c08c08",
X"f0050883",
X"c08c08e0",
X"050c83c0",
X"8c08fc05",
X"0c83c08c",
X"08f00508",
X"89278a38",
X"890b83c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"860587ff",
X"fc0683c0",
X"8c08e005",
X"0c0283c0",
X"8c08e005",
X"08310d85",
X"3d705583",
X"c08c08ec",
X"05085483",
X"c08c08f0",
X"05085383",
X"c08c08f4",
X"05085283",
X"c08c08e4",
X"050c80d9",
X"f23f83c0",
X"800881ff",
X"0683c08c",
X"08e40508",
X"83c08c08",
X"ec050c83",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08802e8c",
X"3883c08c",
X"08f80508",
X"0d89c839",
X"83c08c08",
X"f0050880",
X"2e89a638",
X"83c08c08",
X"ec050881",
X"053383c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"842ea938",
X"840b83c0",
X"8c08e005",
X"082588c7",
X"3883c08c",
X"08e00508",
X"852e859b",
X"3883c08c",
X"08e00508",
X"a12e87ad",
X"3888ac39",
X"800b83c0",
X"8c08ec05",
X"08850533",
X"83c08c08",
X"e0050c83",
X"c08c08fc",
X"050c83c0",
X"8c08e005",
X"08832e09",
X"81068883",
X"3883c08c",
X"08e80508",
X"81053383",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08812687",
X"e638810b",
X"83c08c08",
X"e0050880",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08fc050c",
X"83c08c08",
X"ec050882",
X"053383c0",
X"8c08e005",
X"08870534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088b0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08e005",
X"088c0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088d0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"800b83c0",
X"8c08e005",
X"088e0523",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"800b83c0",
X"8c08e005",
X"088a0534",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"08057094",
X"0508fcff",
X"ff067194",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08ec0508",
X"86053383",
X"c08c08e0",
X"050c83c0",
X"8c08f405",
X"0c83c08c",
X"08e00508",
X"83c08c08",
X"fc05082e",
X"098106b6",
X"3883c08c",
X"08e80508",
X"81053370",
X"80d82983",
X"c08c08e8",
X"05080583",
X"c08c08e0",
X"050c83c0",
X"8c08e405",
X"0c83c08c",
X"08fc0508",
X"83c08c08",
X"e005088b",
X"053483c0",
X"8c08ec05",
X"08870533",
X"83c08c08",
X"e0050c83",
X"c08c08e0",
X"0508812e",
X"8f3883c0",
X"8c08e005",
X"08822eb7",
X"38848c39",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"820b83c0",
X"8c08e005",
X"088a0534",
X"83d93983",
X"c08c08e8",
X"05088105",
X"337080d8",
X"2983c08c",
X"08e80508",
X"0583c08c",
X"08e0050c",
X"83c08c08",
X"e4050c83",
X"c08c08fc",
X"050883c0",
X"8c08e005",
X"088a0534",
X"83a13983",
X"c08c08fc",
X"0508802e",
X"83953883",
X"c08c08ec",
X"05088305",
X"33830683",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08832e09",
X"810682f3",
X"3883c08c",
X"08ec0508",
X"82053370",
X"982b83c0",
X"8c08e005",
X"0c83c08c",
X"08e4050c",
X"83c08c08",
X"e0050880",
X"2582cc38",
X"83c08c08",
X"e8050881",
X"05337080",
X"d82983c0",
X"8c08e805",
X"080583c0",
X"8c08e005",
X"0c83c08c",
X"08f4050c",
X"83c08c08",
X"ec050886",
X"053383c0",
X"8c08e005",
X"0880d605",
X"3483c08c",
X"08e00508",
X"840583c0",
X"8c08ec05",
X"08820533",
X"8f0683c0",
X"8c08e405",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"e4050883",
X"c08c08e0",
X"05083483",
X"c08c08ec",
X"05088405",
X"3383c08c",
X"08e00508",
X"81053480",
X"0b83c08c",
X"08e00508",
X"82053483",
X"c08c08e0",
X"050808ff",
X"83ff0682",
X"800783c0",
X"8c08e005",
X"080c83c0",
X"8c08e805",
X"08810533",
X"810583c0",
X"8c08e005",
X"0c83c08c",
X"08e00508",
X"83c08c08",
X"e8050881",
X"05348183",
X"3983c08c",
X"08fc0508",
X"802e80f7",
X"3883c08c",
X"08ec0508",
X"86053383",
X"c08c08e0",
X"050c83c0",
X"8c08e005",
X"08a22e09",
X"810680d7",
X"3883c08c",
X"08ec0508",
X"88053383",
X"c08c08ec",
X"05088705",
X"33718280",
X"290583c0",
X"8c08e805",
X"08810533",
X"7080d829",
X"83c08c08",
X"e8050805",
X"83c08c08",
X"e0050c52",
X"83c08c08",
X"e4050c83",
X"c08c08f4",
X"050c83c0",
X"8c08e405",
X"0883c08c",
X"08e00508",
X"88052383",
X"c08c08ec",
X"05083383",
X"c08c08f0",
X"05087131",
X"7083ffff",
X"0683c08c",
X"08f0050c",
X"83c08c08",
X"e0050c83",
X"c08c08ec",
X"05080583",
X"c08c08ec",
X"050cf6d0",
X"3983c08c",
X"08f80508",
X"0d83c08c",
X"08f00508",
X"83c08c08",
X"e0050c83",
X"c08c08f8",
X"05080d83",
X"c08c08e0",
X"050883c0",
X"800c8d3d",
X"0d83c08c",
X"0c0483c0",
X"8c080283",
X"c08c0ce6",
X"3d0d83c0",
X"8c088805",
X"08028405",
X"83c08c08",
X"e8050c83",
X"c08c08d4",
X"050c800b",
X"83cb8434",
X"83c08c08",
X"d4050890",
X"0583c08c",
X"08c0050c",
X"800b83c0",
X"8c08c005",
X"0834800b",
X"83c08c08",
X"c0050881",
X"0534800b",
X"83c08c08",
X"c4050c83",
X"c08c08c4",
X"050880d8",
X"2983c08c",
X"08c00508",
X"0583c08c",
X"08ffb405",
X"0c800b83",
X"c08c08ff",
X"b4050880",
X"d8050c83",
X"c08c08ff",
X"b4050884",
X"0583c08c",
X"08ffb405",
X"0c83c08c",
X"08c40508",
X"83c08c08",
X"ffb40508",
X"34880b83",
X"c08c08ff",
X"b4050881",
X"0534800b",
X"83c08c08",
X"ffb40508",
X"82053483",
X"c08c08ff",
X"b4050808",
X"ffa1ff06",
X"a0800783",
X"c08c08ff",
X"b405080c",
X"83c08c08",
X"c4050881",
X"057081ff",
X"0683c08c",
X"08c4050c",
X"83c08c08",
X"ffb4050c",
X"810b83c0",
X"8c08c405",
X"0827fedb",
X"3883c08c",
X"08ec0570",
X"5483c08c",
X"08c8050c",
X"925283c0",
X"8c08d405",
X"085180cd",
X"993f83c0",
X"800881ff",
X"067083c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb8",
X"05088dea",
X"3883c08c",
X"08f40551",
X"f18c3f83",
X"c0800883",
X"ffff0683",
X"c08c08f6",
X"055283c0",
X"8c08e405",
X"0cf0f33f",
X"83c08008",
X"83ffff06",
X"83c08c08",
X"fd053383",
X"c08c08ff",
X"b8050883",
X"c08c08c4",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08e005",
X"0c83c08c",
X"08c40508",
X"83c08c08",
X"ffbc0508",
X"2780fe38",
X"83c08c08",
X"c8050854",
X"83c08c08",
X"c4050853",
X"895283c0",
X"8c08d405",
X"085180cc",
X"9e3f83c0",
X"800881ff",
X"0683c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"0880f238",
X"83c08c08",
X"ee0551ef",
X"f13f83c0",
X"800883ff",
X"ff065383",
X"c08c08c4",
X"05085283",
X"c08c08d4",
X"050851f0",
X"b33f83c0",
X"8c08c405",
X"08810570",
X"81ff0683",
X"c08c08c4",
X"050c83c0",
X"8c08ffb4",
X"050cfef1",
X"3983c08c",
X"08c00508",
X"81053383",
X"c08c08ff",
X"b4050c81",
X"db0b83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb4",
X"0508802e",
X"8be03894",
X"3983c08c",
X"08ffb805",
X"0883c08c",
X"08ffbc05",
X"0c8bcb39",
X"83c08c08",
X"f1053352",
X"83c08c08",
X"d4050851",
X"80cb9c3f",
X"800b83c0",
X"8c08c005",
X"08810533",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"c4050c83",
X"c08c08c4",
X"050883c0",
X"8c08ffb4",
X"05082789",
X"e63883c0",
X"8c08c405",
X"0880d829",
X"7083c08c",
X"08c00508",
X"05708805",
X"70830533",
X"83c08c08",
X"cc050c83",
X"c08c08c8",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08d805",
X"0c83c08c",
X"08cc0508",
X"87a63883",
X"c08c08c8",
X"05082202",
X"84057186",
X"0587fffc",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08dc050c",
X"83c08c08",
X"ffb8050c",
X"0283c08c",
X"08ffb405",
X"08310d89",
X"3d705983",
X"c08c08ff",
X"b8050858",
X"83c08c08",
X"ffbc0508",
X"87053357",
X"83c08c08",
X"ffb4050c",
X"a25583c0",
X"8c08cc05",
X"08548653",
X"81815283",
X"c08c08d4",
X"050851be",
X"933f83c0",
X"800881ff",
X"0683c08c",
X"08d0050c",
X"83c08c08",
X"d0050881",
X"c13883c0",
X"8c08ffbc",
X"05089605",
X"5383c08c",
X"08ffb805",
X"085283c0",
X"8c08ffb4",
X"050851a1",
X"c63f83c0",
X"800881ff",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb405",
X"08802e81",
X"853883c0",
X"8c08ffbc",
X"05089405",
X"83c08c08",
X"ffbc0508",
X"96053370",
X"862a83c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08cc05",
X"0c83c08c",
X"08ffb405",
X"08832e09",
X"810680c6",
X"3883c08c",
X"08ffb405",
X"0883c08c",
X"08c80508",
X"82053483",
X"cae83370",
X"810583c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb4",
X"050883ca",
X"e83483c0",
X"8c08ffb8",
X"050883c0",
X"8c08cc05",
X"083483c0",
X"8c08dc05",
X"080d83c0",
X"8c08d005",
X"0881ff06",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb80508",
X"fbff3883",
X"c08c08d8",
X"050883c0",
X"8c08c005",
X"08058805",
X"70820533",
X"5183c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb405",
X"08832e09",
X"810680e3",
X"3883c08c",
X"08ffb805",
X"0883c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb405",
X"08810570",
X"81ff0651",
X"83c08c08",
X"ffb4050c",
X"810b83c0",
X"8c08ffb4",
X"050827dd",
X"38800b83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b4050881",
X"057081ff",
X"065183c0",
X"8c08ffb4",
X"050c970b",
X"83c08c08",
X"ffb40508",
X"27dd3883",
X"c08c08e4",
X"050880f9",
X"32703070",
X"80255151",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"e0050891",
X"2e098106",
X"80f93883",
X"c08c08ff",
X"b4050880",
X"2e80ec38",
X"83c08c08",
X"c4050880",
X"e238850b",
X"83c08c08",
X"c00508a6",
X"0534a00b",
X"83c08c08",
X"c00508a7",
X"0534850b",
X"83c08c08",
X"c00508a8",
X"053480c0",
X"0b83c08c",
X"08c00508",
X"a9053486",
X"0b83c08c",
X"08c00508",
X"aa053490",
X"0b83c08c",
X"08c00508",
X"ab053486",
X"0b83c08c",
X"08c00508",
X"ac0534a0",
X"0b83c08c",
X"08c00508",
X"ad053483",
X"c08c08e4",
X"050889d8",
X"32703070",
X"80255151",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"e0050883",
X"edec2e09",
X"810680f6",
X"38817083",
X"c08c08ff",
X"b4050806",
X"83c08c08",
X"ffb4050c",
X"83c08c08",
X"ffb8050c",
X"83c08c08",
X"ffb40508",
X"802e80ce",
X"3883c08c",
X"08c40508",
X"80c43884",
X"0b83c08c",
X"08c00508",
X"aa053480",
X"c00b83c0",
X"8c08c005",
X"08ab0534",
X"840b83c0",
X"8c08c005",
X"08ac0534",
X"900b83c0",
X"8c08c005",
X"08ad0534",
X"83c08c08",
X"ffb80508",
X"83c08c08",
X"c005088c",
X"053483c0",
X"8c08e405",
X"0880f932",
X"70307080",
X"25515183",
X"c08c08ff",
X"b4050c83",
X"c08c08e0",
X"0508862e",
X"09810680",
X"c3388170",
X"83c08c08",
X"ffb40508",
X"0683c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb405",
X"08802e9c",
X"3883c08c",
X"08c40508",
X"933883c0",
X"8c08ffb8",
X"050883c0",
X"8c08c005",
X"088d0534",
X"83c08c08",
X"c4050880",
X"d82983c0",
X"8c08c005",
X"08057084",
X"05708305",
X"3383c08c",
X"08ffb405",
X"0c83c08c",
X"08c8050c",
X"83c08c08",
X"ffbc050c",
X"80588057",
X"83c08c08",
X"ffb40508",
X"56805580",
X"548a53a1",
X"5283c08c",
X"08d40508",
X"51b78d3f",
X"83c08008",
X"81ff0670",
X"30709f2a",
X"5183c08c",
X"08ffb405",
X"0c83c08c",
X"08ffb805",
X"0c83c08c",
X"08ffb805",
X"08a02e8c",
X"3883c08c",
X"08ffb405",
X"08f6c238",
X"83c08c08",
X"ffbc0508",
X"8b053383",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"b4050880",
X"2eb33883",
X"c08c08c8",
X"05088305",
X"3383c08c",
X"08ffb405",
X"0c805880",
X"5783c08c",
X"08ffb405",
X"08568055",
X"80548b53",
X"a15283c0",
X"8c08d405",
X"0851b688",
X"3f83c08c",
X"08c40508",
X"81057081",
X"ff0683c0",
X"8c08c005",
X"08810533",
X"5283c08c",
X"08c4050c",
X"83c08c08",
X"ffb4050c",
X"f6893980",
X"0b83c08c",
X"08c4050c",
X"83c08c08",
X"c4050880",
X"d82983c0",
X"8c08d405",
X"0805709a",
X"053383c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffb8",
X"050c83c0",
X"8c08ffb4",
X"0508822e",
X"098106a9",
X"3883cb84",
X"56815580",
X"5483c08c",
X"08ffb405",
X"085383c0",
X"8c08ffb8",
X"05089705",
X"335283c0",
X"8c08d405",
X"0851e48a",
X"3f83c08c",
X"08c40508",
X"81057081",
X"ff0683c0",
X"8c08c405",
X"0c83c08c",
X"08ffb405",
X"0c810b83",
X"c08c08c4",
X"050827fe",
X"fb38810b",
X"83c08c08",
X"c0050834",
X"800b83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08e805",
X"080d83c0",
X"8c08ffbc",
X"050883c0",
X"800c9c3d",
X"0d83c08c",
X"0c04f53d",
X"0d901e57",
X"800b8118",
X"33545978",
X"7327819d",
X"387880d8",
X"29178a11",
X"33545472",
X"832e0981",
X"0680f838",
X"9414335b",
X"a98c3f83",
X"c080085a",
X"80567581",
X"c4291a87",
X"11335454",
X"72802e80",
X"c0387308",
X"81d4e82e",
X"098106b5",
X"38807459",
X"557480d8",
X"29189a11",
X"33545472",
X"832e0981",
X"069238a4",
X"14703354",
X"547a7327",
X"8738ff13",
X"53727434",
X"81157081",
X"ff065653",
X"817527d1",
X"38811670",
X"81ff0657",
X"538f7627",
X"ffa43883",
X"cae833ff",
X"05537283",
X"cae83481",
X"197081ff",
X"06811933",
X"5e5a537b",
X"7926fee5",
X"38800b83",
X"c0800c8d",
X"3d0d0483",
X"c08c0802",
X"83c08c0c",
X"e63d0d83",
X"c08c0888",
X"05080284",
X"05719005",
X"70337083",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08c8",
X"050c83c0",
X"8c08dc05",
X"0c83c08c",
X"08e0050c",
X"83c08c08",
X"ffa40508",
X"802e94b5",
X"38800b83",
X"c08c08c8",
X"05088105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08d4050c",
X"83c08c08",
X"d4050883",
X"c08c08ff",
X"a4050825",
X"93fd3883",
X"c08c08d4",
X"050880d8",
X"2983c08c",
X"08c80508",
X"05840570",
X"86053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b8050c83",
X"c08c08ff",
X"a4050880",
X"2e938938",
X"a6b23f83",
X"c08c08ff",
X"b8050880",
X"d4050883",
X"c0800826",
X"92f23802",
X"83c08c08",
X"ffb80508",
X"81053383",
X"c08c08ff",
X"a4050c83",
X"c08c08d8",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08fc05",
X"2383c08c",
X"08ffa405",
X"08860583",
X"fc0683c0",
X"8c08ffa4",
X"050c0283",
X"c08c08ff",
X"a4050831",
X"0d853d70",
X"5583c08c",
X"08fc0554",
X"83c08c08",
X"ffb80508",
X"5383c08c",
X"08e00508",
X"5283c08c",
X"08c0050c",
X"ae8a3f83",
X"c0800881",
X"ff0683c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"050891bb",
X"3883c08c",
X"08ffb805",
X"08870533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"802e80d5",
X"3883c08c",
X"08ffb805",
X"08860533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"822e0981",
X"06b33883",
X"c08c08fc",
X"052283c0",
X"8c08ffa4",
X"050c870b",
X"83c08c08",
X"ffa40508",
X"27973883",
X"c08c08c0",
X"05088205",
X"5283c08c",
X"08c00508",
X"3351dba6",
X"3f83c08c",
X"08ffb805",
X"08860533",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"832e0981",
X"0690a438",
X"83c08c08",
X"ffb80508",
X"92057082",
X"053383c0",
X"8c08fc05",
X"2283c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08c4050c",
X"83c08c08",
X"ffa40508",
X"83c08c08",
X"ffa80508",
X"268fe438",
X"800b83c0",
X"8c08e405",
X"0c800b83",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"b0050810",
X"83c08c08",
X"05f80583",
X"c08c08ff",
X"b0050884",
X"2983c08c",
X"08ffb005",
X"08100583",
X"c08c08c4",
X"05080570",
X"84057033",
X"83c08c08",
X"c0050805",
X"703383c0",
X"8c08ffb4",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffbc",
X"05082383",
X"c08c08ff",
X"a8050881",
X"053383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508902e",
X"098106be",
X"3883c08c",
X"08ffa805",
X"083383c0",
X"8c08c005",
X"08058105",
X"70337082",
X"802983c0",
X"8c08ffb4",
X"05080551",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffbc05",
X"082383c0",
X"8c08ffac",
X"05088605",
X"2283c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa805",
X"08a23883",
X"c08c08ff",
X"ac050888",
X"052283c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"050881ff",
X"2e80e538",
X"83c08c08",
X"ffbc0508",
X"227083c0",
X"8c08ffa8",
X"05083170",
X"82802971",
X"3183c08c",
X"08ffac05",
X"08880522",
X"7083c08c",
X"08ffa805",
X"08317073",
X"355383c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffac",
X"050c5183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050883",
X"c08c08ff",
X"bc050823",
X"83c08c08",
X"ffb00508",
X"81057081",
X"ff0683c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa4",
X"050c810b",
X"83c08c08",
X"ffb00508",
X"27fce038",
X"83c08c08",
X"f8052283",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a40508bf",
X"26913883",
X"c08c08e4",
X"05088207",
X"83c08c08",
X"e4050c81",
X"c00b83c0",
X"8c08ffa4",
X"05082791",
X"3883c08c",
X"08e40508",
X"810783c0",
X"8c08e405",
X"0c83c08c",
X"08fa0522",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffa40508",
X"bf269138",
X"83c08c08",
X"e4050888",
X"0783c08c",
X"08e4050c",
X"81c00b83",
X"c08c08ff",
X"a4050827",
X"913883c0",
X"8c08e405",
X"08840783",
X"c08c08e4",
X"050c800b",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffb00508",
X"1083c08c",
X"08c40508",
X"05709005",
X"703383c0",
X"8c08c005",
X"08057033",
X"72810533",
X"70720651",
X"535183c0",
X"8c08ffa8",
X"050c5183",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e9b3890",
X"0b83c08c",
X"08ffb005",
X"082b83c0",
X"8c08e405",
X"080783c0",
X"8c08e405",
X"0c83c08c",
X"08ffb005",
X"08810570",
X"81ff0683",
X"c08c08ff",
X"b0050c83",
X"c08c08ff",
X"a4050c97",
X"0b83c08c",
X"08ffb005",
X"0827fef4",
X"3883c08c",
X"08ffb805",
X"08900533",
X"83c08c08",
X"e4050883",
X"c08c08ff",
X"b4050c83",
X"c08c08c4",
X"050c83c0",
X"8c08ffb4",
X"050883c0",
X"8c08ffb8",
X"05088c05",
X"082e83ff",
X"3883c08c",
X"08ffb405",
X"0883c08c",
X"08ffb805",
X"088c050c",
X"83c08c08",
X"ffb80508",
X"89053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e83b938",
X"83c08c08",
X"e40583c0",
X"8c08ffb4",
X"05088f06",
X"83c08c08",
X"e4050c83",
X"c08c08cc",
X"050c800b",
X"83c08c08",
X"f0050c80",
X"0b83c08c",
X"08f40523",
X"800b81d6",
X"e43383c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffbc",
X"050c83c0",
X"8c08ffa4",
X"050883c0",
X"8c08ffbc",
X"05082e82",
X"d33883c0",
X"8c08f005",
X"81d6e40b",
X"83c08c08",
X"ffac050c",
X"83c08c08",
X"d0050c83",
X"c08c08ff",
X"ac050833",
X"83c08c08",
X"ffac0508",
X"81053381",
X"722b8172",
X"2b077083",
X"c08c08ff",
X"b4050806",
X"5283c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb005",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffa805",
X"082e0981",
X"0681be38",
X"83c08c08",
X"ffbc0508",
X"852680f6",
X"3883c08c",
X"08ffac05",
X"08820533",
X"7081ff06",
X"83c08c08",
X"ffa4050c",
X"83c08c08",
X"ffb0050c",
X"83c08c08",
X"ffa40508",
X"802e80ca",
X"3883c08c",
X"08ffbc05",
X"0883c08c",
X"08ffbc05",
X"08810570",
X"81ff0683",
X"c08c08d0",
X"05087305",
X"5383c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb005",
X"0883c08c",
X"08ffa405",
X"083483c0",
X"8c08ffac",
X"05088305",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e9d",
X"38810b83",
X"c08c08ff",
X"a405082b",
X"83c08c08",
X"cc050808",
X"0783c08c",
X"08cc0508",
X"0c83c08c",
X"08ffac05",
X"08840570",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa405",
X"08fdc838",
X"83c08c08",
X"f0055280",
X"51d0c33f",
X"83c08c08",
X"e4050852",
X"83c08c08",
X"c4050851",
X"d1fe3f83",
X"c08c08fb",
X"05337081",
X"800a2981",
X"0a057098",
X"2c5583c0",
X"8c08ffa4",
X"050c83c0",
X"8c08f905",
X"33708180",
X"0a29810a",
X"0570982c",
X"5583c08c",
X"08ffa405",
X"0c83c08c",
X"08c40508",
X"5383c08c",
X"08ffac05",
X"0c83c08c",
X"08ffa805",
X"0cd1d43f",
X"83c08c08",
X"ffb80508",
X"88053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050880",
X"2e84e038",
X"83c08c08",
X"ffb80508",
X"90053383",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a4050881",
X"2684c038",
X"807081d7",
X"980b81d7",
X"980b8105",
X"3383c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa805",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffb405",
X"0c83c08c",
X"08ffa405",
X"0883c08c",
X"08ffb405",
X"082e81ae",
X"3883c08c",
X"08ffac05",
X"08842983",
X"c08c08ff",
X"a8050805",
X"703383c0",
X"8c08c005",
X"08057033",
X"72810533",
X"70720651",
X"535183c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa4",
X"0508802e",
X"aa38810b",
X"83c08c08",
X"ffac0508",
X"2b83c08c",
X"08ffb405",
X"08077083",
X"ffff0683",
X"c08c08ff",
X"b4050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"ac050881",
X"057081ff",
X"0681d798",
X"71842971",
X"05708105",
X"33515383",
X"c08c08ff",
X"a8050c83",
X"c08c08ff",
X"ac050c83",
X"c08c08ff",
X"a4050c83",
X"c08c08ff",
X"a40508fe",
X"d43883c0",
X"8c08ffb8",
X"05088a05",
X"2283c08c",
X"08c0050c",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"c005082e",
X"82ad3880",
X"0b83c08c",
X"08e8050c",
X"800b83c0",
X"8c08ec05",
X"23807083",
X"c08c08e8",
X"0583c08c",
X"08ffbc05",
X"0c83c08c",
X"08ffac05",
X"0c83c08c",
X"08ffb005",
X"0c81af39",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffac0508",
X"2c708106",
X"5183c08c",
X"08ffa405",
X"0c83c08c",
X"08ffa405",
X"08802e80",
X"e73883c0",
X"8c08ffb0",
X"050883c0",
X"8c08ffb0",
X"05088105",
X"7081ff06",
X"83c08c08",
X"ffbc0508",
X"730583c0",
X"8c08ffb8",
X"05089005",
X"3383c08c",
X"08ffac05",
X"08842905",
X"535383c0",
X"8c08ffb0",
X"050c83c0",
X"8c08ffa8",
X"050c83c0",
X"8c08ffa4",
X"050c83c0",
X"8c08ffa8",
X"050881d7",
X"9a053383",
X"c08c08ff",
X"a4050834",
X"83c08c08",
X"ffac0508",
X"81057081",
X"ff0683c0",
X"8c08ffac",
X"050c83c0",
X"8c08ffa4",
X"050c8f0b",
X"83c08c08",
X"ffac0508",
X"2783c08c",
X"08ffa405",
X"0c83c08c",
X"08ffb005",
X"0885268c",
X"3883c08c",
X"08ffa405",
X"08fea938",
X"83c08c08",
X"e8055280",
X"51caf33f",
X"83c08c08",
X"ffb40508",
X"83c08c08",
X"ffb80508",
X"8a052383",
X"c08c08ff",
X"b8050880",
X"d2053383",
X"c08c08ff",
X"b8050880",
X"d4050805",
X"83c08c08",
X"ffb80508",
X"80d4050c",
X"83c08c08",
X"d805080d",
X"83c08c08",
X"d4050881",
X"800a2981",
X"800a0570",
X"982c83c0",
X"8c08c805",
X"08810533",
X"83c08c08",
X"ffa8050c",
X"5183c08c",
X"08d4050c",
X"83c08c08",
X"ffa80508",
X"83c08c08",
X"d4050824",
X"ec853880",
X"0b83c08c",
X"08ffa805",
X"0c83c08c",
X"08dc0508",
X"0d83c08c",
X"08ffa805",
X"0883c080",
X"0c9c3d0d",
X"83c08c0c",
X"04f33d0d",
X"02bf0533",
X"02840580",
X"c3053383",
X"cb84335a",
X"5b597980",
X"2e8d3878",
X"78065776",
X"802e8e38",
X"81893978",
X"78065776",
X"802e80ff",
X"3883cb84",
X"33707a07",
X"58587988",
X"38780970",
X"79065157",
X"7683cb84",
X"3492973f",
X"83c08008",
X"5e805c8f",
X"5d7d1c87",
X"11335858",
X"76802e80",
X"c1387708",
X"81d4e82e",
X"098106b6",
X"38805b81",
X"5a7d1c70",
X"1c9a1133",
X"59595976",
X"822e0981",
X"06943883",
X"cb845681",
X"55805476",
X"53971833",
X"527851cb",
X"c53fff1a",
X"80d81c5c",
X"5a798025",
X"d038ff1d",
X"81c41d5d",
X"5d7c8025",
X"ffa7388f",
X"3d0d04e9",
X"3d0d696c",
X"02880580",
X"ea05225c",
X"5a5b8070",
X"71415e58",
X"ff78797a",
X"7b7c7d46",
X"4c4a4540",
X"5d436299",
X"3d346202",
X"840580dd",
X"05347779",
X"2280ffff",
X"06544572",
X"79237978",
X"2e888738",
X"7a708105",
X"5c337084",
X"2a718c06",
X"70822a5a",
X"56568306",
X"ff1b7083",
X"ffff065c",
X"54568054",
X"75742e91",
X"387a7081",
X"055c33ff",
X"1b7083ff",
X"ff065c54",
X"54817627",
X"9b387381",
X"ff067b70",
X"81055d33",
X"55748280",
X"2905ff1b",
X"7083ffff",
X"065c5454",
X"827627aa",
X"387383ff",
X"ff067b70",
X"81055d33",
X"70902b72",
X"077d7081",
X"055f3370",
X"982b7207",
X"fe1f7083",
X"ffff0640",
X"52525252",
X"54547e80",
X"2e80c438",
X"7686f738",
X"748a2e09",
X"81069438",
X"811f7081",
X"ff06811e",
X"7081ff06",
X"5f524053",
X"86dc3974",
X"8c2e0981",
X"0686d338",
X"ff1f7081",
X"ff06ff1e",
X"7081ff06",
X"5f524053",
X"7b632586",
X"bd38ff43",
X"86b83976",
X"812e83bb",
X"38768124",
X"89387680",
X"2e8d3886",
X"a5397682",
X"2e84a638",
X"869c39f8",
X"15537284",
X"26849538",
X"72842981",
X"d7d80553",
X"72080464",
X"802e80cd",
X"38782283",
X"80800653",
X"72838080",
X"2e098106",
X"bc388056",
X"756427a4",
X"38751e70",
X"83ffff06",
X"77101b90",
X"1172832a",
X"58515751",
X"53737534",
X"72870681",
X"712b5153",
X"72811634",
X"81167081",
X"ff065753",
X"977627cc",
X"387f8407",
X"40800b99",
X"3d435661",
X"16703370",
X"982b7098",
X"2c515151",
X"53807324",
X"80fb3860",
X"73291e70",
X"83ffff06",
X"7a228380",
X"80065258",
X"53728380",
X"802e0981",
X"0680de38",
X"60883270",
X"30707207",
X"80256390",
X"32703070",
X"72078025",
X"73075354",
X"58515553",
X"73802ebd",
X"38768706",
X"5372b638",
X"75842976",
X"10057911",
X"84117983",
X"2a575751",
X"53737534",
X"60811634",
X"65861423",
X"66881423",
X"7587387f",
X"8107408d",
X"3975812e",
X"09810685",
X"387f8207",
X"40811670",
X"81ff0657",
X"53817627",
X"fee53863",
X"61291e70",
X"83ffff06",
X"5f538070",
X"4642ff02",
X"840580dd",
X"0534ff0b",
X"993d3483",
X"f539811c",
X"7081ff06",
X"5d538042",
X"73812e09",
X"81068e38",
X"7781800a",
X"2981800a",
X"055880d3",
X"3973802e",
X"89387382",
X"2e098106",
X"8d387c81",
X"800a2981",
X"800a055d",
X"a439815f",
X"83b839ff",
X"1c7081ff",
X"065d537b",
X"63258338",
X"ff437c80",
X"2e92387c",
X"81800a29",
X"81ff0a05",
X"5d7c982c",
X"5d839339",
X"77802e92",
X"38778180",
X"0a2981ff",
X"0a055877",
X"982c5882",
X"fd397753",
X"839e3974",
X"892680f4",
X"38748429",
X"81d7ec05",
X"53720804",
X"73872e82",
X"e1387385",
X"2e82db38",
X"73882e82",
X"d538738c",
X"2e82cf38",
X"73892e09",
X"81068638",
X"814582c2",
X"3973812e",
X"09810682",
X"b9386280",
X"2582b338",
X"7b982b70",
X"982c5143",
X"82a83973",
X"83ffff06",
X"46829f39",
X"7383ffff",
X"06478296",
X"397381ff",
X"0641828e",
X"3973811a",
X"34828739",
X"7381ff06",
X"4481ff39",
X"7e5382a0",
X"3974812e",
X"81e33874",
X"81248938",
X"74802e8d",
X"3881e739",
X"74822e81",
X"d83881de",
X"3974567b",
X"83388156",
X"74537386",
X"2e098106",
X"97387581",
X"06537280",
X"2e8e3878",
X"2282ffff",
X"06fe8080",
X"0753b639",
X"7b833881",
X"5373822e",
X"09810697",
X"38728106",
X"5372802e",
X"8e387822",
X"81ffff06",
X"81808007",
X"5393397b",
X"9638fc14",
X"53728126",
X"8e387822",
X"ff808007",
X"53727923",
X"80e53980",
X"5573812e",
X"09810683",
X"38735577",
X"5377802e",
X"89387481",
X"06537280",
X"ca3872d0",
X"15545572",
X"81268338",
X"81557780",
X"2eb93874",
X"81065372",
X"802eb038",
X"78228380",
X"80065372",
X"8380802e",
X"0981069f",
X"3873b02e",
X"09810687",
X"3861993d",
X"34913973",
X"b12e0981",
X"06893861",
X"02840580",
X"dd053461",
X"8105538c",
X"39617431",
X"81055384",
X"39611453",
X"7283ffff",
X"064279f7",
X"fb387d83",
X"2a537282",
X"1a347822",
X"83808006",
X"53728380",
X"802e0981",
X"06883881",
X"537f872e",
X"83388053",
X"7283c080",
X"0c993d0d",
X"04fd3d0d",
X"75831133",
X"82123371",
X"982b7190",
X"2b078114",
X"3370882b",
X"72077533",
X"710783c0",
X"800c5253",
X"54565452",
X"853d0d04",
X"f63d0d02",
X"b7053302",
X"8405bb05",
X"33028805",
X"bf05335b",
X"5b5b8058",
X"80577888",
X"2b7a0756",
X"80557a54",
X"8153a352",
X"7c5192cc",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8c3d0d04",
X"f63d0d02",
X"b7053302",
X"8405bb05",
X"33028805",
X"bf05335b",
X"5b5b8058",
X"80577888",
X"2b7a0756",
X"80557a54",
X"8353a352",
X"7c519290",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8c3d0d04",
X"f73d0d02",
X"b3053302",
X"8405b605",
X"22605a58",
X"56805580",
X"54805381",
X"a3527b51",
X"91e23f83",
X"c0800881",
X"ff0683c0",
X"800c8b3d",
X"0d04ee3d",
X"0d649011",
X"5c5c807b",
X"34800b84",
X"1c0c800b",
X"881c3481",
X"0b891c34",
X"880b8a1c",
X"34800b8b",
X"1c34881b",
X"08c10681",
X"07881c0c",
X"8f3d7054",
X"5d88527b",
X"519beb3f",
X"83c08008",
X"81ff0670",
X"5b597881",
X"a938903d",
X"335e81db",
X"5a7d892e",
X"09810681",
X"99387c53",
X"92527b51",
X"9bc43f83",
X"c0800881",
X"ff06705b",
X"59788182",
X"387c5888",
X"577856a9",
X"55785486",
X"5381a052",
X"7b5190d0",
X"3f83c080",
X"0881ff06",
X"705b5978",
X"80e03802",
X"ba05337b",
X"347c5478",
X"537d527b",
X"519bac3f",
X"83c08008",
X"81ff0670",
X"5b597880",
X"c13802bd",
X"0533527b",
X"519bc43f",
X"83c08008",
X"81ff0670",
X"5b5978aa",
X"38817b33",
X"5a5a7979",
X"26993880",
X"54795388",
X"527b51fd",
X"bb3f811a",
X"7081ff06",
X"7c33525b",
X"59e43981",
X"0b881c34",
X"805a7983",
X"c0800c94",
X"3d0d0480",
X"0b83c080",
X"0c04f93d",
X"0d790284",
X"05ab0533",
X"8e3d7054",
X"585858ff",
X"beb03f8a",
X"3d8a0551",
X"ffbea73f",
X"7551fc8d",
X"3f83c080",
X"08848681",
X"2ebe3883",
X"c0800884",
X"86812699",
X"3883c080",
X"08848280",
X"2e80e638",
X"83c08008",
X"8482812e",
X"9f3881b4",
X"3983c080",
X"0880c082",
X"832e80f4",
X"3883c080",
X"0880c086",
X"832e80e8",
X"38819939",
X"83c09c33",
X"55805674",
X"762e0981",
X"06818b38",
X"74547653",
X"91527751",
X"fbd63f74",
X"54765390",
X"527751fb",
X"cb3f7454",
X"76538452",
X"7751fbfc",
X"3f810b83",
X"c09c3481",
X"b15680de",
X"39805476",
X"53915277",
X"51fba93f",
X"80547653",
X"90527751",
X"fb9e3f80",
X"0b83c09c",
X"34765287",
X"18335197",
X"963fb539",
X"80547653",
X"94527751",
X"fb823f80",
X"54765390",
X"527751fa",
X"f73f7551",
X"ffbcdb3f",
X"83c08008",
X"892a8106",
X"53765287",
X"18335190",
X"cd3f800b",
X"83c09c34",
X"80567583",
X"c0800c89",
X"3d0d04f2",
X"3d0d6090",
X"115a5880",
X"0b881a33",
X"71595656",
X"74762e82",
X"a53882ac",
X"3f841908",
X"83c08008",
X"26829538",
X"78335a81",
X"0b8e3d23",
X"903df811",
X"55f40553",
X"99185277",
X"518ae53f",
X"83c08008",
X"81ff0670",
X"57557477",
X"2e098106",
X"81d93886",
X"39745681",
X"d2398156",
X"82578e3d",
X"33770655",
X"74802ebb",
X"38800b8d",
X"3d34903d",
X"f0055484",
X"53755277",
X"51facd3f",
X"83c08008",
X"81ff0655",
X"749d387b",
X"53755277",
X"51fce73f",
X"83c08008",
X"81ff0655",
X"7481b12e",
X"818b3874",
X"ffb33876",
X"1081fc06",
X"81177081",
X"ff065856",
X"57877627",
X"ffa83881",
X"56757a26",
X"80eb3880",
X"0b8d3d34",
X"8c3d7055",
X"57845375",
X"527751f9",
X"f73f83c0",
X"800881ff",
X"06557480",
X"c1387651",
X"ffbad73f",
X"83c08008",
X"82870655",
X"7482812e",
X"098106aa",
X"3802ae05",
X"33810755",
X"74028405",
X"ae05347b",
X"53755277",
X"51fbeb3f",
X"83c08008",
X"81ff0655",
X"7481b12e",
X"903874fe",
X"b8388116",
X"7081ff06",
X"5755ff91",
X"39805675",
X"81ff0656",
X"973f83c0",
X"80088fd0",
X"05841a0c",
X"75577683",
X"c0800c90",
X"3d0d0404",
X"9080a008",
X"83c0800c",
X"04ff3d0d",
X"7387e829",
X"51ff91cc",
X"3f833d0d",
X"040483cb",
X"880b83c0",
X"800c04fd",
X"3d0d7577",
X"5454800b",
X"83cae834",
X"728a3890",
X"90800b84",
X"150c9039",
X"72812e09",
X"81068838",
X"9098800b",
X"84150c84",
X"140883cb",
X"800c800b",
X"88150c80",
X"0b8c150c",
X"83cb8008",
X"53820b87",
X"80143481",
X"51ff9e3f",
X"83cb8008",
X"53800b88",
X"143483cb",
X"80085381",
X"0b878014",
X"3483cb80",
X"0853800b",
X"8c143483",
X"cb800853",
X"800ba414",
X"34917434",
X"800b83c0",
X"a034800b",
X"83c0a434",
X"800b83c0",
X"a8348054",
X"7381c429",
X"83cb8c05",
X"53800b83",
X"14348114",
X"7081ff06",
X"55538f74",
X"27e63885",
X"3d0d04fe",
X"3d0d7476",
X"82113370",
X"bf068171",
X"2bff0556",
X"51515253",
X"90712783",
X"38ff5276",
X"51717123",
X"83cb8008",
X"51871333",
X"90123480",
X"0b83c0a4",
X"34800b83",
X"c0a83488",
X"13338a14",
X"33525271",
X"802eaa38",
X"7081ff06",
X"51845270",
X"83387052",
X"7183c0a4",
X"348a1333",
X"70307080",
X"25842b70",
X"88075151",
X"52537083",
X"c0a83490",
X"397081ff",
X"06517083",
X"38985271",
X"83c0a834",
X"800b83c0",
X"800c843d",
X"0d04f13d",
X"0d616568",
X"028c0580",
X"cb053302",
X"900580ce",
X"05220294",
X"0580d605",
X"22424041",
X"5a4040fd",
X"8b3f83c0",
X"8008a788",
X"055b8070",
X"715b5b52",
X"83943983",
X"cb800851",
X"7d941234",
X"83c0a433",
X"81075580",
X"7054567f",
X"862680ea",
X"387f8429",
X"81d8a005",
X"83cb8008",
X"53517008",
X"04800b84",
X"1334a139",
X"77337030",
X"70802583",
X"71315151",
X"52537084",
X"13348d39",
X"810b8413",
X"34b83983",
X"0b841334",
X"81705456",
X"ad39810b",
X"841334a2",
X"39773370",
X"30708025",
X"83713151",
X"51525370",
X"84133480",
X"78335252",
X"70833881",
X"52717834",
X"81537488",
X"075583c0",
X"a83383cb",
X"80085257",
X"810b81d0",
X"123483cb",
X"80085181",
X"0b819012",
X"347e802e",
X"ae387280",
X"2ea9387e",
X"ff1e5254",
X"7083ffff",
X"06537283",
X"ffff2e97",
X"38737081",
X"05553383",
X"cb800853",
X"517081c0",
X"1334ff13",
X"51de3983",
X"cb8008a8",
X"11335351",
X"76881234",
X"83cb8008",
X"51747134",
X"81ff5291",
X"3983cb80",
X"08a01133",
X"70810651",
X"5253708f",
X"38fafd3f",
X"7a83c080",
X"0826e638",
X"81883981",
X"0ba01434",
X"83cb8008",
X"a8113380",
X"ff067078",
X"07525351",
X"70802e80",
X"ed387186",
X"2a708106",
X"51517080",
X"2e913880",
X"78335253",
X"70833881",
X"53727834",
X"80e03971",
X"842a7081",
X"06515170",
X"802e9b38",
X"81197083",
X"ffff067d",
X"30709f2a",
X"51525a51",
X"787c2e09",
X"8106af38",
X"a4397183",
X"2a708106",
X"51517080",
X"2e933881",
X"1a7081ff",
X"065b5179",
X"832e0981",
X"0690388a",
X"3971a306",
X"5170802e",
X"85387151",
X"9239f9e4",
X"3f7a83c0",
X"800826fc",
X"e2387181",
X"bf065170",
X"83c0800c",
X"913d0d04",
X"f63d0d02",
X"b3053302",
X"8405b705",
X"33028805",
X"ba052259",
X"5959800b",
X"8c3d348c",
X"3dfc0556",
X"80558054",
X"76537752",
X"7851fbf2",
X"3f83c080",
X"0881ff06",
X"83c0800c",
X"8c3d0d04",
X"f33d0d7f",
X"6264028c",
X"0580c205",
X"22722281",
X"1533425f",
X"415e5959",
X"8078237d",
X"53783352",
X"8151ffa0",
X"3f83c080",
X"0881ff06",
X"5675802e",
X"86387554",
X"81ad3983",
X"cb8008a8",
X"1133821b",
X"3370862a",
X"70810673",
X"982b5351",
X"575c5657",
X"79802583",
X"38815673",
X"762e8738",
X"81f05481",
X"8239818c",
X"17337081",
X"ff067922",
X"7d713190",
X"2b70902c",
X"7009709f",
X"2c720670",
X"52525351",
X"53575754",
X"75742483",
X"38755574",
X"84808029",
X"fc808005",
X"70902c51",
X"5574ff2e",
X"943883cb",
X"80088180",
X"11335154",
X"737c7081",
X"055e34db",
X"39772276",
X"05547378",
X"23790970",
X"9f2a7081",
X"06821c33",
X"81bf0671",
X"862b0751",
X"51515473",
X"821a347c",
X"76268a38",
X"7722547a",
X"7426febb",
X"38805473",
X"83c0800c",
X"8f3d0d04",
X"f93d0d7a",
X"57800b89",
X"3d23893d",
X"fc055376",
X"527951f8",
X"da3f83c0",
X"800881ff",
X"06705755",
X"7496387c",
X"547b5388",
X"3d225276",
X"51fde53f",
X"83c08008",
X"81ff0656",
X"7583c080",
X"0c893d0d",
X"04f03d0d",
X"62660288",
X"0580ce05",
X"22415d5e",
X"80028405",
X"80d20522",
X"7f810533",
X"ff115a5d",
X"5a5d81da",
X"5876bf26",
X"80e93878",
X"802e80e1",
X"387a5878",
X"7b278338",
X"7858821e",
X"3370872a",
X"585a7692",
X"3d34923d",
X"fc055677",
X"557b547e",
X"537d3352",
X"8251f8de",
X"3f83c080",
X"0881ff06",
X"5d800b92",
X"3d33585a",
X"76802e83",
X"38815a82",
X"1e3380ff",
X"067a872b",
X"07577682",
X"1f347c91",
X"38787831",
X"7083ffff",
X"06791e5e",
X"5a57ff9b",
X"397c5877",
X"83c0800c",
X"923d0d04",
X"f83d0d7b",
X"028405b2",
X"05225858",
X"800b8a3d",
X"238a3dfc",
X"05537752",
X"7a51f6f7",
X"3f83c080",
X"0881ff06",
X"70575574",
X"96387d54",
X"7653893d",
X"22527751",
X"feaf3f83",
X"c0800881",
X"ff065675",
X"83c0800c",
X"8a3d0d04",
X"ec3d0d66",
X"6e028805",
X"80df0533",
X"028c0580",
X"e3053302",
X"900580e7",
X"05330294",
X"0580eb05",
X"33029805",
X"80ee0522",
X"4143415f",
X"5c405702",
X"80f20522",
X"963d2396",
X"3df00553",
X"84177053",
X"775259f6",
X"863f83c0",
X"800881ff",
X"06587781",
X"e538777a",
X"81800658",
X"40807725",
X"83388140",
X"79943d34",
X"7b028405",
X"80c90534",
X"7c028405",
X"80ca0534",
X"7d028405",
X"80cb0534",
X"7a953d34",
X"7a882a57",
X"76028405",
X"80cd0534",
X"953d2257",
X"76028405",
X"80ce0534",
X"76882a57",
X"76028405",
X"80cf0534",
X"77923d34",
X"963dec11",
X"57578855",
X"f4175492",
X"3d225377",
X"527751f6",
X"953f83c0",
X"800881ff",
X"06587780",
X"ed387e80",
X"2e80cb38",
X"923d2279",
X"0858587f",
X"802e9c38",
X"76818080",
X"07790c7e",
X"54963dfc",
X"05537783",
X"ffff0652",
X"7851f9fc",
X"3f993976",
X"82808007",
X"790c7e54",
X"953d2253",
X"7783ffff",
X"06527851",
X"fc8f3f83",
X"c0800881",
X"ff065877",
X"9d38923d",
X"22538052",
X"7f307080",
X"25847131",
X"535157f9",
X"873f83c0",
X"800881ff",
X"06587783",
X"c0800c96",
X"3d0d04f6",
X"3d0d7c02",
X"8405b705",
X"335b5b80",
X"58805780",
X"56805579",
X"54855380",
X"527a51fd",
X"a33f83c0",
X"800881ff",
X"06597885",
X"3879871c",
X"347883c0",
X"800c8c3d",
X"0d04f93d",
X"0d02a705",
X"33028405",
X"ab053302",
X"8805af05",
X"33585957",
X"800b83cb",
X"8f335454",
X"72742e9f",
X"38811470",
X"81ff0655",
X"53738f26",
X"81b63873",
X"81c42983",
X"cb8c0583",
X"11335153",
X"72e33873",
X"81c42983",
X"cb880555",
X"800b8716",
X"34768816",
X"34758a16",
X"34778916",
X"3480750c",
X"83cb8008",
X"8c160c80",
X"0b841634",
X"880b8516",
X"34800b86",
X"16348415",
X"08ffa1ff",
X"06a08007",
X"84160c81",
X"147081ff",
X"06535374",
X"51febc3f",
X"83c08008",
X"81ff0670",
X"55537280",
X"cd388a39",
X"7308750c",
X"725480c2",
X"397281dd",
X"bc555681",
X"ddbc0880",
X"2eb23875",
X"84291470",
X"08765370",
X"08515454",
X"722d83c0",
X"800881ff",
X"06537280",
X"2ece3881",
X"167081ff",
X"0681ddbc",
X"71842911",
X"53565753",
X"7208d038",
X"80547383",
X"c0800c89",
X"3d0d04f9",
X"3d0d7957",
X"800b8418",
X"0883cb80",
X"0c58f088",
X"3f881708",
X"83c08008",
X"2783ed38",
X"effa3f83",
X"c0800881",
X"0588180c",
X"83cb8008",
X"b8113370",
X"81ff0651",
X"51547381",
X"2ea43873",
X"81248838",
X"73782e8a",
X"38b83973",
X"822e9538",
X"b1397633",
X"81f00654",
X"73902ea6",
X"38917734",
X"a1397358",
X"763381f0",
X"06547390",
X"2e098106",
X"9138efa8",
X"3f83c080",
X"0881c805",
X"8c180ca0",
X"77348056",
X"7581c429",
X"83cb8f11",
X"33555573",
X"802eaa38",
X"83cb8815",
X"70085654",
X"74802e9d",
X"38881508",
X"802e9638",
X"8c140883",
X"cb80082e",
X"09810689",
X"38735188",
X"15085473",
X"2d811670",
X"81ff0657",
X"548f7627",
X"ffba3876",
X"335473b0",
X"2e819938",
X"73b0248f",
X"3873912e",
X"ab3873a0",
X"2e80f538",
X"82a63973",
X"80d02e81",
X"e4387380",
X"d0248b38",
X"7380c02e",
X"81993882",
X"8f397381",
X"802e81fb",
X"38828539",
X"80567581",
X"c42983cb",
X"8c118311",
X"33565955",
X"73802ea8",
X"3883cb88",
X"15700856",
X"5474802e",
X"9b388c14",
X"0883cb80",
X"082e0981",
X"068e3873",
X"51841508",
X"54732d80",
X"0b831934",
X"81167081",
X"ff065754",
X"8f7627ff",
X"b9389277",
X"3481b539",
X"edc23f8c",
X"170883c0",
X"80082781",
X"a738b077",
X"3481a139",
X"83cb8008",
X"54800b8c",
X"153483cb",
X"80085484",
X"0b881534",
X"80c07734",
X"ed963f83",
X"c08008b2",
X"058c180c",
X"80fa39ed",
X"873f8c17",
X"0883c080",
X"082780ec",
X"3883cb80",
X"0854810b",
X"8c153483",
X"cb800854",
X"800b8815",
X"3483cb80",
X"0854880b",
X"a01534ec",
X"db3f83c0",
X"80089405",
X"8c180c80",
X"d07734bc",
X"3983cb80",
X"08a01133",
X"70832a70",
X"81065151",
X"55557380",
X"2ea63888",
X"0ba01634",
X"ecae3f8c",
X"170883c0",
X"80082794",
X"38ff8077",
X"348e3977",
X"53805280",
X"51fa8b3f",
X"ff907734",
X"83cb8008",
X"a0113370",
X"832a7081",
X"06515155",
X"5573802e",
X"8638880b",
X"a0163489",
X"3d0d04f6",
X"3d0d02b3",
X"05330284",
X"05b70533",
X"5b5b800b",
X"83cb8c70",
X"84127274",
X"5d59575b",
X"58568315",
X"33537280",
X"2e80f338",
X"7333537a",
X"732e0981",
X"0680e738",
X"81143353",
X"79732e09",
X"810680da",
X"38805574",
X"81c42983",
X"cb900570",
X"33831b33",
X"58555373",
X"762e0981",
X"068a3881",
X"13335273",
X"51ff9c3f",
X"81157081",
X"ff065653",
X"8f7527d3",
X"38800b83",
X"cb881970",
X"08565455",
X"73752e91",
X"38725184",
X"14085372",
X"2d83c080",
X"0881ff06",
X"55800b83",
X"18347453",
X"a0398116",
X"81c41981",
X"c41781c4",
X"1781c41d",
X"81c41c5c",
X"5d575759",
X"568f7625",
X"fee83880",
X"537283c0",
X"800c8c3d",
X"0d04f83d",
X"0d02ae05",
X"227d5957",
X"80568155",
X"80548653",
X"8180527a",
X"51f5953f",
X"83c08008",
X"81ff0683",
X"c0800c8a",
X"3d0d04f7",
X"3d0d02b2",
X"05220284",
X"05b70533",
X"605a5b57",
X"80568255",
X"79548653",
X"8180527b",
X"51f4e53f",
X"83c08008",
X"81ff0683",
X"c0800c8b",
X"3d0d04f8",
X"3d0d02af",
X"05335980",
X"58805780",
X"56805578",
X"54895380",
X"527a51f4",
X"bb3f83c0",
X"800881ff",
X"0683c080",
X"0c8a3d0d",
X"04000000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002b0a",
X"00002b4b",
X"00002b6d",
X"00002b93",
X"00002b93",
X"00002b93",
X"00002b93",
X"00002c04",
X"00002c55",
X"0000417a",
X"000049be",
X"00004a77",
X"00ff00ff",
X"00ff00ff",
X"001c0032",
X"00210023",
X"0024002b",
X"00340033",
X"0043003b",
X"0042004b",
X"003a0031",
X"0044004d",
X"0015002d",
X"001b002c",
X"003c002a",
X"001d0022",
X"0035001a",
X"0016001e",
X"00260025",
X"002e0036",
X"003d003e",
X"00460045",
X"005a0076",
X"0066000d",
X"0029004e",
X"00550054",
X"005b005d",
X"005d004c",
X"0052000e",
X"00410049",
X"004a0058",
X"00050006",
X"0004000c",
X"0003000b",
X"0083000a",
X"00010009",
X"00780207",
X"107c0800",
X"00771070",
X"106c107d",
X"10711069",
X"107a1074",
X"106b1072",
X"10750800",
X"104a007c",
X"007b0079",
X"105a0069",
X"0072007a",
X"006b0073",
X"0074006c",
X"0075007d",
X"00700071",
X"0061102f",
X"1037000f",
X"00080010",
X"00180020",
X"00280030",
X"00380040",
X"00140012",
X"0011101f",
X"10140059",
X"10111027",
X"0d0d3f00",
X"0c0c4000",
X"0a0a4100",
X"0b0b4100",
X"07074100",
X"0a0b4300",
X"080b4200",
X"04044500",
X"05054400",
X"06060004",
X"08080004",
X"09090004",
X"00000000",
X"04103a3d",
X"04203b3e",
X"04403c3f",
X"05011e21",
X"05021f22",
X"05042023",
X"05081415",
X"05101a17",
X"0520081c",
X"05400409",
X"0580160a",
X"0601070b",
X"06021d19",
X"06041b05",
X"06080611",
X"00000000",
X"00005703",
X"00005a0a",
X"00005816",
X"00005a0a",
X"00005853",
X"000058a4",
X"000058e3",
X"000058ec",
X"00005a0a",
X"00005a0a",
X"00005a0a",
X"00005a0a",
X"000058f5",
X"000058fd",
X"00005904",
X"00005b0a",
X"00005c03",
X"00005d17",
X"0000600d",
X"00006028",
X"00006014",
X"00006028",
X"0000602f",
X"0000603a",
X"00006041",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"66726565",
X"7a65722e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00006c7c",
X"00006c80",
X"00006c88",
X"00006c94",
X"00006ca0",
X"00006cac",
X"00006cb8",
X"00006cbc",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00006c14",
X"00006a68",
X"00000000",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"69383030",
X"00000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
