
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80e9",
X"b4738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80ec",
X"ec0c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580e6",
X"ec2d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580e6ab",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80d08c04",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"775193b0",
X"3f83e080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3380ecf4",
X"0b80ecf4",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"52775192",
X"df3f83e0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583e0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"55b3963f",
X"83e08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"811451b2",
X"ae3f83e0",
X"80083070",
X"83e08008",
X"07802583",
X"e0800c53",
X"863d0d04",
X"fc3d0d76",
X"70525599",
X"cd3f83e0",
X"80085481",
X"5383e080",
X"0880c738",
X"74519990",
X"3f83e080",
X"080b0b80",
X"eaf45383",
X"e0800852",
X"53ff8f3f",
X"83e08008",
X"a5380b0b",
X"80eaf852",
X"7251fefe",
X"3f83e080",
X"0894380b",
X"0b80eafc",
X"527251fe",
X"ed3f83e0",
X"8008802e",
X"83388154",
X"73537283",
X"e0800c86",
X"3d0d04fd",
X"3d0d7570",
X"525498e6",
X"3f815383",
X"e0800898",
X"38735198",
X"af3f83e0",
X"a0085283",
X"e0800851",
X"feb43f83",
X"e0800853",
X"7283e080",
X"0c853d0d",
X"04e03d0d",
X"a33d0870",
X"525e8ed1",
X"3f83e080",
X"0833943d",
X"56547394",
X"3880eff0",
X"52745184",
X"c6397d52",
X"785191d6",
X"3f84d039",
X"7d518eb9",
X"3f83e080",
X"08527451",
X"8de93f83",
X"e0a80852",
X"933d7052",
X"5d94c73f",
X"83e08008",
X"59800b83",
X"e0800855",
X"5b83e080",
X"087b2e94",
X"38811b74",
X"525b97c9",
X"3f83e080",
X"085483e0",
X"8008ee38",
X"805aff7a",
X"437a427a",
X"415f7909",
X"709f2c7b",
X"065b547a",
X"7a248438",
X"ff1b5af6",
X"1a700970",
X"9f2c7206",
X"7bff125a",
X"5a525555",
X"80752595",
X"38765197",
X"883f83e0",
X"800876ff",
X"18585557",
X"738024ed",
X"38747f2e",
X"8638b8a0",
X"3f745f78",
X"ff1b7058",
X"5d58807a",
X"25953877",
X"5196de3f",
X"83e08008",
X"76ff1858",
X"55587380",
X"24ed3880",
X"0b83e3a8",
X"0c800b83",
X"e3c80c0b",
X"0b80eb80",
X"518bad3f",
X"81800b83",
X"e3c80c0b",
X"0b80eb88",
X"518b9d3f",
X"a80b83e3",
X"a80c7680",
X"2e80e838",
X"83e3a808",
X"77793270",
X"30707207",
X"80257087",
X"2b83e3c8",
X"0c515678",
X"53565696",
X"913f83e0",
X"8008802e",
X"8a380b0b",
X"80eb9051",
X"8ae23f76",
X"5195d13f",
X"83e08008",
X"520b0b80",
X"ec9c518a",
X"cf3f7651",
X"95d73f83",
X"e0800883",
X"e3a80855",
X"57757425",
X"8638a816",
X"56f73975",
X"83e3a80c",
X"86f07624",
X"ff943887",
X"980b83e3",
X"a80c7780",
X"2eb73877",
X"51958d3f",
X"83e08008",
X"78525595",
X"ad3f0b0b",
X"80eb9854",
X"83e08008",
X"8f388739",
X"807634fd",
X"96390b0b",
X"80eb9454",
X"74537352",
X"0b0b80ea",
X"e85189e8",
X"3f80540b",
X"0b80ece8",
X"5189dd3f",
X"81145473",
X"a82e0981",
X"06ed3886",
X"8da051b4",
X"a23f8052",
X"903d7052",
X"5480d4f4",
X"3f835273",
X"5180d4ec",
X"3f61802e",
X"80ff387b",
X"5473ff2e",
X"96387880",
X"2e818038",
X"785194ad",
X"3f83e080",
X"08ff1555",
X"59e73978",
X"802e80eb",
X"38785194",
X"a93f83e0",
X"8008802e",
X"fc843878",
X"5193f13f",
X"83e08008",
X"520b0b80",
X"eaf051ab",
X"d13f83e0",
X"8008a438",
X"7c51ad89",
X"3f83e080",
X"085574ff",
X"16565480",
X"7425fbef",
X"38741d70",
X"33555673",
X"af2efec8",
X"38e83978",
X"5193af3f",
X"83e08008",
X"527c51ac",
X"c03ffbcf",
X"397f8829",
X"6010057a",
X"0561055a",
X"fc8039a2",
X"3d0d0480",
X"3d0d9080",
X"f8337081",
X"ff067084",
X"2a813270",
X"81065151",
X"51517080",
X"2e8d38a8",
X"0b9080f8",
X"34b80b90",
X"80f83470",
X"83e0800c",
X"823d0d04",
X"803d0d90",
X"80f83370",
X"81ff0670",
X"852a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"980b9080",
X"f834b80b",
X"9080f834",
X"7083e080",
X"0c823d0d",
X"04930b90",
X"80fc34ff",
X"0b9080e8",
X"3404ff3d",
X"0d028f05",
X"3352800b",
X"9080fc34",
X"8a51b1f7",
X"3fdf3f80",
X"f80b9080",
X"e034800b",
X"9080c834",
X"fa125271",
X"9080c034",
X"800b9080",
X"d8347190",
X"80d03490",
X"80f85280",
X"7234b872",
X"34833d0d",
X"04803d0d",
X"028b0533",
X"51709080",
X"f434febf",
X"3f83e080",
X"08802ef6",
X"38823d0d",
X"04803d0d",
X"8439bbb6",
X"3ffed93f",
X"83e08008",
X"802ef338",
X"9080f433",
X"7081ff06",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"a30b9080",
X"fc34ff0b",
X"9080e834",
X"9080f851",
X"a87134b8",
X"7134823d",
X"0d04803d",
X"0d9080fc",
X"337081c0",
X"06703070",
X"802583e0",
X"800c5151",
X"51823d0d",
X"04803d0d",
X"9080f833",
X"7081ff06",
X"70832a81",
X"32708106",
X"51515151",
X"70802ee8",
X"38b00b90",
X"80f834b8",
X"0b9080f8",
X"34823d0d",
X"04803d0d",
X"9080ac08",
X"810683e0",
X"800c823d",
X"0d04fd3d",
X"0d757754",
X"54807325",
X"94387370",
X"81055533",
X"5280eb9c",
X"5185a13f",
X"ff1353e9",
X"39853d0d",
X"04f63d0d",
X"7c7e6062",
X"5a5d5b56",
X"80598155",
X"8539747a",
X"29557452",
X"755180d1",
X"d63f83e0",
X"80087a27",
X"ed387480",
X"2e80e038",
X"74527551",
X"80d1c03f",
X"83e08008",
X"75537652",
X"5480d1c3",
X"3f83e080",
X"087a5375",
X"525680d1",
X"a63f83e0",
X"80087930",
X"707b079f",
X"2a707780",
X"24075151",
X"54557287",
X"3883e080",
X"08c23876",
X"8118b016",
X"55585889",
X"74258b38",
X"b714537a",
X"853880d7",
X"14537278",
X"34811959",
X"ff9c3980",
X"77348c3d",
X"0d04f73d",
X"0d7b7d7f",
X"62029005",
X"bb053357",
X"59565a5a",
X"b0587283",
X"38a05875",
X"70708105",
X"52337159",
X"54559039",
X"8074258e",
X"38ff1477",
X"70810559",
X"33545472",
X"ef3873ff",
X"15555380",
X"73258938",
X"77527951",
X"782def39",
X"75337557",
X"5372802e",
X"90387252",
X"7951782d",
X"75708105",
X"573353ed",
X"398b3d0d",
X"04ee3d0d",
X"64666969",
X"70708105",
X"52335b4a",
X"5c5e5e76",
X"802e82f9",
X"3876a52e",
X"09810682",
X"e0388070",
X"41677070",
X"81055233",
X"714a5957",
X"5f76b02e",
X"0981068c",
X"38757081",
X"05573376",
X"4857815f",
X"d0175675",
X"892680da",
X"3876675c",
X"59805c93",
X"39778a24",
X"80c3387b",
X"8a29187b",
X"7081055d",
X"335a5cd0",
X"197081ff",
X"06585889",
X"7727a438",
X"ff9f1970",
X"81ff06ff",
X"a91b5a51",
X"56857627",
X"9238ffbf",
X"197081ff",
X"06515675",
X"85268a38",
X"c9195877",
X"8025ffb9",
X"387a477b",
X"407881ff",
X"06577680",
X"e42e80e5",
X"387680e4",
X"24a73876",
X"80d82e81",
X"86387680",
X"d8249038",
X"76802e81",
X"cc3876a5",
X"2e81b638",
X"81b93976",
X"80e32e81",
X"8c3881af",
X"397680f5",
X"2e9b3876",
X"80f5248b",
X"387680f3",
X"2e818138",
X"81993976",
X"80f82e80",
X"ca38818f",
X"39913d70",
X"55578053",
X"8a527984",
X"1b710853",
X"5b56fbfd",
X"3f7655ab",
X"3979841b",
X"7108943d",
X"705b5b52",
X"5b567580",
X"258c3875",
X"3056ad78",
X"340280c1",
X"05577654",
X"80538a52",
X"7551fbd1",
X"3f77557e",
X"54b83991",
X"3d705577",
X"80d83270",
X"30708025",
X"56515856",
X"90527984",
X"1b710853",
X"5b57fbad",
X"3f7555db",
X"3979841b",
X"83123354",
X"5b569839",
X"79841b71",
X"08575b56",
X"80547f53",
X"7c527d51",
X"fc9c3f87",
X"3976527d",
X"517c2d66",
X"70335881",
X"0547fd83",
X"39943d0d",
X"047283e0",
X"900c7183",
X"e0940c04",
X"fb3d0d88",
X"3d707084",
X"05520857",
X"54755383",
X"e0900852",
X"83e09408",
X"51fcc63f",
X"873d0d04",
X"ff3d0d73",
X"70085351",
X"02930533",
X"72347008",
X"8105710c",
X"833d0d04",
X"fc3d0d87",
X"3d881155",
X"785499d0",
X"5351fc99",
X"3f805287",
X"3d51d13f",
X"863d0d04",
X"fd3d0d75",
X"705254a3",
X"c83f83e0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83e0",
X"8008732e",
X"a13883e0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183e0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83e2d408",
X"248b3880",
X"cde63fff",
X"0b83e2d4",
X"0c800b83",
X"e0800c04",
X"ff3d0d73",
X"5283e0b0",
X"08722e8d",
X"38d83f71",
X"51969c3f",
X"7183e0b0",
X"0c833d0d",
X"04f43d0d",
X"7e60625c",
X"5a558154",
X"bc150881",
X"92387451",
X"cf3f7958",
X"807a2580",
X"f83883e3",
X"84087089",
X"2a5783ff",
X"06788480",
X"72315656",
X"57737825",
X"83387355",
X"7583e2d4",
X"082e8438",
X"ff883f83",
X"e2d40880",
X"25a63875",
X"892b5198",
X"df3f83e3",
X"84088f3d",
X"fc11555c",
X"548152f8",
X"1b5196c9",
X"3f761483",
X"e3840c75",
X"83e2d40c",
X"74537652",
X"785180cb",
X"f83f83e0",
X"800883e3",
X"84081683",
X"e3840c78",
X"7631761b",
X"5b595677",
X"8024ff8a",
X"38617a71",
X"0c547554",
X"75802e83",
X"38815473",
X"83e0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"993f7651",
X"feae3f86",
X"3dfc0553",
X"78527751",
X"95eb3f79",
X"75710c54",
X"83e08008",
X"5483e080",
X"08802e83",
X"38815473",
X"83e0800c",
X"863d0d04",
X"fe3d0d75",
X"83e2d408",
X"53538072",
X"24893871",
X"732e8438",
X"fdd43f74",
X"51fde93f",
X"725197b0",
X"3f83e080",
X"085283e0",
X"8008802e",
X"83388152",
X"7183e080",
X"0c843d0d",
X"04803d0d",
X"7280c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d72bc11",
X"0883e080",
X"0c51823d",
X"0d0480c4",
X"0b83e080",
X"0c04fd3d",
X"0d757771",
X"54705355",
X"539f9e3f",
X"82c81308",
X"bc150c82",
X"c0130880",
X"c0150cfc",
X"e93f7351",
X"93ad3f73",
X"83e0b00c",
X"83e08008",
X"5383e080",
X"08802e83",
X"38815372",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"775553fc",
X"bd3f7280",
X"2ea538bc",
X"13085273",
X"519ea83f",
X"83e08008",
X"8f387752",
X"7251ff9a",
X"3f83e080",
X"08538a39",
X"82cc1308",
X"53d83981",
X"537283e0",
X"800c853d",
X"0d04fe3d",
X"0dff0b83",
X"e2d40c74",
X"83e0b40c",
X"7583e2d0",
X"0c80c8bb",
X"3f83e080",
X"0881ff06",
X"52815371",
X"993883e2",
X"ec518e96",
X"3f83e080",
X"085283e0",
X"8008802e",
X"83387252",
X"71537283",
X"e0800c84",
X"3d0d04fa",
X"3d0d787a",
X"82c41208",
X"82c41208",
X"70722459",
X"56565757",
X"73732e09",
X"81069138",
X"80c01652",
X"80c01751",
X"9c983f83",
X"e0800855",
X"7483e080",
X"0c883d0d",
X"04f63d0d",
X"7c5b807b",
X"715c5457",
X"7a772e8c",
X"38811a82",
X"cc140854",
X"5a72f638",
X"805980d9",
X"397a5481",
X"5780707b",
X"7b315a57",
X"55ff1853",
X"74732580",
X"c13882cc",
X"14085273",
X"51ff8c3f",
X"800b83e0",
X"800825a1",
X"3882cc14",
X"0882cc11",
X"0882cc16",
X"0c7482cc",
X"120c5375",
X"802e8638",
X"7282cc17",
X"0c725480",
X"577382cc",
X"15088117",
X"575556ff",
X"b8398119",
X"59800bff",
X"1b545478",
X"73258338",
X"81547681",
X"32707506",
X"515372ff",
X"90388c3d",
X"0d04f73d",
X"0d7b7d5a",
X"5a82d052",
X"83e2d008",
X"5180c4db",
X"3f83e080",
X"0857f9de",
X"3f795283",
X"e2d85195",
X"b63f83e0",
X"80085480",
X"5383e080",
X"08732e09",
X"81068283",
X"3883e0b4",
X"080b0b80",
X"eaf05370",
X"52569bd5",
X"3f0b0b80",
X"eaf05280",
X"c016519b",
X"c83f75bc",
X"170c7382",
X"c0170c81",
X"0b82c417",
X"0c810b82",
X"c8170c73",
X"82cc170c",
X"ff1782d0",
X"17555781",
X"913983e0",
X"c0337082",
X"2a708106",
X"51545572",
X"81803874",
X"812a8106",
X"587780f6",
X"3874842a",
X"810682c4",
X"150c83e0",
X"c0338106",
X"82c8150c",
X"79527351",
X"9aef3f73",
X"519b863f",
X"83e08008",
X"1453af73",
X"70810555",
X"3472bc15",
X"0c83e0c1",
X"5272519a",
X"d03f83e0",
X"b80882c0",
X"150c83e0",
X"ce5280c0",
X"14519abd",
X"3f78802e",
X"8d387351",
X"782d83e0",
X"8008802e",
X"99387782",
X"cc150c75",
X"802e8638",
X"7382cc17",
X"0c7382d0",
X"15ff1959",
X"55567680",
X"2e9b3883",
X"e0b85283",
X"e2d85194",
X"ac3f83e0",
X"80088a38",
X"83e0c133",
X"5372fed2",
X"3878802e",
X"893883e0",
X"b40851fc",
X"b83f83e0",
X"b4085372",
X"83e0800c",
X"8b3d0d04",
X"ff3d0d80",
X"527351fd",
X"b53f833d",
X"0d04f03d",
X"0d627052",
X"54f68d3f",
X"83e08008",
X"7453873d",
X"70535555",
X"f6ad3ff7",
X"8d3f7351",
X"d33f6353",
X"745283e0",
X"800851fa",
X"b73f923d",
X"0d047183",
X"e0800c04",
X"80c01283",
X"e0800c04",
X"803d0d72",
X"82c01108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"7282cc11",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282c4",
X"110883e0",
X"800c5182",
X"3d0d04f9",
X"3d0d7983",
X"e0980857",
X"57817727",
X"81983876",
X"88170827",
X"81903875",
X"33557482",
X"2e893874",
X"832eb438",
X"81803974",
X"54761083",
X"fe065376",
X"882a8c17",
X"08055289",
X"3dfc0551",
X"80c2d53f",
X"83e08008",
X"80e03802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d23984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"5180c2a4",
X"3f83e080",
X"08b03802",
X"9f053302",
X"84059e05",
X"3371982b",
X"71902b07",
X"028c059d",
X"05337088",
X"2b72078d",
X"3d337180",
X"fffffe80",
X"06075152",
X"53575856",
X"83398155",
X"7483e080",
X"0c893d0d",
X"04fb3d0d",
X"83e09808",
X"fe198812",
X"08fe0555",
X"56548056",
X"7473278d",
X"38821433",
X"75712994",
X"16080557",
X"537583e0",
X"800c873d",
X"0d04fc3d",
X"0d765280",
X"0b83e098",
X"08703351",
X"52537083",
X"2e098106",
X"91389512",
X"33941333",
X"71982b71",
X"902b0755",
X"55519b12",
X"339a1333",
X"71882b07",
X"740783e0",
X"800c5586",
X"3d0d04fc",
X"3d0d7683",
X"e0980855",
X"55807523",
X"88150853",
X"72812e88",
X"38881408",
X"73268538",
X"8152b239",
X"72903873",
X"33527183",
X"2e098106",
X"85389014",
X"0853728c",
X"160c7280",
X"2e8d3872",
X"51fed63f",
X"83e08008",
X"52853990",
X"14085271",
X"90160c80",
X"527183e0",
X"800c863d",
X"0d04fa3d",
X"0d7883e0",
X"98087122",
X"81057083",
X"ffff0657",
X"54575573",
X"802e8838",
X"90150853",
X"72863883",
X"5280e739",
X"738f0652",
X"7180da38",
X"81139016",
X"0c8c1508",
X"53729038",
X"830b8417",
X"22575273",
X"762780c6",
X"38bf3982",
X"1633ff05",
X"74842a06",
X"5271b238",
X"7251fcaf",
X"3f815271",
X"83e08008",
X"27a83883",
X"5283e080",
X"08881708",
X"279c3883",
X"e080088c",
X"160c83e0",
X"800851fd",
X"bc3f83e0",
X"80089016",
X"0c737523",
X"80527183",
X"e0800c88",
X"3d0d04f2",
X"3d0d6062",
X"64585e5b",
X"75335574",
X"a02e0981",
X"06883881",
X"16704456",
X"ef396270",
X"33565674",
X"af2e0981",
X"06843881",
X"1643800b",
X"881c0c62",
X"70335155",
X"749f2691",
X"387a51fd",
X"d23f83e0",
X"80085680",
X"7d348381",
X"39933d84",
X"1c087058",
X"595f8a55",
X"a0767081",
X"055834ff",
X"155574ff",
X"2e098106",
X"ef388070",
X"5a5c887f",
X"085f5a7b",
X"811d7081",
X"ff066013",
X"703370af",
X"327030a0",
X"73277180",
X"25075151",
X"525b535e",
X"57557480",
X"e73876ae",
X"2e098106",
X"83388155",
X"787a2775",
X"07557480",
X"2e9f3879",
X"88327030",
X"78ae3270",
X"30707307",
X"9f2a5351",
X"57515675",
X"bb388859",
X"8b5affab",
X"3976982b",
X"55748025",
X"873880e8",
X"c4173357",
X"ff9f1755",
X"74992689",
X"38e01770",
X"81ff0658",
X"5578811a",
X"7081ff06",
X"721b535b",
X"57557675",
X"34fef839",
X"7b1e7f0c",
X"805576a0",
X"26833881",
X"55748b19",
X"347a51fc",
X"823f83e0",
X"800880f5",
X"38a0547a",
X"2270852b",
X"83e00654",
X"55901b08",
X"527c51bc",
X"df3f83e0",
X"80085783",
X"e0800881",
X"81387c33",
X"5574802e",
X"80f4388b",
X"1d337083",
X"2a708106",
X"51565674",
X"b4388b7d",
X"841d0883",
X"e0800859",
X"5b5b58ff",
X"185877ff",
X"2e9a3879",
X"7081055b",
X"33797081",
X"055b3371",
X"71315256",
X"5675802e",
X"e2388639",
X"75802e96",
X"387a51fb",
X"e53fff86",
X"3983e080",
X"085683e0",
X"8008b638",
X"83397656",
X"841b088b",
X"11335155",
X"74a7388b",
X"1d337084",
X"2a708106",
X"51565674",
X"89388356",
X"94398156",
X"90397c51",
X"fa943f83",
X"e0800888",
X"1c0cfd81",
X"397583e0",
X"800c903d",
X"0d04f83d",
X"0d7a7c59",
X"57825483",
X"fe537752",
X"7651bba4",
X"3f835683",
X"e0800880",
X"ec388117",
X"33773371",
X"882b0756",
X"56825674",
X"82d4d52e",
X"09810680",
X"d4387554",
X"b6537752",
X"7651baf8",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"ac388254",
X"80d25377",
X"527651ba",
X"cf3f83e0",
X"80089838",
X"81173377",
X"3371882b",
X"0783e080",
X"08525656",
X"748182c6",
X"2e833881",
X"567583e0",
X"800c8a3d",
X"0d04eb3d",
X"0d675a80",
X"0b83e098",
X"0cba843f",
X"83e08008",
X"81065582",
X"567483ee",
X"38747553",
X"8f3d7053",
X"5759feca",
X"3f83e080",
X"0881ff06",
X"5776812e",
X"09810680",
X"d4389054",
X"83be5374",
X"527551b9",
X"e33f83e0",
X"800880c9",
X"388f3d33",
X"5574802e",
X"80c93802",
X"bf053302",
X"8405be05",
X"3371982b",
X"71902b07",
X"028c05bd",
X"05337088",
X"2b720795",
X"3d337107",
X"70587b57",
X"5e525e57",
X"5957fdee",
X"3f83e080",
X"0881ff06",
X"5776832e",
X"09810686",
X"38815682",
X"f1397680",
X"2e863886",
X"5682e739",
X"a4548d53",
X"78527551",
X"b8fa3f81",
X"5683e080",
X"0882d338",
X"02be0533",
X"028405bd",
X"05337188",
X"2b07595d",
X"77ab3802",
X"80ce0533",
X"02840580",
X"cd053371",
X"982b7190",
X"2b07973d",
X"3370882b",
X"72070294",
X"0580cb05",
X"33710754",
X"525e5759",
X"5602b705",
X"33787129",
X"028805b6",
X"0533028c",
X"05b50533",
X"71882b07",
X"701d707f",
X"8c050c5f",
X"5957595d",
X"8e3d3382",
X"1b3402b9",
X"0533903d",
X"3371882b",
X"075a5c78",
X"841b2302",
X"bb053302",
X"8405ba05",
X"3371882b",
X"07565c74",
X"ab380280",
X"ca053302",
X"840580c9",
X"05337198",
X"2b71902b",
X"07963d33",
X"70882b72",
X"07029405",
X"80c70533",
X"71075152",
X"53575e5c",
X"74763178",
X"3179842a",
X"903d3354",
X"71713153",
X"5656b5bf",
X"3f83e080",
X"08820570",
X"881c0c83",
X"e08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83e0980c",
X"80567583",
X"e0800c97",
X"3d0d04e9",
X"3d0d83e0",
X"98085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e63f83e0",
X"80085483",
X"e0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f48a",
X"3f83e080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383e080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83e09808",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0e83f",
X"83e08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"843f83e0",
X"80085583",
X"e0800880",
X"2eff8938",
X"83e08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"51b3a13f",
X"83e08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83e0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83e09808",
X"55568555",
X"73802e81",
X"e1388114",
X"33810653",
X"84557280",
X"2e81d338",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b7388214",
X"3370892b",
X"56537680",
X"2eb53874",
X"52ff1651",
X"b0c13f83",
X"e08008ff",
X"18765470",
X"535853b0",
X"b23f83e0",
X"80087326",
X"96387430",
X"70780670",
X"98170c77",
X"7131a417",
X"08525851",
X"538939a0",
X"140870a4",
X"160c5374",
X"7627b938",
X"7251eed7",
X"3f83e080",
X"0853810b",
X"83e08008",
X"278b3888",
X"140883e0",
X"80082688",
X"38800b81",
X"1534b039",
X"83e08008",
X"a4150c98",
X"14081598",
X"150c7575",
X"3156c439",
X"98140816",
X"7098160c",
X"735256ef",
X"c83f83e0",
X"80088c38",
X"83e08008",
X"81153481",
X"55943982",
X"1433ff05",
X"76892a06",
X"83e08008",
X"05a8150c",
X"80557483",
X"e0800c88",
X"3d0d04ef",
X"3d0d6356",
X"855583e0",
X"9808802e",
X"80d23893",
X"3df40584",
X"170c6453",
X"883d7053",
X"765257f1",
X"d23f83e0",
X"80085583",
X"e08008b4",
X"38883d33",
X"5473802e",
X"a13802a7",
X"05337084",
X"2a708106",
X"51555583",
X"5573802e",
X"97387651",
X"eef83f83",
X"e0800888",
X"170c7551",
X"efa93f83",
X"e0800855",
X"7483e080",
X"0c933d0d",
X"04e43d0d",
X"6ea13d08",
X"405e8556",
X"83e09808",
X"802e8485",
X"389e3df4",
X"05841f0c",
X"7e98387d",
X"51eef83f",
X"83e08008",
X"5683ee39",
X"814181f6",
X"39834181",
X"f139933d",
X"7f960541",
X"59807f82",
X"95055e56",
X"756081ff",
X"05348341",
X"901e0876",
X"2e81d338",
X"a0547d22",
X"70852b83",
X"e0065458",
X"901e0852",
X"7851afac",
X"3f83e080",
X"084183e0",
X"8008ffb8",
X"3878335c",
X"7b802eff",
X"b4388b19",
X"3370bf06",
X"71810652",
X"43557480",
X"2e80de38",
X"7b81bf06",
X"55748f24",
X"80d3389a",
X"19335574",
X"80cb38f3",
X"1d70585d",
X"8156758b",
X"2e098106",
X"85388e56",
X"8b39759a",
X"2e098106",
X"83389c56",
X"75197070",
X"81055233",
X"7133811a",
X"821a5f5b",
X"525b5574",
X"86387977",
X"34853980",
X"df773477",
X"7b57577a",
X"a02e0981",
X"06c03881",
X"567b81e5",
X"32703070",
X"9f2a5151",
X"557bae2e",
X"93387480",
X"2e8e3861",
X"832a7081",
X"06515574",
X"802e9738",
X"7d51ede2",
X"3f83e080",
X"084183e0",
X"80088738",
X"901e08fe",
X"af388060",
X"3475802e",
X"88387c52",
X"7f5183a5",
X"3f60802e",
X"8638800b",
X"901f0c60",
X"5660832e",
X"85386081",
X"d038891f",
X"57901e08",
X"802e81a8",
X"38805675",
X"19703351",
X"5574a02e",
X"a0387485",
X"2e098106",
X"843881e5",
X"55747770",
X"81055934",
X"81167081",
X"ff065755",
X"877627d7",
X"38881933",
X"5574a02e",
X"a938ae77",
X"70810559",
X"34885675",
X"19703351",
X"5574a02e",
X"95387477",
X"70810559",
X"34811670",
X"81ff0657",
X"558a7627",
X"e2388b19",
X"337f8805",
X"349f1933",
X"9e1a3371",
X"982b7190",
X"2b079d1c",
X"3370882b",
X"72079c1e",
X"33710764",
X"0c52991d",
X"33981e33",
X"71882b07",
X"53515357",
X"5956747f",
X"84052397",
X"1933961a",
X"3371882b",
X"07565674",
X"7f860523",
X"8077347d",
X"51ebf33f",
X"83e08008",
X"83327030",
X"7072079f",
X"2c83e080",
X"08065256",
X"56961f33",
X"55748a38",
X"891f5296",
X"1f5181b1",
X"3f7583e0",
X"800c9e3d",
X"0d04fd3d",
X"0d757753",
X"54733351",
X"70893871",
X"33517080",
X"2ea13873",
X"33723352",
X"53727127",
X"8538ff51",
X"94397073",
X"27853881",
X"518b3981",
X"14811353",
X"54d33980",
X"517083e0",
X"800c853d",
X"0d04fd3d",
X"0d757754",
X"54723370",
X"81ff0652",
X"5270802e",
X"a3387181",
X"ff068114",
X"ffbf1253",
X"54527099",
X"268938a0",
X"127081ff",
X"06535171",
X"74708105",
X"5634d239",
X"80743485",
X"3d0d04ff",
X"bd3d0d80",
X"c63d0852",
X"a53d7052",
X"54ffb33f",
X"80c73d08",
X"52853d70",
X"5253ffa6",
X"3f725273",
X"51fedf3f",
X"80c53d0d",
X"04fe3d0d",
X"74765353",
X"71708105",
X"53335170",
X"73708105",
X"553470f0",
X"38843d0d",
X"04fe3d0d",
X"74528072",
X"33525370",
X"732e8d38",
X"81128114",
X"71335354",
X"5270f538",
X"7283e080",
X"0c843d0d",
X"047183e3",
X"9c0c8880",
X"800b83e3",
X"980c8480",
X"800b83e3",
X"a00c04fd",
X"3d0d7770",
X"17557705",
X"ff1a5353",
X"71ff2e94",
X"38737081",
X"05553351",
X"70737081",
X"055534ff",
X"1252e939",
X"853d0d04",
X"fc3d0d87",
X"a6815574",
X"3383e3a4",
X"34a05483",
X"a0805383",
X"e39c0852",
X"83e39808",
X"51ffb83f",
X"a05483a4",
X"805383e3",
X"9c085283",
X"e3980851",
X"ffa53f90",
X"5483a880",
X"5383e39c",
X"085283e3",
X"980851ff",
X"923fa053",
X"805283e3",
X"a00883a0",
X"80055185",
X"8b3fa053",
X"805283e3",
X"a00883a4",
X"80055184",
X"fb3f9053",
X"805283e3",
X"a00883a8",
X"80055184",
X"eb3fff75",
X"3483a080",
X"54805383",
X"e39c0852",
X"83e3a008",
X"51fecc3f",
X"80d08054",
X"83b08053",
X"83e39c08",
X"5283e3a0",
X"0851feb7",
X"3f86913f",
X"a2548053",
X"83e3a008",
X"8c800552",
X"80ede851",
X"fea13f86",
X"0b87a883",
X"34800b87",
X"a8823480",
X"0b87a09a",
X"34af0b87",
X"a09634bf",
X"0b87a097",
X"34800b87",
X"a098349f",
X"0b87a099",
X"34800b87",
X"a09b34e0",
X"0b87a889",
X"34a20b87",
X"a8803483",
X"0b87a48f",
X"34820b87",
X"a8813486",
X"3d0d04fd",
X"3d0d83a0",
X"80548053",
X"83e3a008",
X"5283e39c",
X"0851fdbf",
X"3f80d080",
X"5483b080",
X"5383e3a0",
X"085283e3",
X"9c0851fd",
X"aa3fa054",
X"83a08053",
X"83e3a008",
X"5283e39c",
X"0851fd97",
X"3fa05483",
X"a4805383",
X"e3a00852",
X"83e39c08",
X"51fd843f",
X"905483a8",
X"805383e3",
X"a0085283",
X"e39c0851",
X"fcf13f83",
X"e3a43387",
X"a6813485",
X"3d0d0480",
X"3d0d9080",
X"90088106",
X"83e0800c",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fe0676",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70812c81",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870fd",
X"06761007",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"822cbf06",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fe83",
X"0676822b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70882c87",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870f1",
X"ff067688",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"08708b2c",
X"bf0683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"f88fff06",
X"768b2b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"912cbf06",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fc87",
X"ffff0676",
X"912b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"80087088",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"892c8106",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708a2c81",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708b2c",
X"810683e0",
X"800c5182",
X"3d0d04fe",
X"3d0d7481",
X"e629872a",
X"9080a00c",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708105",
X"5434ff11",
X"51f03984",
X"3d0d04fe",
X"3d0d7575",
X"ff195353",
X"5370ff2e",
X"8d387272",
X"70840554",
X"0cff1151",
X"f039843d",
X"0d04fe3d",
X"0d848080",
X"53805288",
X"800a51ff",
X"b33f8180",
X"80538052",
X"82800a51",
X"c63f843d",
X"0d04803d",
X"0d8151fc",
X"bf3f7280",
X"2e8338d2",
X"3f8151fc",
X"dd3f8051",
X"fcd83f80",
X"51fca93f",
X"823d0d04",
X"fd3d0d75",
X"52805480",
X"ff722588",
X"38810bff",
X"80135354",
X"ffbf1251",
X"70992686",
X"38e01252",
X"9e39ff9f",
X"12519971",
X"279538d0",
X"12e01370",
X"54545189",
X"71278838",
X"8f732783",
X"38805273",
X"802e8538",
X"81801252",
X"7181ff06",
X"83e0800c",
X"853d0d04",
X"803d0d84",
X"d8c05180",
X"71708105",
X"53347084",
X"e0c02e09",
X"8106f038",
X"823d0d04",
X"fe3d0d02",
X"97053351",
X"ff863f83",
X"e0800881",
X"ff0683e3",
X"a8085452",
X"8073249b",
X"3883e3c4",
X"08137283",
X"e3c80807",
X"53537173",
X"3483e3a8",
X"08810583",
X"e3a80c84",
X"3d0d04fa",
X"3d0d8280",
X"0a1b5580",
X"57883dfc",
X"05547953",
X"74527851",
X"d69e3f88",
X"3d0d04fe",
X"3d0d83e3",
X"c0085274",
X"51dd833f",
X"83e08008",
X"8c387653",
X"755283e3",
X"c00851c7",
X"3f843d0d",
X"04fe3d0d",
X"83e3c008",
X"53755274",
X"51d7c13f",
X"83e08008",
X"8d387753",
X"765283e3",
X"c00851ff",
X"a23f843d",
X"0d04fe3d",
X"0d83e3c0",
X"0851d6b5",
X"3f83e080",
X"08818080",
X"2e098106",
X"883883c1",
X"8080539b",
X"3983e3c0",
X"0851d699",
X"3f83e080",
X"0880d080",
X"2e098106",
X"933883c1",
X"b0805383",
X"e0800852",
X"83e3c008",
X"51fed83f",
X"843d0d04",
X"803d0dfa",
X"b43f83e0",
X"80088429",
X"80ee8c05",
X"700883e0",
X"800c5182",
X"3d0d04ee",
X"3d0d8043",
X"80428041",
X"80705a5b",
X"fdd23f80",
X"0b83e3a8",
X"0c800b83",
X"e3c80c80",
X"ebe851d1",
X"833f8180",
X"0b83e3c8",
X"0c80ebec",
X"51d0f53f",
X"80d00b83",
X"e3a80c78",
X"30707a07",
X"80257087",
X"2b83e3c8",
X"0c5155f9",
X"a73f83e0",
X"80085280",
X"ebf451d0",
X"cf3f80f8",
X"0b83e3a8",
X"0c788132",
X"70307072",
X"07802570",
X"872b83e3",
X"c80c5156",
X"56fef13f",
X"83e08008",
X"5280ec80",
X"51d0a53f",
X"81a00b83",
X"e3a80c78",
X"82327030",
X"70720780",
X"2570872b",
X"83e3c80c",
X"515683e3",
X"c0085256",
X"d1bf3f83",
X"e0800852",
X"80ec8851",
X"cff63f81",
X"f00b83e3",
X"a80c810b",
X"83e3ac5b",
X"5883e3a8",
X"0882197a",
X"32703070",
X"72078025",
X"70872b83",
X"e3c80c51",
X"578e3d70",
X"55ff1b54",
X"57575799",
X"863f7970",
X"84055b08",
X"51d0f63f",
X"745483e0",
X"80085377",
X"5280ec90",
X"51cfa93f",
X"a81783e3",
X"a80c8118",
X"5877852e",
X"098106ff",
X"b0388390",
X"0b83e3a8",
X"0c788732",
X"70307072",
X"07802570",
X"872b83e3",
X"c80c5156",
X"56f8cd3f",
X"80eca055",
X"83e08008",
X"802e8e38",
X"83e3bc08",
X"51d0a23f",
X"83e08008",
X"55745280",
X"eca851ce",
X"d73f83e0",
X"0b83e3a8",
X"0c788832",
X"70307072",
X"07802570",
X"872b83e3",
X"c80c5157",
X"80ecb452",
X"55ceb53f",
X"868da051",
X"f9853f80",
X"52913d70",
X"525599d8",
X"3f835274",
X"5199d13f",
X"61195978",
X"80258538",
X"80599039",
X"88792585",
X"38885987",
X"39788826",
X"82db3878",
X"822b5580",
X"eac41508",
X"04f6c13f",
X"83e08008",
X"61575575",
X"812e0981",
X"06893883",
X"e0800810",
X"55903975",
X"ff2e0981",
X"06883883",
X"e0800881",
X"2c559075",
X"25853890",
X"55883974",
X"80248338",
X"81557451",
X"f69b3f82",
X"9039f6ad",
X"3f83e080",
X"08610555",
X"74802585",
X"38805588",
X"39877525",
X"83388755",
X"7451f6a6",
X"3f81ee39",
X"60873862",
X"802e81e5",
X"3883e0a4",
X"0883e0a0",
X"0c8bdf0b",
X"83e0a80c",
X"83e3c008",
X"51ffbfd5",
X"3ffae73f",
X"81c73960",
X"56807625",
X"99388af8",
X"0b83e0a8",
X"0c83e3a0",
X"15700852",
X"55ffbfb5",
X"3f740852",
X"91397580",
X"25913883",
X"e3a01508",
X"51ce903f",
X"8052fd19",
X"51b83962",
X"802e818d",
X"3883e3a0",
X"15700883",
X"e3ac0872",
X"0c83e3ac",
X"0cfd1a70",
X"5351558a",
X"f73f83e0",
X"80085680",
X"518aed3f",
X"83e08008",
X"52745187",
X"8b3f7552",
X"80518784",
X"3f80d639",
X"60558075",
X"25b83883",
X"e0ac0883",
X"e0a00c8b",
X"df0b83e0",
X"a80c83e3",
X"bc0851ff",
X"bebf3f83",
X"e3bc0851",
X"ffbbd93f",
X"83e08008",
X"81ff0670",
X"5255f5b1",
X"3f74802e",
X"9c388155",
X"a0397480",
X"25933883",
X"e3bc0851",
X"cd813f80",
X"51f5963f",
X"84396287",
X"387a802e",
X"fa8a3880",
X"557483e0",
X"800c943d",
X"0d04fe3d",
X"0df5943f",
X"83e08008",
X"802e8638",
X"805180f7",
X"39f5993f",
X"83e08008",
X"80eb38f5",
X"b93f83e0",
X"8008802e",
X"aa388151",
X"f2f63fef",
X"ef3f800b",
X"83e3a80c",
X"f9b93f83",
X"e0800853",
X"ff0b83e3",
X"a80cf1db",
X"3f72be38",
X"7251f2d4",
X"3fbc39f4",
X"f03f83e0",
X"8008802e",
X"b1388151",
X"f2c23fef",
X"bb3f8af8",
X"0b83e0a8",
X"0c83e3ac",
X"0851ffbd",
X"843fff0b",
X"83e3a80c",
X"f1a53f83",
X"e3ac0852",
X"80518594",
X"3f8151f5",
X"d13f843d",
X"0d04fc3d",
X"0d908080",
X"52868480",
X"8051cfd6",
X"3f83e080",
X"0880c338",
X"88df3f80",
X"efe051d4",
X"973f83e0",
X"8008559c",
X"800a5480",
X"c0805380",
X"ecbc5283",
X"e0800851",
X"f79f3f83",
X"e3c00853",
X"80eccc52",
X"7451cee0",
X"3f83e080",
X"088438f7",
X"ad3f8151",
X"f4f83f92",
X"ea3f8151",
X"f4f03ffe",
X"913ffc39",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"0280ecd8",
X"0b83e0a4",
X"0c80ecdc",
X"0b83e09c",
X"0c80ece0",
X"0b83e0ac",
X"0c83e08c",
X"08fc050c",
X"800b83e3",
X"ac0b83e0",
X"8c08f805",
X"0c83e08c",
X"08f4050c",
X"cdb83f83",
X"e0800886",
X"05fc0683",
X"e08c08f0",
X"050c0283",
X"e08c08f0",
X"0508310d",
X"833d7083",
X"e08c08f8",
X"05087084",
X"0583e08c",
X"08f8050c",
X"0c51c9ff",
X"3f83e08c",
X"08f40508",
X"810583e0",
X"8c08f405",
X"0c83e08c",
X"08f40508",
X"862e0981",
X"06ffad38",
X"86948080",
X"51ecd23f",
X"ff0b83e3",
X"a80c800b",
X"83e3c80c",
X"84d8c00b",
X"83e3c40c",
X"8151effc",
X"3f8151f0",
X"a13f8051",
X"f09c3f81",
X"51f0c23f",
X"8151f197",
X"3f8251f0",
X"e53f8051",
X"f1bb3f80",
X"c6885280",
X"51c7be3f",
X"fdc03f83",
X"e08c08fc",
X"05080d80",
X"0b83e080",
X"0c873d0d",
X"83e08c0c",
X"04803d0d",
X"81ff5180",
X"0b83e3d4",
X"1234ff11",
X"5170f438",
X"823d0d04",
X"ff3d0d73",
X"70335351",
X"81113371",
X"34718112",
X"34833d0d",
X"04fb3d0d",
X"77795656",
X"80707155",
X"55527175",
X"25ac3872",
X"16703370",
X"147081ff",
X"06555151",
X"51717427",
X"89388112",
X"7081ff06",
X"53517181",
X"147083ff",
X"ff065552",
X"54747324",
X"d6387183",
X"e0800c87",
X"3d0d04fc",
X"3d0d7655",
X"c0eb3f83",
X"e0800880",
X"2ef63883",
X"e5f00886",
X"057081ff",
X"065253ff",
X"beec3f84",
X"39fb833f",
X"c0cb3f83",
X"e0800881",
X"2ef33880",
X"54731553",
X"ffbfb23f",
X"83e08008",
X"73348114",
X"5473852e",
X"098106e9",
X"388439fa",
X"d93fc0a1",
X"3f83e080",
X"08802ef3",
X"38743383",
X"e3d43481",
X"153383e3",
X"d5348215",
X"3383e3d6",
X"34831533",
X"83e3d734",
X"845283e3",
X"d451febd",
X"3f83e080",
X"0881ff06",
X"84163356",
X"5372752e",
X"0981068d",
X"38ffbf96",
X"3f83e080",
X"08802e9a",
X"3883e5f0",
X"08a82e09",
X"81068938",
X"860b83e5",
X"f00c8739",
X"a80b83e5",
X"f00c80e4",
X"51efd83f",
X"863d0d04",
X"f43d0d7e",
X"60595580",
X"5d807582",
X"2b7183e5",
X"f4120c83",
X"e688175b",
X"5b577679",
X"3477772e",
X"83b23876",
X"527751c8",
X"cf3f8e3d",
X"fc055490",
X"5383e5dc",
X"527751c8",
X"8b3f7c56",
X"75902e09",
X"81068390",
X"3883e5dc",
X"51fd993f",
X"83e5de51",
X"fd923f83",
X"e5e051fd",
X"8b3f7683",
X"e5ec0c77",
X"51c5d63f",
X"80eaf852",
X"83e08008",
X"51ffb592",
X"3f83e080",
X"08812e09",
X"810680d3",
X"387683e6",
X"840c820b",
X"83e5dc34",
X"ff960b83",
X"e5dd3477",
X"51c89e3f",
X"83e08008",
X"5583e080",
X"08772588",
X"3883e080",
X"088f0555",
X"74842c70",
X"83ffff06",
X"70882a58",
X"51557583",
X"e5de3474",
X"83e5df34",
X"7683e5e0",
X"34ff800b",
X"83e5e134",
X"818f3983",
X"e5dc3383",
X"e5dd3371",
X"882b0756",
X"5b7483ff",
X"ff2e0981",
X"0680e738",
X"fe800b83",
X"e6840c81",
X"0b83e5ec",
X"0cff0b83",
X"e5dc34ff",
X"0b83e5dd",
X"347751c7",
X"ac3f83e0",
X"800883e6",
X"8c0c83e0",
X"80085583",
X"e0800880",
X"25883883",
X"e080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583e5de",
X"347483e5",
X"df347683",
X"e5e034ff",
X"800b83e5",
X"e134810b",
X"83e5eb34",
X"a4397485",
X"962e0981",
X"0680fd38",
X"7583e684",
X"0c7751c6",
X"e13f83e5",
X"eb3383e0",
X"80080755",
X"7483e5eb",
X"3483e5eb",
X"33810655",
X"74802e83",
X"38845783",
X"e5e03383",
X"e5e13371",
X"882b0756",
X"5c748180",
X"2e098106",
X"a13883e5",
X"de3383e5",
X"df337188",
X"2b07565b",
X"ad807527",
X"87387682",
X"07579c39",
X"76810757",
X"96397482",
X"802e0981",
X"06873876",
X"83075787",
X"397481ff",
X"268a3877",
X"83e5f41b",
X"0c767934",
X"8e3d0d04",
X"803d0d72",
X"842983e5",
X"f4057008",
X"83e0800c",
X"51823d0d",
X"04fe3d0d",
X"800b83e5",
X"d80c800b",
X"83e5d40c",
X"ff0b83e3",
X"d00ca80b",
X"83e5f00c",
X"ae51ffb9",
X"bd3f800b",
X"83e5f454",
X"52807370",
X"8405550c",
X"81125271",
X"842e0981",
X"06ef3884",
X"3d0d04fe",
X"3d0d7402",
X"84059605",
X"22535371",
X"802e9738",
X"72708105",
X"543351ff",
X"b9c73fff",
X"127083ff",
X"ff065152",
X"e639843d",
X"0d04fe3d",
X"0d029205",
X"225382ac",
X"51eaf03f",
X"80c351ff",
X"b9a33f81",
X"9651eae3",
X"3f725283",
X"e3d451ff",
X"b23f7252",
X"83e3d451",
X"f8f73f83",
X"e0800881",
X"ff0651ff",
X"b8ff3f84",
X"3d0d04ff",
X"b13d0d80",
X"d13df805",
X"51f9a03f",
X"83e5d808",
X"810583e5",
X"d80c80cf",
X"3d33cf11",
X"7081ff06",
X"51565674",
X"832688ec",
X"38758f06",
X"ff055675",
X"83e3d008",
X"2e9b3875",
X"83269638",
X"7583e3d0",
X"0c758429",
X"83e5f405",
X"70085355",
X"7551fa9c",
X"3f807624",
X"88c83875",
X"842983e5",
X"f4055574",
X"08802e88",
X"b93883e3",
X"d0088429",
X"83e5f405",
X"70080288",
X"0582b905",
X"33525b55",
X"7480d22e",
X"84b03874",
X"80d22490",
X"3874bf2e",
X"9c387480",
X"d02e81d7",
X"3887f739",
X"7480d32e",
X"80d23874",
X"80d72e81",
X"c63887e6",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055656",
X"ffb7fa3f",
X"80c151ff",
X"b7b33ff6",
X"f03f860b",
X"83e3d434",
X"815283e3",
X"d451ffb8",
X"d53f8151",
X"fde43f74",
X"8938860b",
X"83e5f00c",
X"8739a80b",
X"83e5f00c",
X"ffb7c63f",
X"80c151ff",
X"b6ff3ff6",
X"bc3f900b",
X"83e5eb33",
X"81065656",
X"74802e83",
X"38985683",
X"e5e03383",
X"e5e13371",
X"882b0756",
X"59748180",
X"2e098106",
X"9c3883e5",
X"de3383e5",
X"df337188",
X"2b075657",
X"ad807527",
X"8c387581",
X"80075685",
X"3975a007",
X"567583e3",
X"d434ff0b",
X"83e3d534",
X"e00b83e3",
X"d634800b",
X"83e3d734",
X"845283e3",
X"d451ffb7",
X"c93f8451",
X"869d3902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"5659ffb6",
X"b83f7951",
X"c1a83f83",
X"e0800880",
X"2e8b3880",
X"ce51ffb5",
X"e43f85f2",
X"3980c151",
X"ffb5da3f",
X"ffb6ce3f",
X"ffb5823f",
X"83e68408",
X"58837525",
X"9b3883e5",
X"e03383e5",
X"e1337188",
X"2b07fc17",
X"71297a05",
X"8380055a",
X"51578d39",
X"74818029",
X"18ff8005",
X"58818057",
X"80567676",
X"2e9338ff",
X"b5b33f83",
X"e0800883",
X"e3d41734",
X"811656ea",
X"39ffb5a1",
X"3f83e080",
X"0881ff06",
X"775383e3",
X"d45256f4",
X"e03f83e0",
X"800881ff",
X"06557575",
X"2e098106",
X"818a38ff",
X"b59f3f80",
X"c151ffb4",
X"d83fffb5",
X"cc3f7752",
X"7951ffbf",
X"b73f805e",
X"80d13dfd",
X"f4055476",
X"5383e3d4",
X"527951ff",
X"bdc33f02",
X"82b90533",
X"55815874",
X"80d72e09",
X"8106bd38",
X"80d13dfd",
X"f0055476",
X"538f3d70",
X"537a5259",
X"ffbec93f",
X"80567676",
X"2ea23875",
X"1983e3d4",
X"17337133",
X"70723270",
X"30708025",
X"70307e06",
X"811d5d5e",
X"51515152",
X"5b55db39",
X"82ac51e5",
X"aa3f7780",
X"2e863880",
X"c3518439",
X"80ce51ff",
X"b3d33fff",
X"b4c73fff",
X"b2fb3f83",
X"dd390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290559",
X"5580705d",
X"59ffb3ed",
X"3f80c151",
X"ffb3a63f",
X"83e5ec08",
X"792e82de",
X"3883e68c",
X"0880fc05",
X"5580fd52",
X"745186d7",
X"3f83e080",
X"085b7782",
X"24b238ff",
X"1870872b",
X"83ffff80",
X"0680eeac",
X"0583e3d4",
X"59575581",
X"80557570",
X"81055733",
X"77708105",
X"5934ff15",
X"7081ff06",
X"515574ea",
X"38828d39",
X"7782e82e",
X"81ab3877",
X"82e92e09",
X"810681b2",
X"3880ece4",
X"51ffb9a8",
X"3f785877",
X"87327030",
X"70720780",
X"257a8a32",
X"70307072",
X"07802573",
X"0753545a",
X"51575575",
X"802e9738",
X"78782692",
X"38a00b83",
X"e3d41a34",
X"81197081",
X"ff065a55",
X"eb398118",
X"7081ff06",
X"59558a78",
X"27ffbc38",
X"8f5883e3",
X"cf183383",
X"e3d41934",
X"ff187081",
X"ff065955",
X"778426ea",
X"38905880",
X"0b83e3d4",
X"19348118",
X"7081ff06",
X"70982b52",
X"59557480",
X"25e93880",
X"c6557a85",
X"8f248438",
X"80c25574",
X"83e3d434",
X"80f10b83",
X"e3d73481",
X"0b83e3d8",
X"347a83e3",
X"d5347a88",
X"2c557483",
X"e3d63480",
X"cb3982f0",
X"782580c4",
X"387780fd",
X"29fd97d3",
X"05527951",
X"ffbbe53f",
X"80d13dfd",
X"ec055480",
X"fd5383e3",
X"d4527951",
X"ffbb9d3f",
X"7b811959",
X"567580fc",
X"24833878",
X"5877882c",
X"557483e4",
X"d1347783",
X"e4d23475",
X"83e4d334",
X"81805980",
X"cc3983e6",
X"84085783",
X"78259b38",
X"83e5e033",
X"83e5e133",
X"71882b07",
X"fc1a7129",
X"79058380",
X"05595159",
X"8d397781",
X"802917ff",
X"80055781",
X"80597652",
X"7951ffba",
X"f33f80d1",
X"3dfdec05",
X"54785383",
X"e3d45279",
X"51ffbaac",
X"3f7851f6",
X"b93fffb0",
X"e43fffaf",
X"983f8b39",
X"83e5d408",
X"810583e5",
X"d40c80d1",
X"3d0d04f6",
X"da3febaa",
X"3ff939fc",
X"3d0d7678",
X"71842983",
X"e5f40570",
X"08515353",
X"53709e38",
X"80ce7234",
X"80cf0b81",
X"133480ce",
X"0b821334",
X"80c50b83",
X"13347084",
X"133480e7",
X"3983e688",
X"13335480",
X"d2723473",
X"822a7081",
X"06515180",
X"cf537084",
X"3880d753",
X"72811334",
X"a00b8213",
X"34738306",
X"5170812e",
X"9e387081",
X"24883870",
X"802e8f38",
X"9f397082",
X"2e923870",
X"832e9238",
X"933980d8",
X"558e3980",
X"d3558939",
X"80cd5584",
X"3980c455",
X"74831334",
X"80c40b84",
X"1334800b",
X"85133486",
X"3d0d04fd",
X"3d0d7553",
X"80730c80",
X"0b84140c",
X"800b8814",
X"0c87a680",
X"337081ff",
X"0670812a",
X"81327181",
X"32718106",
X"71810631",
X"84180c55",
X"5670832a",
X"81327182",
X"2a813271",
X"81067181",
X"0631770c",
X"52545151",
X"87a09033",
X"70098106",
X"88150c51",
X"853d0d04",
X"fe3d0d74",
X"76545271",
X"51ffa03f",
X"72812ea2",
X"38817326",
X"8d387282",
X"2eab3872",
X"832e9f38",
X"e6397108",
X"e2388412",
X"08dd3888",
X"1208d838",
X"a0398812",
X"08812e09",
X"8106cc38",
X"94398812",
X"08812e8d",
X"38710889",
X"38841208",
X"802effb7",
X"38843d0d",
X"04fc3d0d",
X"76785354",
X"81538055",
X"87397110",
X"73105452",
X"73722651",
X"72802ea7",
X"3870802e",
X"86387180",
X"25e83872",
X"802e9838",
X"71742689",
X"38737231",
X"75740756",
X"5472812a",
X"72812a53",
X"53e53973",
X"51788338",
X"74517083",
X"e0800c86",
X"3d0d04fe",
X"3d0d8053",
X"75527451",
X"ffa33f84",
X"3d0d04fe",
X"3d0d8153",
X"75527451",
X"ff933f84",
X"3d0d04fb",
X"3d0d7779",
X"55558056",
X"74762586",
X"38743055",
X"81567380",
X"25883873",
X"30768132",
X"57548053",
X"73527451",
X"fee73f83",
X"e0800854",
X"75802e87",
X"3883e080",
X"08305473",
X"83e0800c",
X"873d0d04",
X"fa3d0d78",
X"7a575580",
X"57747725",
X"86387430",
X"55815775",
X"9f2c5481",
X"53757432",
X"74315274",
X"51feaa3f",
X"83e08008",
X"5476802e",
X"873883e0",
X"80083054",
X"7383e080",
X"0c883d0d",
X"04ff3d0d",
X"73527183",
X"e694082e",
X"a63871a0",
X"0a079080",
X"9c0c9080",
X"8c085170",
X"802ef738",
X"800b9080",
X"9c0c9080",
X"8c085170",
X"f9387183",
X"e6940c83",
X"3d0d04ff",
X"0b83e694",
X"0c818080",
X"0b83e690",
X"0c800b83",
X"e0800c04",
X"fc3d0d76",
X"028405a2",
X"05220288",
X"05a60522",
X"7a545555",
X"55ff9e3f",
X"72802ea3",
X"3883e690",
X"08145271",
X"33757081",
X"05573481",
X"147083ff",
X"ff06ff15",
X"7083ffff",
X"06565255",
X"52da3980",
X"0b83e080",
X"0c863d0d",
X"04f73d0d",
X"7b7d7f11",
X"58555980",
X"5573762e",
X"b13883e6",
X"90088b3d",
X"59577419",
X"703375fc",
X"06197008",
X"5d768306",
X"7b075354",
X"54517271",
X"3479720c",
X"81148116",
X"56547376",
X"2e098106",
X"d938800b",
X"83e0800c",
X"8b3d0d04",
X"803d0d83",
X"e6940890",
X"0a079080",
X"9c0c9080",
X"8c085170",
X"802ef738",
X"800b9080",
X"9c0c9080",
X"8c085170",
X"f938823d",
X"0d040000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"000025b9",
X"000025fa",
X"0000261c",
X"00002643",
X"00002643",
X"00002643",
X"00002643",
X"000026b4",
X"00002706",
X"25732025",
X"73000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"6e616d65",
X"20000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"000035a4",
X"000035a8",
X"000035b0",
X"000035bc",
X"000035c8",
X"000035d4",
X"000035e0",
X"000035e4",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
