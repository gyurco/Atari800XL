-- megafunction wizard: %ALTIOBUF%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altiobuf_bidir 

-- ============================================================
-- File Name: altiobuf.vhd
-- Megafunction Name(s):
-- 			altiobuf_bidir
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 14.0.0 Build 200 06/17/2014 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus II License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


--altiobuf_bidir CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" ENABLE_BUS_HOLD="FALSE" NUMBER_OF_CHANNELS=4 OPEN_DRAIN_OUTPUT="FALSE" USE_DIFFERENTIAL_MODE="TRUE" USE_DYNAMIC_TERMINATION_CONTROL="FALSE" USE_TERMINATION_CONTROL="FALSE" datain dataio dataio_b dataout oe oe_b
--VERSION_BEGIN 14.0 cbx_altiobuf_bidir 2014:06:05:09:45:41:SJ cbx_mgl 2014:06:05:10:17:12:SJ cbx_stratixiii 2014:06:05:09:45:41:SJ cbx_stratixv 2014:06:05:09:45:41:SJ  VERSION_END

 LIBRARY cyclonev;
 USE cyclonev.all;

--synthesis_resources = cyclonev_io_ibuf 4 cyclonev_io_obuf 8 cyclonev_pseudo_diff_out 4 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altiobuf_iobuf_bidir_lup IS 
	 PORT 
	 ( 
		 datain	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 dataio	:	INOUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 dataio_b	:	INOUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 dataout	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 oe	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 oe_b	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '1')
	 ); 
 END altiobuf_iobuf_bidir_lup;

 ARCHITECTURE RTL OF altiobuf_iobuf_bidir_lup IS

	 SIGNAL  wire_ibufa_i	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_ibufa_ibar	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_ibufa_o	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_obuf_ba_o	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_obuf_ba_oe	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_obufa_o	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_obufa_oe	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_pseudo_diffa_w_lg_oebout3w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_pseudo_diffa_w_lg_oeout2w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_pseudo_diffa_i	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_pseudo_diffa_o	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_pseudo_diffa_obar	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_pseudo_diffa_oebout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_pseudo_diffa_oein	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_pseudo_diffa_oeout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_oe1w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 COMPONENT  cyclonev_io_ibuf
	 GENERIC 
	 (
		bus_hold	:	STRING := "false";
		differential_mode	:	STRING := "false";
		simulate_z_as	:	STRING := "z";
		lpm_type	:	STRING := "cyclonev_io_ibuf"
	 );
	 PORT
	 ( 
		dynamicterminationcontrol	:	IN STD_LOGIC := '0';
		i	:	IN STD_LOGIC := '0';
		ibar	:	IN STD_LOGIC := '0';
		o	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  cyclonev_io_obuf
	 GENERIC 
	 (
		bus_hold	:	STRING := "false";
		open_drain_output	:	STRING := "false";
		shift_series_termination_control	:	STRING := "false";
		lpm_type	:	STRING := "cyclonev_io_obuf"
	 );
	 PORT
	 ( 
		dynamicterminationcontrol	:	IN STD_LOGIC := '0';
		i	:	IN STD_LOGIC := '0';
		o	:	OUT STD_LOGIC;
		obar	:	OUT STD_LOGIC;
		oe	:	IN STD_LOGIC := '1';
		parallelterminationcontrol	:	IN STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
		seriesterminationcontrol	:	IN STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  cyclonev_pseudo_diff_out
	 PORT
	 ( 
		dtc	:	OUT STD_LOGIC;
		dtcbar	:	OUT STD_LOGIC;
		dtcin	:	IN STD_LOGIC := '0';
		i	:	IN STD_LOGIC := '0';
		o	:	OUT STD_LOGIC;
		obar	:	OUT STD_LOGIC;
		oebout	:	OUT STD_LOGIC;
		oein	:	IN STD_LOGIC := '0';
		oeout	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	loop0 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_oe1w(i) <= NOT oe(i);
	END GENERATE loop0;
	dataio <= wire_obufa_o;
	dataio_b <= wire_obuf_ba_o;
	dataout <= wire_ibufa_o;
	wire_ibufa_i <= dataio;
	wire_ibufa_ibar <= dataio_b;
	loop1 : FOR i IN 0 TO 3 GENERATE 
	  ibufa :  cyclonev_io_ibuf
	  GENERIC MAP (
		bus_hold => "false",
		differential_mode => "true"
	  )
	  PORT MAP ( 
		i => wire_ibufa_i(i),
		ibar => wire_ibufa_ibar(i),
		o => wire_ibufa_o(i)
	  );
	END GENERATE loop1;
	wire_obuf_ba_oe <= wire_pseudo_diffa_w_lg_oebout3w;
	loop2 : FOR i IN 0 TO 3 GENERATE 
	  obuf_ba :  cyclonev_io_obuf
	  GENERIC MAP (
		bus_hold => "false",
		open_drain_output => "false"
	  )
	  PORT MAP ( 
		i => wire_pseudo_diffa_obar(i),
		o => wire_obuf_ba_o(i),
		oe => wire_obuf_ba_oe(i)
	  );
	END GENERATE loop2;
	wire_obufa_oe <= wire_pseudo_diffa_w_lg_oeout2w;
	loop3 : FOR i IN 0 TO 3 GENERATE 
	  obufa :  cyclonev_io_obuf
	  GENERIC MAP (
		bus_hold => "false",
		open_drain_output => "false"
	  )
	  PORT MAP ( 
		i => wire_pseudo_diffa_o(i),
		o => wire_obufa_o(i),
		oe => wire_obufa_oe(i)
	  );
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 3 GENERATE 
		wire_pseudo_diffa_w_lg_oebout3w(i) <= NOT wire_pseudo_diffa_oebout(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 3 GENERATE 
		wire_pseudo_diffa_w_lg_oeout2w(i) <= NOT wire_pseudo_diffa_oeout(i);
	END GENERATE loop5;
	wire_pseudo_diffa_i <= datain;
	wire_pseudo_diffa_oein <= wire_w_lg_oe1w;
	loop6 : FOR i IN 0 TO 3 GENERATE 
	  pseudo_diffa :  cyclonev_pseudo_diff_out
	  PORT MAP ( 
		i => wire_pseudo_diffa_i(i),
		o => wire_pseudo_diffa_o(i),
		obar => wire_pseudo_diffa_obar(i),
		oebout => wire_pseudo_diffa_oebout(i),
		oein => wire_pseudo_diffa_oein(i),
		oeout => wire_pseudo_diffa_oeout(i)
	  );
	END GENERATE loop6;

 END RTL; --altiobuf_iobuf_bidir_lup
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY altiobuf IS
	PORT
	(
		datain		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		oe		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		oe_b		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		dataio		: INOUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		dataio_b		: INOUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		dataout		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
END altiobuf;


ARCHITECTURE RTL OF altiobuf IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (3 DOWNTO 0);



	COMPONENT altiobuf_iobuf_bidir_lup
	PORT (
			datain	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			oe	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			oe_b	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			dataout	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			dataio	: INOUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			dataio_b	: INOUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	dataout    <= sub_wire0(3 DOWNTO 0);

	altiobuf_iobuf_bidir_lup_component : altiobuf_iobuf_bidir_lup
	PORT MAP (
		datain => datain,
		oe => oe,
		oe_b => oe_b,
		dataout => sub_wire0,
		dataio => dataio,
		dataio_b => dataio_b
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: enable_bus_hold STRING "FALSE"
-- Retrieval info: CONSTANT: left_shift_series_termination_control STRING "FALSE"
-- Retrieval info: CONSTANT: number_of_channels NUMERIC "4"
-- Retrieval info: CONSTANT: open_drain_output STRING "FALSE"
-- Retrieval info: CONSTANT: use_differential_mode STRING "TRUE"
-- Retrieval info: CONSTANT: use_dynamic_termination_control STRING "FALSE"
-- Retrieval info: CONSTANT: use_termination_control STRING "FALSE"
-- Retrieval info: USED_PORT: datain 0 0 4 0 INPUT NODEFVAL "datain[3..0]"
-- Retrieval info: USED_PORT: dataio 0 0 4 0 BIDIR NODEFVAL "dataio[3..0]"
-- Retrieval info: USED_PORT: dataio_b 0 0 4 0 BIDIR NODEFVAL "dataio_b[3..0]"
-- Retrieval info: USED_PORT: dataout 0 0 4 0 OUTPUT NODEFVAL "dataout[3..0]"
-- Retrieval info: USED_PORT: oe 0 0 4 0 INPUT NODEFVAL "oe[3..0]"
-- Retrieval info: USED_PORT: oe_b 0 0 4 0 INPUT NODEFVAL "oe_b[3..0]"
-- Retrieval info: CONNECT: @datain 0 0 4 0 datain 0 0 4 0
-- Retrieval info: CONNECT: @oe 0 0 4 0 oe 0 0 4 0
-- Retrieval info: CONNECT: @oe_b 0 0 4 0 oe_b 0 0 4 0
-- Retrieval info: CONNECT: dataio 0 0 4 0 @dataio 0 0 4 0
-- Retrieval info: CONNECT: dataio_b 0 0 4 0 @dataio_b 0 0 4 0
-- Retrieval info: CONNECT: dataout 0 0 4 0 @dataout 0 0 4 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altiobuf.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altiobuf.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altiobuf.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altiobuf.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altiobuf_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
