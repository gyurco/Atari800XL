
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f2",
X"dc738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80f6",
X"a00c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f2",
X"9d2d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580f1dc",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80dbac04",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"775193b0",
X"3f83e080",
X"0880d638",
X"78902e09",
X"810680cd",
X"3802ab05",
X"3380f6a8",
X"0b80f6a8",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ac388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"5696800a",
X"52775192",
X"df3f83e0",
X"80088638",
X"78752e85",
X"38805685",
X"39811733",
X"567583e0",
X"800c8e3d",
X"0d04fc3d",
X"0d767052",
X"55b3943f",
X"83e08008",
X"15ff0554",
X"73752e8e",
X"38733353",
X"72ae2e86",
X"38ff1454",
X"ef397752",
X"811451b2",
X"ac3f83e0",
X"80083070",
X"83e08008",
X"07802583",
X"e0800c53",
X"863d0d04",
X"fc3d0d76",
X"70525599",
X"cc3f83e0",
X"80085481",
X"5383e080",
X"0880c738",
X"7451998f",
X"3f83e080",
X"080b0b80",
X"f49c5383",
X"e0800852",
X"53ff8f3f",
X"83e08008",
X"a5380b0b",
X"80f4a052",
X"7251fefe",
X"3f83e080",
X"0894380b",
X"0b80f4a4",
X"527251fe",
X"ed3f83e0",
X"8008802e",
X"83388154",
X"73537283",
X"e0800c86",
X"3d0d04fd",
X"3d0d7570",
X"525498e5",
X"3f815383",
X"e0800898",
X"38735198",
X"ae3f83e0",
X"a0085283",
X"e0800851",
X"feb43f83",
X"e0800853",
X"7283e080",
X"0c853d0d",
X"04e03d0d",
X"a33d0870",
X"525e8ed3",
X"3f83e080",
X"0833943d",
X"56547394",
X"3880f9ac",
X"52745184",
X"c7397d52",
X"785191d6",
X"3f84d139",
X"7d518ebb",
X"3f83e080",
X"08527451",
X"8deb3f83",
X"e0a80852",
X"933d7052",
X"5d94c63f",
X"83e08008",
X"59800b83",
X"e0800855",
X"5b83e080",
X"087b2e94",
X"38811b74",
X"525b97c8",
X"3f83e080",
X"085483e0",
X"8008ee38",
X"805aff7a",
X"437a427a",
X"415f7909",
X"709f2c7b",
X"065b547a",
X"7a248438",
X"ff1b5af6",
X"1a700970",
X"9f2c7206",
X"7bff125a",
X"5a525555",
X"80752595",
X"38765197",
X"873f83e0",
X"800876ff",
X"18585557",
X"738024ed",
X"38747f2e",
X"873880c2",
X"d53f745f",
X"78ff1b70",
X"585d5880",
X"7a259538",
X"775196dc",
X"3f83e080",
X"0876ff18",
X"58555873",
X"8024ed38",
X"800b83e7",
X"c00c800b",
X"83e7e40c",
X"0b0b80f4",
X"a8518bae",
X"3f81800b",
X"83e7e40c",
X"0b0b80f4",
X"b0518b9e",
X"3fa80b83",
X"e7c00c76",
X"802e80e8",
X"3883e7c0",
X"08777932",
X"70307072",
X"07802570",
X"872b83e7",
X"e40c5156",
X"78535656",
X"968f3f83",
X"e0800880",
X"2e8a380b",
X"0b80f4b8",
X"518ae33f",
X"765195cf",
X"3f83e080",
X"08520b0b",
X"80f5c451",
X"8ad03f76",
X"5195d53f",
X"83e08008",
X"83e7c008",
X"55577574",
X"258638a8",
X"1656f739",
X"7583e7c0",
X"0c86f076",
X"24ff9438",
X"87980b83",
X"e7c00c77",
X"802eb738",
X"7751958b",
X"3f83e080",
X"08785255",
X"95ab3f0b",
X"0b80f4c0",
X"5483e080",
X"088f3887",
X"39807634",
X"fd95390b",
X"0b80f4bc",
X"54745373",
X"520b0b80",
X"f4905189",
X"e93f8054",
X"0b0b80f6",
X"9c5189de",
X"3f811454",
X"73a82e09",
X"8106ed38",
X"868da051",
X"beca3f80",
X"52903d70",
X"525480e0",
X"a43f8352",
X"735180e0",
X"9c3f6180",
X"2e80ff38",
X"7b5473ff",
X"2e963878",
X"802e8180",
X"38785194",
X"ab3f83e0",
X"8008ff15",
X"5559e739",
X"78802e80",
X"eb387851",
X"94a73f83",
X"e0800880",
X"2efc8338",
X"785193ef",
X"3f83e080",
X"08520b0b",
X"80f49851",
X"abce3f83",
X"e08008a4",
X"387c51ad",
X"863f83e0",
X"80085574",
X"ff165654",
X"807425fb",
X"ee38741d",
X"70335556",
X"73af2efe",
X"c838e839",
X"785193ad",
X"3f83e080",
X"08527c51",
X"acbd3ffb",
X"ce397f88",
X"29601005",
X"7a056105",
X"5afbff39",
X"a23d0d04",
X"803d0d90",
X"80f83370",
X"81ff0670",
X"842a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"a80b9080",
X"f834b80b",
X"9080f834",
X"7083e080",
X"0c823d0d",
X"04803d0d",
X"9080f833",
X"7081ff06",
X"70852a81",
X"32708106",
X"51515151",
X"70802e8d",
X"38980b90",
X"80f834b8",
X"0b9080f8",
X"347083e0",
X"800c823d",
X"0d04930b",
X"9080fc34",
X"ff0b9080",
X"e83404ff",
X"3d0d028f",
X"05335280",
X"0b9080fc",
X"348a51bc",
X"9f3fdf3f",
X"80f80b90",
X"80e03480",
X"0b9080c8",
X"34fa1252",
X"719080c0",
X"34800b90",
X"80d83471",
X"9080d034",
X"9080f852",
X"807234b8",
X"7234833d",
X"0d04803d",
X"0d028b05",
X"33517090",
X"80f434fe",
X"bf3f83e0",
X"8008802e",
X"f638823d",
X"0d04803d",
X"0d853980",
X"c5ea3ffe",
X"d83f83e0",
X"8008802e",
X"f2389080",
X"f4337081",
X"ff0683e0",
X"800c5182",
X"3d0d0480",
X"3d0da30b",
X"9080fc34",
X"ff0b9080",
X"e8349080",
X"f851a871",
X"34b87134",
X"823d0d04",
X"803d0d90",
X"80fc3370",
X"81c00670",
X"30708025",
X"83e0800c",
X"51515182",
X"3d0d0480",
X"3d0d9080",
X"f8337081",
X"ff067083",
X"2a813270",
X"81065151",
X"51517080",
X"2ee838b0",
X"0b9080f8",
X"34b80b90",
X"80f83482",
X"3d0d0480",
X"3d0d9080",
X"ac088106",
X"83e0800c",
X"823d0d04",
X"fd3d0d75",
X"77545480",
X"73259438",
X"73708105",
X"55335280",
X"f4c45185",
X"a13fff13",
X"53e93985",
X"3d0d04f6",
X"3d0d7c7e",
X"60625a5d",
X"5b568059",
X"81558539",
X"747a2955",
X"74527551",
X"80dd853f",
X"83e08008",
X"7a27ed38",
X"74802e80",
X"e0387452",
X"755180dc",
X"ef3f83e0",
X"80087553",
X"76525480",
X"dcf23f83",
X"e080087a",
X"53755256",
X"80dcd53f",
X"83e08008",
X"7930707b",
X"079f2a70",
X"77802407",
X"51515455",
X"72873883",
X"e08008c2",
X"38768118",
X"b0165558",
X"58897425",
X"8b38b714",
X"537a8538",
X"80d71453",
X"72783481",
X"1959ff9c",
X"39807734",
X"8c3d0d04",
X"f73d0d7b",
X"7d7f6202",
X"9005bb05",
X"33575956",
X"5a5ab058",
X"728338a0",
X"58757070",
X"81055233",
X"71595455",
X"90398074",
X"258e38ff",
X"14777081",
X"05593354",
X"5472ef38",
X"73ff1555",
X"53807325",
X"89387752",
X"7951782d",
X"ef397533",
X"75575372",
X"802e9038",
X"72527951",
X"782d7570",
X"81055733",
X"53ed398b",
X"3d0d04ee",
X"3d0d6466",
X"69697070",
X"81055233",
X"5b4a5c5e",
X"5e76802e",
X"82f93876",
X"a52e0981",
X"0682e038",
X"80704167",
X"70708105",
X"5233714a",
X"59575f76",
X"b02e0981",
X"068c3875",
X"70810557",
X"33764857",
X"815fd017",
X"56758926",
X"80da3876",
X"675c5980",
X"5c933977",
X"8a2480c3",
X"387b8a29",
X"187b7081",
X"055d335a",
X"5cd01970",
X"81ff0658",
X"58897727",
X"a438ff9f",
X"197081ff",
X"06ffa91b",
X"5a515685",
X"76279238",
X"ffbf1970",
X"81ff0651",
X"56758526",
X"8a38c919",
X"58778025",
X"ffb9387a",
X"477b4078",
X"81ff0657",
X"7680e42e",
X"80e53876",
X"80e424a7",
X"387680d8",
X"2e818638",
X"7680d824",
X"90387680",
X"2e81cc38",
X"76a52e81",
X"b63881b9",
X"397680e3",
X"2e818c38",
X"81af3976",
X"80f52e9b",
X"387680f5",
X"248b3876",
X"80f32e81",
X"81388199",
X"397680f8",
X"2e80ca38",
X"818f3991",
X"3d705557",
X"80538a52",
X"79841b71",
X"08535b56",
X"fbfd3f76",
X"55ab3979",
X"841b7108",
X"943d705b",
X"5b525b56",
X"7580258c",
X"38753056",
X"ad783402",
X"80c10557",
X"76548053",
X"8a527551",
X"fbd13f77",
X"557e54b8",
X"39913d70",
X"557780d8",
X"32703070",
X"80255651",
X"58569052",
X"79841b71",
X"08535b57",
X"fbad3f75",
X"55db3979",
X"841b8312",
X"33545b56",
X"98397984",
X"1b710857",
X"5b568054",
X"7f537c52",
X"7d51fc9c",
X"3f873976",
X"527d517c",
X"2d667033",
X"58810547",
X"fd833994",
X"3d0d0472",
X"83e0900c",
X"7183e094",
X"0c04fb3d",
X"0d883d70",
X"70840552",
X"08575475",
X"5383e090",
X"085283e0",
X"940851fc",
X"c63f873d",
X"0d04ff3d",
X"0d737008",
X"53510293",
X"05337234",
X"70088105",
X"710c833d",
X"0d04fc3d",
X"0d873d88",
X"11557854",
X"99d25351",
X"fc993f80",
X"52873d51",
X"d13f863d",
X"0d04fd3d",
X"0d757052",
X"54a3c43f",
X"83e08008",
X"14537274",
X"2e9238ff",
X"13703353",
X"5371af2e",
X"098106ee",
X"38811353",
X"7283e080",
X"0c853d0d",
X"04fd3d0d",
X"75777053",
X"5454c73f",
X"83e08008",
X"732ea138",
X"83e08008",
X"733152ff",
X"125271ff",
X"2e8f3872",
X"70810554",
X"33747081",
X"055634eb",
X"39ff1454",
X"80743485",
X"3d0d0480",
X"3d0d7251",
X"ff903f82",
X"3d0d0471",
X"83e0800c",
X"04803d0d",
X"72518071",
X"34810bbc",
X"120c800b",
X"80c0120c",
X"823d0d04",
X"800b83e2",
X"d408248a",
X"38a4ae3f",
X"ff0b83e2",
X"d40c800b",
X"83e0800c",
X"04ff3d0d",
X"735283e0",
X"b008722e",
X"8d38d93f",
X"71519699",
X"3f7183e0",
X"b00c833d",
X"0d04f43d",
X"0d7e6062",
X"5c5a5581",
X"54bc1508",
X"81913874",
X"51cf3f79",
X"58807a25",
X"80f73883",
X"e3840870",
X"892a5783",
X"ff067884",
X"80723156",
X"56577378",
X"25833873",
X"557583e2",
X"d4082e84",
X"38ff893f",
X"83e2d408",
X"8025a638",
X"75892b51",
X"98dc3f83",
X"e384088f",
X"3dfc1155",
X"5c548152",
X"f81b5196",
X"c63f7614",
X"83e3840c",
X"7583e2d4",
X"0c745376",
X"527851a2",
X"df3f83e0",
X"800883e3",
X"84081683",
X"e3840c78",
X"7631761b",
X"5b595677",
X"8024ff8b",
X"38617a71",
X"0c547554",
X"75802e83",
X"38815473",
X"83e0800c",
X"8e3d0d04",
X"fc3d0dfe",
X"9b3f7651",
X"feaf3f86",
X"3dfc0553",
X"78527751",
X"95e93f79",
X"75710c54",
X"83e08008",
X"5483e080",
X"08802e83",
X"38815473",
X"83e0800c",
X"863d0d04",
X"fe3d0d75",
X"83e2d408",
X"53538072",
X"24893871",
X"732e8438",
X"fdd63f74",
X"51fdea3f",
X"725197ae",
X"3f83e080",
X"085283e0",
X"8008802e",
X"83388152",
X"7183e080",
X"0c843d0d",
X"04803d0d",
X"7280c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d72bc11",
X"0883e080",
X"0c51823d",
X"0d0480c4",
X"0b83e080",
X"0c04fd3d",
X"0d757771",
X"54705355",
X"539f9c3f",
X"82c81308",
X"bc150c82",
X"c0130880",
X"c0150cfc",
X"eb3f7351",
X"93ab3f73",
X"83e0b00c",
X"83e08008",
X"5383e080",
X"08802e83",
X"38815372",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"775553fc",
X"bf3f7280",
X"2ea538bc",
X"13085273",
X"519ea63f",
X"83e08008",
X"8f387752",
X"7251ff9a",
X"3f83e080",
X"08538a39",
X"82cc1308",
X"53d83981",
X"537283e0",
X"800c853d",
X"0d04fe3d",
X"0dff0b83",
X"e2d40c74",
X"83e0b40c",
X"7583e2d0",
X"0c9f933f",
X"83e08008",
X"81ff0652",
X"81537199",
X"3883e2ec",
X"518e943f",
X"83e08008",
X"5283e080",
X"08802e83",
X"38725271",
X"537283e0",
X"800c843d",
X"0d04fa3d",
X"0d787a82",
X"c4120882",
X"c4120870",
X"72245956",
X"56575773",
X"732e0981",
X"06913880",
X"c0165280",
X"c017519c",
X"973f83e0",
X"80085574",
X"83e0800c",
X"883d0d04",
X"f63d0d7c",
X"5b807b71",
X"5c54577a",
X"772e8c38",
X"811a82cc",
X"1408545a",
X"72f63880",
X"5980d939",
X"7a548157",
X"80707b7b",
X"315a5755",
X"ff185374",
X"732580c1",
X"3882cc14",
X"08527351",
X"ff8c3f80",
X"0b83e080",
X"0825a138",
X"82cc1408",
X"82cc1108",
X"82cc160c",
X"7482cc12",
X"0c537580",
X"2e863872",
X"82cc170c",
X"72548057",
X"7382cc15",
X"08811757",
X"5556ffb8",
X"39811959",
X"800bff1b",
X"54547873",
X"25833881",
X"54768132",
X"70750651",
X"5372ff90",
X"388c3d0d",
X"04f73d0d",
X"7b7d5a5a",
X"82d05283",
X"e2d00851",
X"80d08d3f",
X"83e08008",
X"57f9e13f",
X"795283e2",
X"d85195b5",
X"3f83e080",
X"08548053",
X"83e08008",
X"732e0981",
X"06828338",
X"83e0b408",
X"0b0b80f4",
X"98537052",
X"569bd43f",
X"0b0b80f4",
X"985280c0",
X"16519bc7",
X"3f75bc17",
X"0c7382c0",
X"170c810b",
X"82c4170c",
X"810b82c8",
X"170c7382",
X"cc170cff",
X"1782d017",
X"55578191",
X"3983e0c0",
X"3370822a",
X"70810651",
X"54557281",
X"80387481",
X"2a810658",
X"7780f638",
X"74842a81",
X"0682c415",
X"0c83e0c0",
X"33810682",
X"c8150c79",
X"5273519a",
X"ee3f7351",
X"9b853f83",
X"e0800814",
X"53af7370",
X"81055534",
X"72bc150c",
X"83e0c152",
X"72519acf",
X"3f83e0b8",
X"0882c015",
X"0c83e0ce",
X"5280c014",
X"519abc3f",
X"78802e8d",
X"38735178",
X"2d83e080",
X"08802e99",
X"387782cc",
X"150c7580",
X"2e863873",
X"82cc170c",
X"7382d015",
X"ff195955",
X"5676802e",
X"9b3883e0",
X"b85283e2",
X"d85194ab",
X"3f83e080",
X"088a3883",
X"e0c13353",
X"72fed238",
X"78802e89",
X"3883e0b4",
X"0851fcb8",
X"3f83e0b4",
X"08537283",
X"e0800c8b",
X"3d0d04ff",
X"3d0d8052",
X"7351fdb5",
X"3f833d0d",
X"04f03d0d",
X"62705254",
X"f6903f83",
X"e0800874",
X"53873d70",
X"535555f6",
X"b03ff790",
X"3f7351d3",
X"3f635374",
X"5283e080",
X"0851fab8",
X"3f923d0d",
X"047183e0",
X"800c0480",
X"c01283e0",
X"800c0480",
X"3d0d7282",
X"c0110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"82cc1108",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"7282c411",
X"0883e080",
X"0c51823d",
X"0d04f93d",
X"0d7983e0",
X"98085757",
X"81772781",
X"96387688",
X"17082781",
X"8e387533",
X"5574822e",
X"89387483",
X"2eb33880",
X"fe397454",
X"761083fe",
X"06537688",
X"2a8c1708",
X"0552893d",
X"fc055199",
X"c13f83e0",
X"800880df",
X"38029d05",
X"33893d33",
X"71882b07",
X"565680d1",
X"39845476",
X"822b83fc",
X"06537687",
X"2a8c1708",
X"0552893d",
X"fc055199",
X"913f83e0",
X"8008b038",
X"029f0533",
X"0284059e",
X"05337198",
X"2b71902b",
X"07028c05",
X"9d053370",
X"882b7207",
X"8d3d3371",
X"80fffffe",
X"80060751",
X"52535758",
X"56833981",
X"557483e0",
X"800c893d",
X"0d04fb3d",
X"0d83e098",
X"08fe1988",
X"1208fe05",
X"55565480",
X"56747327",
X"8d388214",
X"33757129",
X"94160805",
X"57537583",
X"e0800c87",
X"3d0d04fc",
X"3d0d7652",
X"800b83e0",
X"98087033",
X"51525370",
X"832e0981",
X"06913895",
X"12339413",
X"3371982b",
X"71902b07",
X"5555519b",
X"12339a13",
X"3371882b",
X"07740783",
X"e0800c55",
X"863d0d04",
X"fc3d0d76",
X"83e09808",
X"55558075",
X"23881508",
X"5372812e",
X"88388814",
X"08732685",
X"388152b2",
X"39729038",
X"73335271",
X"832e0981",
X"06853890",
X"14085372",
X"8c160c72",
X"802e8d38",
X"7251fed6",
X"3f83e080",
X"08528539",
X"90140852",
X"7190160c",
X"80527183",
X"e0800c86",
X"3d0d04fa",
X"3d0d7883",
X"e0980871",
X"22810570",
X"83ffff06",
X"57545755",
X"73802e88",
X"38901508",
X"53728638",
X"835280e7",
X"39738f06",
X"527180da",
X"38811390",
X"160c8c15",
X"08537290",
X"38830b84",
X"17225752",
X"73762780",
X"c638bf39",
X"821633ff",
X"0574842a",
X"065271b2",
X"387251fc",
X"b13f8152",
X"7183e080",
X"0827a838",
X"835283e0",
X"80088817",
X"08279c38",
X"83e08008",
X"8c160c83",
X"e0800851",
X"fdbc3f83",
X"e0800890",
X"160c7375",
X"23805271",
X"83e0800c",
X"883d0d04",
X"f23d0d60",
X"6264585e",
X"5b753355",
X"74a02e09",
X"81068838",
X"81167044",
X"56ef3962",
X"70335656",
X"74af2e09",
X"81068438",
X"81164380",
X"0b881c0c",
X"62703351",
X"55749f26",
X"91387a51",
X"fdd23f83",
X"e0800856",
X"807d3483",
X"8139933d",
X"841c0870",
X"58595f8a",
X"55a07670",
X"81055834",
X"ff155574",
X"ff2e0981",
X"06ef3880",
X"705a5c88",
X"7f085f5a",
X"7b811d70",
X"81ff0660",
X"13703370",
X"af327030",
X"a0732771",
X"80250751",
X"51525b53",
X"5e575574",
X"80e73876",
X"ae2e0981",
X"06833881",
X"55787a27",
X"75075574",
X"802e9f38",
X"79883270",
X"3078ae32",
X"70307073",
X"079f2a53",
X"51575156",
X"75bb3888",
X"598b5aff",
X"ab397698",
X"2b557480",
X"25873880",
X"f1ec1733",
X"57ff9f17",
X"55749926",
X"8938e017",
X"7081ff06",
X"58557881",
X"1a7081ff",
X"06721b53",
X"5b575576",
X"7534fef8",
X"397b1e7f",
X"0c805576",
X"a0268338",
X"8155748b",
X"19347a51",
X"fc823f83",
X"e0800880",
X"f538a054",
X"7a227085",
X"2b83e006",
X"5455901b",
X"08527c51",
X"93cc3f83",
X"e0800857",
X"83e08008",
X"8181387c",
X"33557480",
X"2e80f438",
X"8b1d3370",
X"832a7081",
X"06515656",
X"74b4388b",
X"7d841d08",
X"83e08008",
X"595b5b58",
X"ff185877",
X"ff2e9a38",
X"79708105",
X"5b337970",
X"81055b33",
X"71713152",
X"56567580",
X"2ee23886",
X"3975802e",
X"96387a51",
X"fbe53fff",
X"863983e0",
X"80085683",
X"e08008b6",
X"38833976",
X"56841b08",
X"8b113351",
X"5574a738",
X"8b1d3370",
X"842a7081",
X"06515656",
X"74893883",
X"56943981",
X"5690397c",
X"51fa943f",
X"83e08008",
X"881c0cfd",
X"81397583",
X"e0800c90",
X"3d0d04f8",
X"3d0d7a7c",
X"59578254",
X"83fe5377",
X"52765192",
X"913f8356",
X"83e08008",
X"80ec3881",
X"17337733",
X"71882b07",
X"56568256",
X"7482d4d5",
X"2e098106",
X"80d43875",
X"54b65377",
X"52765191",
X"e53f83e0",
X"80089838",
X"81173377",
X"3371882b",
X"0783e080",
X"08525656",
X"748182c6",
X"2eac3882",
X"5480d253",
X"77527651",
X"91bc3f83",
X"e0800898",
X"38811733",
X"77337188",
X"2b0783e0",
X"80085256",
X"56748182",
X"c62e8338",
X"81567583",
X"e0800c8a",
X"3d0d04eb",
X"3d0d675a",
X"800b83e0",
X"980c90de",
X"3f83e080",
X"08810655",
X"82567483",
X"ef387475",
X"538f3d70",
X"535759fe",
X"ca3f83e0",
X"800881ff",
X"06577681",
X"2e098106",
X"80d43890",
X"5483be53",
X"74527551",
X"90d03f83",
X"e0800880",
X"c9388f3d",
X"33557480",
X"2e80c938",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"0770587b",
X"575e525e",
X"575957fd",
X"ee3f83e0",
X"800881ff",
X"06577683",
X"2e098106",
X"86388156",
X"82f23976",
X"802e8638",
X"865682e8",
X"39a4548d",
X"53785275",
X"518fe73f",
X"815683e0",
X"800882d4",
X"3802be05",
X"33028405",
X"bd053371",
X"882b0759",
X"5d77ab38",
X"0280ce05",
X"33028405",
X"80cd0533",
X"71982b71",
X"902b0797",
X"3d337088",
X"2b720702",
X"940580cb",
X"05337107",
X"54525e57",
X"595602b7",
X"05337871",
X"29028805",
X"b6053302",
X"8c05b505",
X"3371882b",
X"07701d70",
X"7f8c050c",
X"5f595759",
X"5d8e3d33",
X"821b3402",
X"b9053390",
X"3d337188",
X"2b075a5c",
X"78841b23",
X"02bb0533",
X"028405ba",
X"05337188",
X"2b07565c",
X"74ab3802",
X"80ca0533",
X"02840580",
X"c9053371",
X"982b7190",
X"2b07963d",
X"3370882b",
X"72070294",
X"0580c705",
X"33710751",
X"5253575e",
X"5c747631",
X"78317984",
X"2a903d33",
X"54717131",
X"53565680",
X"c0f23f83",
X"e0800882",
X"0570881c",
X"0c83e080",
X"08e08a05",
X"56567483",
X"dffe2683",
X"38825783",
X"fff67627",
X"85388357",
X"89398656",
X"76802e80",
X"db38767a",
X"3476832e",
X"098106b0",
X"380280d6",
X"05330284",
X"0580d505",
X"3371982b",
X"71902b07",
X"993d3370",
X"882b7207",
X"02940580",
X"d3053371",
X"077f9005",
X"0c525e57",
X"58568639",
X"771b901b",
X"0c841a22",
X"8c1b0819",
X"71842a05",
X"941c0c5d",
X"800b811b",
X"347983e0",
X"980c8056",
X"7583e080",
X"0c973d0d",
X"04e93d0d",
X"83e09808",
X"56855475",
X"802e8182",
X"38800b81",
X"1734993d",
X"e011466a",
X"548a3d70",
X"5458ec05",
X"51f6e53f",
X"83e08008",
X"5483e080",
X"0880df38",
X"893d3354",
X"73802e91",
X"3802ab05",
X"3370842a",
X"81065155",
X"74802e86",
X"38835480",
X"c1397651",
X"f4893f83",
X"e08008a0",
X"170c02bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"3371079c",
X"1c0c5278",
X"981b0c53",
X"56595781",
X"0b811734",
X"74547383",
X"e0800c99",
X"3d0d04f5",
X"3d0d7d7f",
X"617283e0",
X"98085a5d",
X"5d595c80",
X"7b0c8557",
X"75802e81",
X"e0388116",
X"33810655",
X"84577480",
X"2e81d238",
X"91397481",
X"17348639",
X"800b8117",
X"34815781",
X"c0399c16",
X"08981708",
X"31557478",
X"27833874",
X"5877802e",
X"81a93898",
X"16087083",
X"ff065657",
X"7480cf38",
X"821633ff",
X"0577892a",
X"067081ff",
X"065a5578",
X"a0387687",
X"38a01608",
X"558d39a4",
X"160851f0",
X"e93f83e0",
X"80085581",
X"7527ffa8",
X"3874a417",
X"0ca41608",
X"51f2833f",
X"83e08008",
X"5583e080",
X"08802eff",
X"893883e0",
X"800819a8",
X"170c9816",
X"0883ff06",
X"84807131",
X"51557775",
X"27833877",
X"557483ff",
X"ff065498",
X"160883ff",
X"0653a816",
X"08527957",
X"7b83387b",
X"5776518a",
X"8d3f83e0",
X"8008fed0",
X"38981608",
X"1598170c",
X"741a7876",
X"317c0817",
X"7d0c595a",
X"fed33980",
X"577683e0",
X"800c8d3d",
X"0d04fa3d",
X"0d7883e0",
X"98085556",
X"85557380",
X"2e81e138",
X"81143381",
X"06538455",
X"72802e81",
X"d3389c14",
X"08537276",
X"27833872",
X"56981408",
X"57800b98",
X"150c7580",
X"2e81b738",
X"82143370",
X"892b5653",
X"76802eb5",
X"387452ff",
X"1651bbf4",
X"3f83e080",
X"08ff1876",
X"54705358",
X"53bbe53f",
X"83e08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed83f83",
X"e0800853",
X"810b83e0",
X"8008278b",
X"38881408",
X"83e08008",
X"26883880",
X"0b811534",
X"b03983e0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc73f",
X"83e08008",
X"8c3883e0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683e0",
X"800805a8",
X"150c8055",
X"7483e080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83e09808",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1d13f",
X"83e08008",
X"5583e080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef7",
X"3f83e080",
X"0888170c",
X"7551efa8",
X"3f83e080",
X"08557483",
X"e0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683e0",
X"9808802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f73f83e0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"86983f83",
X"e0800841",
X"83e08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"ede13f83",
X"e0800841",
X"83e08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"83a53f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f23f83e0",
X"80088332",
X"70307072",
X"079f2c83",
X"e0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"81b13f75",
X"83e0800c",
X"9e3d0d04",
X"fd3d0d75",
X"77535473",
X"33517089",
X"38713351",
X"70802ea1",
X"38733372",
X"33525372",
X"71278538",
X"ff519439",
X"70732785",
X"3881518b",
X"39811481",
X"135354d3",
X"39805170",
X"83e0800c",
X"853d0d04",
X"fd3d0d75",
X"77545472",
X"337081ff",
X"06525270",
X"802ea338",
X"7181ff06",
X"8114ffbf",
X"12535452",
X"70992689",
X"38a01270",
X"81ff0653",
X"51717470",
X"81055634",
X"d2398074",
X"34853d0d",
X"04ffbd3d",
X"0d80c63d",
X"0852a53d",
X"705254ff",
X"b33f80c7",
X"3d085285",
X"3d705253",
X"ffa63f72",
X"527351fe",
X"df3f80c5",
X"3d0d04fe",
X"3d0d7476",
X"53537170",
X"81055333",
X"51707370",
X"81055534",
X"70f03884",
X"3d0d04fe",
X"3d0d7452",
X"80723352",
X"5370732e",
X"8d388112",
X"81147133",
X"53545270",
X"f5387283",
X"e0800c84",
X"3d0d04fc",
X"3d0d7655",
X"7483e398",
X"082eaf38",
X"80537451",
X"87c13f83",
X"e0800881",
X"ff06ff14",
X"7081ff06",
X"7230709f",
X"2a515255",
X"53547280",
X"2e843871",
X"dd3873fe",
X"387483e3",
X"980c863d",
X"0d04ff3d",
X"0dff0b83",
X"e3980c84",
X"a53f8151",
X"87853f83",
X"e0800881",
X"ff065271",
X"ee3881d3",
X"3f7183e0",
X"800c833d",
X"0d04fc3d",
X"0d760284",
X"05a20522",
X"028805a6",
X"05227a54",
X"555555ff",
X"823f7280",
X"2ea03883",
X"e3ac1433",
X"75708105",
X"57348114",
X"7083ffff",
X"06ff1570",
X"83ffff06",
X"56525552",
X"dd39800b",
X"83e0800c",
X"863d0d04",
X"fc3d0d76",
X"787a1156",
X"53558053",
X"71742e93",
X"38721551",
X"703383e3",
X"ac133481",
X"12811454",
X"52ea3980",
X"0b83e080",
X"0c863d0d",
X"04fd3d0d",
X"905483e3",
X"98085186",
X"f43f83e0",
X"800881ff",
X"06ff1571",
X"30713070",
X"73079f2a",
X"729f2a06",
X"52555255",
X"5372db38",
X"853d0d04",
X"803d0d83",
X"e3a40810",
X"83e39c08",
X"079080a8",
X"0c823d0d",
X"04800b83",
X"e3a40ce4",
X"3f04810b",
X"83e3a40c",
X"db3f04ed",
X"3f047183",
X"e3a00c04",
X"803d0d80",
X"51f43f81",
X"0b83e3a4",
X"0c810b83",
X"e39c0cff",
X"bb3f823d",
X"0d04803d",
X"0d723070",
X"74078025",
X"83e39c0c",
X"51ffa53f",
X"823d0d04",
X"803d0d02",
X"8b053390",
X"80a40c90",
X"80a80870",
X"81065151",
X"70f53890",
X"80a40870",
X"81ff0683",
X"e0800c51",
X"823d0d04",
X"803d0d81",
X"ff51d13f",
X"83e08008",
X"81ff0683",
X"e0800c82",
X"3d0d0480",
X"3d0d7390",
X"2b730790",
X"80b40c82",
X"3d0d0404",
X"fb3d0d78",
X"0284059f",
X"05337098",
X"2b555755",
X"7280259b",
X"387580ff",
X"06568052",
X"80f751e0",
X"3f83e080",
X"0881ff06",
X"54738126",
X"80ff3880",
X"51fee73f",
X"ffa23f81",
X"51fedf3f",
X"ff9a3f75",
X"51feed3f",
X"74982a51",
X"fee63f74",
X"902a7081",
X"ff065253",
X"feda3f74",
X"882a7081",
X"ff065253",
X"fece3f74",
X"81ff0651",
X"fec63f81",
X"557580c0",
X"2e098106",
X"86388195",
X"558d3975",
X"80c82e09",
X"81068438",
X"81875574",
X"51fea53f",
X"8a55fec8",
X"3f83e080",
X"0881ff06",
X"70982b54",
X"54728025",
X"8c38ff15",
X"7081ff06",
X"565374e2",
X"387383e0",
X"800c873d",
X"0d04fa3d",
X"0dfdc53f",
X"8051fdda",
X"3f8a54fe",
X"933fff14",
X"7081ff06",
X"555373f3",
X"38737453",
X"5580c051",
X"fea63f83",
X"e0800881",
X"ff065473",
X"812e0981",
X"06829f38",
X"83aa5280",
X"c851fe8c",
X"3f83e080",
X"0881ff06",
X"5372812e",
X"09810681",
X"a8387454",
X"873d7411",
X"5456fdc8",
X"3f83e080",
X"08733481",
X"147081ff",
X"06555383",
X"7427e538",
X"029a0533",
X"5372812e",
X"09810681",
X"d938029b",
X"05335380",
X"ce905472",
X"81aa2e8d",
X"3881c739",
X"80e4518a",
X"b73fff14",
X"5473802e",
X"81b83882",
X"0a5281e9",
X"51fda53f",
X"83e08008",
X"81ff0653",
X"72de3872",
X"5280fa51",
X"fd923f83",
X"e0800881",
X"ff065372",
X"81903872",
X"54731653",
X"fcd63f83",
X"e0800873",
X"34811470",
X"81ff0655",
X"53837427",
X"e838873d",
X"3370862a",
X"70810651",
X"54548c55",
X"7280e338",
X"845580de",
X"39745281",
X"e951fccc",
X"3f83e080",
X"0881ff06",
X"53825581",
X"e9568173",
X"27863873",
X"5580c156",
X"80ce9054",
X"8a3980e4",
X"5189a93f",
X"ff145473",
X"802ea938",
X"80527551",
X"fc9a3f83",
X"e0800881",
X"ff065372",
X"e1388480",
X"5280d051",
X"fc863f83",
X"e0800881",
X"ff065372",
X"802e8338",
X"80557483",
X"e3a83480",
X"51fb873f",
X"fbc23f88",
X"3d0d04fb",
X"3d0d7754",
X"800b83e3",
X"a8337083",
X"2a708106",
X"51555755",
X"72752e09",
X"81068538",
X"73892b54",
X"735280d1",
X"51fbbd3f",
X"83e08008",
X"81ff0653",
X"72bd3882",
X"b8c054fb",
X"833f83e0",
X"800881ff",
X"06537281",
X"ff2e0981",
X"068938ff",
X"145473e7",
X"389f3972",
X"81fe2e09",
X"81069638",
X"83e7ac52",
X"83e3ac51",
X"faed3ffa",
X"d33ffad0",
X"3f833981",
X"558051fa",
X"893ffac4",
X"3f7481ff",
X"0683e080",
X"0c873d0d",
X"04fb3d0d",
X"7783e3ac",
X"56548151",
X"f9ec3f83",
X"e3a83370",
X"832a7081",
X"06515456",
X"72853873",
X"892b5473",
X"5280d851",
X"fab63f83",
X"e0800881",
X"ff065372",
X"80e43881",
X"ff51f9d4",
X"3f81fe51",
X"f9ce3f84",
X"80537470",
X"81055633",
X"51f9c13f",
X"ff137083",
X"ffff0651",
X"5372eb38",
X"7251f9b0",
X"3f7251f9",
X"ab3ff9d0",
X"3f83e080",
X"089f0653",
X"a7885472",
X"852e8c38",
X"993980e4",
X"5186e13f",
X"ff1454f9",
X"b33f83e0",
X"800881ff",
X"2e843873",
X"e9388051",
X"f8e43ff9",
X"9f3f800b",
X"83e0800c",
X"873d0d04",
X"7183e7b0",
X"0c888080",
X"0b83e7ac",
X"0c848080",
X"0b83e7b4",
X"0c04fd3d",
X"0d777017",
X"557705ff",
X"1a535371",
X"ff2e9438",
X"73708105",
X"55335170",
X"73708105",
X"5534ff12",
X"52e93985",
X"3d0d04fc",
X"3d0d87a6",
X"81557433",
X"83e7b834",
X"a05483a0",
X"805383e7",
X"b0085283",
X"e7ac0851",
X"ffb83fa0",
X"5483a480",
X"5383e7b0",
X"085283e7",
X"ac0851ff",
X"a53f9054",
X"83a88053",
X"83e7b008",
X"5283e7ac",
X"0851ff92",
X"3fa05380",
X"5283e7b4",
X"0883a080",
X"055185b9",
X"3fa05380",
X"5283e7b4",
X"0883a480",
X"055185a9",
X"3f905380",
X"5283e7b4",
X"0883a880",
X"05518599",
X"3fff7534",
X"83a08054",
X"805383e7",
X"b0085283",
X"e7b40851",
X"fecc3f80",
X"d0805483",
X"b0805383",
X"e7b00852",
X"83e7b408",
X"51feb73f",
X"86cc3fa2",
X"54805383",
X"e7b4088c",
X"80055280",
X"f79c51fe",
X"a13f860b",
X"87a88334",
X"800b87a8",
X"8234800b",
X"87a09a34",
X"af0b87a0",
X"9634bf0b",
X"87a09734",
X"800b87a0",
X"98349f0b",
X"87a09934",
X"800b87a0",
X"9b34e00b",
X"87a88934",
X"a20b87a8",
X"8034830b",
X"87a48f34",
X"820b87a8",
X"8134863d",
X"0d04fd3d",
X"0d83a080",
X"54805383",
X"e7b40852",
X"83e7b008",
X"51fdbf3f",
X"80d08054",
X"83b08053",
X"83e7b408",
X"5283e7b0",
X"0851fdaa",
X"3fa05483",
X"a0805383",
X"e7b40852",
X"83e7b008",
X"51fd973f",
X"a05483a4",
X"805383e7",
X"b4085283",
X"e7b00851",
X"fd843f90",
X"5483a880",
X"5383e7b4",
X"085283e7",
X"b00851fc",
X"f13f83e7",
X"b83387a6",
X"8134853d",
X"0d04803d",
X"0d908090",
X"08810683",
X"e0800c82",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fe067607",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"812c8106",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fd06",
X"76100772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087082",
X"2cbf0683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fe8306",
X"76822b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"882c8706",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870f1ff",
X"0676882b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"708b2cbf",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870f8",
X"8fff0676",
X"8b2b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"90087091",
X"2cbf0683",
X"e0800c51",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fc87ff",
X"ff067691",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870992c",
X"810683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"ffbf0a06",
X"76992b07",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80800870",
X"882c8106",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"70892c81",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708a2c",
X"810683e0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708b",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"fe3d0d74",
X"81e62987",
X"2a9080a0",
X"0c843d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727081",
X"055434ff",
X"1151f039",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708405",
X"540cff11",
X"51f03984",
X"3d0d04fe",
X"3d0d8480",
X"80538052",
X"88800a51",
X"ffb33f81",
X"80805380",
X"5282800a",
X"51c63f84",
X"3d0d0480",
X"3d0d8151",
X"fc913f72",
X"802e9038",
X"8051fe93",
X"3fcd3f83",
X"e7bc3351",
X"fe893f81",
X"51fca23f",
X"8051fc9d",
X"3f8051fb",
X"ee3f823d",
X"0d04fd3d",
X"0d755280",
X"5480ff72",
X"25883881",
X"0bff8013",
X"5354ffbf",
X"12517099",
X"268638e0",
X"12529e39",
X"ff9f1251",
X"99712795",
X"38d012e0",
X"13705454",
X"51897127",
X"88388f73",
X"27833880",
X"5273802e",
X"85388180",
X"12527181",
X"ff0683e0",
X"800c853d",
X"0d04803d",
X"0d84d8c0",
X"51807170",
X"81055334",
X"7084e0c0",
X"2e098106",
X"f038823d",
X"0d04fe3d",
X"0d029705",
X"3351ff86",
X"3f83e080",
X"0881ff06",
X"83e7c008",
X"54528073",
X"249b3883",
X"e7e00813",
X"7283e7e4",
X"08075353",
X"71733483",
X"e7c00881",
X"0583e7c0",
X"0c843d0d",
X"04fa3d0d",
X"82800a1b",
X"55805788",
X"3dfc0554",
X"79537452",
X"7851cbe8",
X"3f883d0d",
X"04fe3d0d",
X"83e7d808",
X"527451d2",
X"cc3f83e0",
X"80088c38",
X"76537552",
X"83e7d808",
X"51c73f84",
X"3d0d04fe",
X"3d0d83e7",
X"d8085375",
X"527451cd",
X"8b3f83e0",
X"80088d38",
X"77537652",
X"83e7d808",
X"51ffa23f",
X"843d0d04",
X"fe3d0d83",
X"e7d80851",
X"cbff3f83",
X"e0800881",
X"80802e09",
X"81068838",
X"83c18080",
X"539b3983",
X"e7d80851",
X"cbe33f83",
X"e0800880",
X"d0802e09",
X"81069338",
X"83c1b080",
X"5383e080",
X"085283e7",
X"d80851fe",
X"d83f843d",
X"0d04803d",
X"0df9f93f",
X"83e08008",
X"842980f7",
X"c0057008",
X"83e0800c",
X"51823d0d",
X"04ee3d0d",
X"80438042",
X"80418070",
X"5a5bfdd2",
X"3f800b83",
X"e7c00c80",
X"0b83e7e4",
X"0c80f590",
X"51c6cf3f",
X"81800b83",
X"e7e40c80",
X"f59451c6",
X"c13f80d0",
X"0b83e7c0",
X"0c783070",
X"7a078025",
X"70872b83",
X"e7e40c51",
X"55f8ec3f",
X"83e08008",
X"5280f59c",
X"51c69b3f",
X"80f80b83",
X"e7c00c78",
X"81327030",
X"70720780",
X"2570872b",
X"83e7e40c",
X"515656fe",
X"f13f83e0",
X"80085280",
X"f5a851c5",
X"f13f81a0",
X"0b83e7c0",
X"0c788232",
X"70307072",
X"07802570",
X"872b83e7",
X"e40c5156",
X"83e7d808",
X"5256c78b",
X"3f83e080",
X"085280f5",
X"b051c5c2",
X"3f81f00b",
X"83e7c00c",
X"810b83e7",
X"c45b5883",
X"e7c00882",
X"197a3270",
X"30707207",
X"80257087",
X"2b83e7e4",
X"0c51578e",
X"3d7055ff",
X"1b545757",
X"579a813f",
X"79708405",
X"5b0851c6",
X"c23f7454",
X"83e08008",
X"53775280",
X"f5b851c4",
X"f53fa817",
X"83e7c00c",
X"81185877",
X"852e0981",
X"06ffb038",
X"83900b83",
X"e7c00c78",
X"87327030",
X"70720780",
X"2570872b",
X"83e7e40c",
X"515656f8",
X"923f80f5",
X"c85583e0",
X"8008802e",
X"8e3883e7",
X"d40851c5",
X"ee3f83e0",
X"80085574",
X"5280f5d0",
X"51c4a33f",
X"83e00b83",
X"e7c00c78",
X"88327030",
X"70720780",
X"2570872b",
X"83e7e40c",
X"515780f5",
X"dc5255c4",
X"813f868d",
X"a051f8f8",
X"3f805291",
X"3d705255",
X"9ad33f83",
X"5274519a",
X"cc3f6119",
X"59788025",
X"85388059",
X"90398879",
X"25853888",
X"59873978",
X"882682db",
X"3878822b",
X"5580f3ec",
X"150804f6",
X"863f83e0",
X"80086157",
X"5575812e",
X"09810689",
X"3883e080",
X"08105590",
X"3975ff2e",
X"09810688",
X"3883e080",
X"08812c55",
X"90752585",
X"38905588",
X"39748024",
X"83388155",
X"7451f5e0",
X"3f829039",
X"f5f23f83",
X"e0800861",
X"05557480",
X"25853880",
X"55883987",
X"75258338",
X"87557451",
X"f5eb3f81",
X"ee396087",
X"3862802e",
X"81e53883",
X"e0a40883",
X"e0a00c8b",
X"df0b83e0",
X"a80c83e7",
X"d80851ff",
X"b59f3ffa",
X"e73f81c7",
X"39605680",
X"76259938",
X"8af80b83",
X"e0a80c83",
X"e7b81570",
X"085255ff",
X"b4ff3f74",
X"08529139",
X"75802591",
X"3883e7b8",
X"150851c3",
X"dc3f8052",
X"fd1951b8",
X"3962802e",
X"818d3883",
X"e7b81570",
X"0883e7c4",
X"08720c83",
X"e7c40cfd",
X"1a705351",
X"558bf13f",
X"83e08008",
X"5680518b",
X"e73f83e0",
X"80085274",
X"5187ff3f",
X"75528051",
X"87f83f80",
X"d6396055",
X"807525b8",
X"3883e0ac",
X"0883e0a0",
X"0c8bdf0b",
X"83e0a80c",
X"83e7d408",
X"51ffb489",
X"3f83e7d4",
X"0851ffb1",
X"a33f83e0",
X"800881ff",
X"06705255",
X"f4f63f74",
X"802e9c38",
X"8155a039",
X"74802593",
X"3883e7d4",
X"0851c2cd",
X"3f8051f4",
X"db3f8439",
X"6287387a",
X"802efa8a",
X"38805574",
X"83e0800c",
X"943d0d04",
X"fe3d0df5",
X"873f83e0",
X"8008802e",
X"86388051",
X"818b39f5",
X"8c3f83e0",
X"800880ff",
X"38f5ac3f",
X"83e08008",
X"802eb938",
X"8151f2bb",
X"3f8051f4",
X"c23fefaf",
X"3f800b83",
X"e7c00cf9",
X"b43f83e0",
X"800853ff",
X"0b83e7c0",
X"0cf19b3f",
X"7280cc38",
X"83e7bc33",
X"51f49c3f",
X"7251f28b",
X"3f80c139",
X"f4d43f83",
X"e0800880",
X"2eb63881",
X"51f1f83f",
X"8051f3ff",
X"3feeec3f",
X"8af80b83",
X"e0a80c83",
X"e7c40851",
X"ffb2ba3f",
X"ff0b83e7",
X"c00cf0d6",
X"3f83e7c4",
X"08528051",
X"85f43f81",
X"51f5b03f",
X"843d0d04",
X"fb3d0d80",
X"0b83e7bc",
X"34908080",
X"52868480",
X"8051c586",
X"3f83e080",
X"08819338",
X"89bf3f80",
X"f99451c9",
X"c63f83e0",
X"8008559c",
X"800a5480",
X"c0805380",
X"f5e45283",
X"e0800851",
X"f7853f83",
X"e7d80853",
X"80f5f452",
X"7451c490",
X"3f83e080",
X"088438f7",
X"933f83e7",
X"dc085380",
X"f6805274",
X"51c3f93f",
X"83e08008",
X"b538873d",
X"fc055484",
X"80805386",
X"a8808052",
X"83e7dc08",
X"51c2853f",
X"83e08008",
X"93387584",
X"80802e09",
X"81068938",
X"810b83e7",
X"bc348739",
X"800b83e7",
X"bc3483e7",
X"bc3351f2",
X"aa3f8151",
X"f4813f92",
X"fb3f8151",
X"f3f93ffd",
X"a73ffc39",
X"83e08c08",
X"0283e08c",
X"0cfb3d0d",
X"0280f68c",
X"0b83e0a4",
X"0c80f690",
X"0b83e09c",
X"0c80f694",
X"0b83e0ac",
X"0c83e08c",
X"08fc050c",
X"800b83e7",
X"c40b83e0",
X"8c08f805",
X"0c83e08c",
X"08f4050c",
X"c2983f83",
X"e0800886",
X"05fc0683",
X"e08c08f0",
X"050c0283",
X"e08c08f0",
X"0508310d",
X"833d7083",
X"e08c08f8",
X"05087084",
X"0583e08c",
X"08f8050c",
X"0c51ffbe",
X"e03f83e0",
X"8c08f405",
X"08810583",
X"e08c08f4",
X"050c83e0",
X"8c08f405",
X"08872e09",
X"8106ffac",
X"38869480",
X"8051ebac",
X"3fff0b83",
X"e7c00c80",
X"0b83e7e4",
X"0c84d8c0",
X"0b83e7e0",
X"0c8151ee",
X"d63f8151",
X"eefb3f80",
X"51eef63f",
X"8151ef9c",
X"3f8151ef",
X"f13f8251",
X"efbf3f80",
X"51f0953f",
X"8051f0bf",
X"3f80d0be",
X"528051ff",
X"bc993ffc",
X"e33f83e0",
X"8c08fc05",
X"080d800b",
X"83e0800c",
X"873d0d83",
X"e08c0c04",
X"803d0d81",
X"ff51800b",
X"83e7f012",
X"34ff1151",
X"70f43882",
X"3d0d04ff",
X"3d0d7370",
X"33535181",
X"11337134",
X"71811234",
X"833d0d04",
X"fb3d0d77",
X"79565680",
X"70715555",
X"52717525",
X"ac387216",
X"70337014",
X"7081ff06",
X"55515151",
X"71742789",
X"38811270",
X"81ff0653",
X"51718114",
X"7083ffff",
X"06555254",
X"747324d6",
X"387183e0",
X"800c873d",
X"0d04fc3d",
X"0d7655ff",
X"b5c53f83",
X"e0800880",
X"2ef53883",
X"ea8c0886",
X"057081ff",
X"065253ff",
X"b3c53f84",
X"39fa913f",
X"ffb5a43f",
X"83e08008",
X"812ef238",
X"80547315",
X"53ffb48a",
X"3f83e080",
X"08733481",
X"14547385",
X"2e098106",
X"e9388439",
X"f9e63fff",
X"b4f93f83",
X"e0800880",
X"2ef23874",
X"3383e7f0",
X"34811533",
X"83e7f134",
X"82153383",
X"e7f23483",
X"153383e7",
X"f3348452",
X"83e7f051",
X"feba3f83",
X"e0800881",
X"ff068416",
X"33565372",
X"752e0981",
X"068d38ff",
X"b3ee3f83",
X"e0800880",
X"2e9a3883",
X"ea8c08a8",
X"2e098106",
X"8938860b",
X"83ea8c0c",
X"8739a80b",
X"83ea8c0c",
X"80e451ee",
X"d73f863d",
X"0d04f43d",
X"0d7e6059",
X"55805d80",
X"75822b71",
X"83ea9012",
X"0c83eaa4",
X"175b5b57",
X"76793477",
X"772e83b8",
X"38765277",
X"51ffbda4",
X"3f8e3dfc",
X"05549053",
X"83e9f852",
X"7751ffbc",
X"df3f7c56",
X"75902e09",
X"81068394",
X"3883e9f8",
X"51fd943f",
X"83e9fa51",
X"fd8d3f83",
X"e9fc51fd",
X"863f7683",
X"ea880c77",
X"51ffbaab",
X"3f80f4a0",
X"5283e080",
X"0851ffa9",
X"e53f83e0",
X"8008812e",
X"09810680",
X"d4387683",
X"eaa00c82",
X"0b83e9f8",
X"34ff960b",
X"83e9f934",
X"7751ffbc",
X"f03f83e0",
X"80085583",
X"e0800877",
X"25883883",
X"e080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583e9fa",
X"347483e9",
X"fb347683",
X"e9fc34ff",
X"800b83e9",
X"fd348190",
X"3983e9f8",
X"3383e9f9",
X"3371882b",
X"07565b74",
X"83ffff2e",
X"09810680",
X"e838fe80",
X"0b83eaa0",
X"0c810b83",
X"ea880cff",
X"0b83e9f8",
X"34ff0b83",
X"e9f93477",
X"51ffbbfd",
X"3f83e080",
X"0883eaa8",
X"0c83e080",
X"085583e0",
X"80088025",
X"883883e0",
X"80088f05",
X"5574842c",
X"7083ffff",
X"0670882a",
X"58515575",
X"83e9fa34",
X"7483e9fb",
X"347683e9",
X"fc34ff80",
X"0b83e9fd",
X"34810b83",
X"ea8734a5",
X"39748596",
X"2e098106",
X"80fe3875",
X"83eaa00c",
X"7751ffbb",
X"b13f83ea",
X"873383e0",
X"80080755",
X"7483ea87",
X"3483ea87",
X"33810655",
X"74802e83",
X"38845783",
X"e9fc3383",
X"e9fd3371",
X"882b0756",
X"5c748180",
X"2e098106",
X"a13883e9",
X"fa3383e9",
X"fb337188",
X"2b07565b",
X"ad807527",
X"87387682",
X"07579c39",
X"76810757",
X"96397482",
X"802e0981",
X"06873876",
X"83075787",
X"397481ff",
X"268a3877",
X"83ea901b",
X"0c767934",
X"8e3d0d04",
X"803d0d72",
X"842983ea",
X"90057008",
X"83e0800c",
X"51823d0d",
X"04fe3d0d",
X"800b83e9",
X"f40c800b",
X"83e9f00c",
X"ff0b83e7",
X"ec0ca80b",
X"83ea8c0c",
X"ae51ffae",
X"8e3f800b",
X"83ea9054",
X"52807370",
X"8405550c",
X"81125271",
X"842e0981",
X"06ef3884",
X"3d0d04fe",
X"3d0d7402",
X"84059605",
X"22535371",
X"802e9738",
X"72708105",
X"543351ff",
X"ae983fff",
X"127083ff",
X"ff065152",
X"e639843d",
X"0d04fe3d",
X"0d029205",
X"225382ac",
X"51e9e93f",
X"80c351ff",
X"adf43f81",
X"9651e9dc",
X"3f725283",
X"e7f051ff",
X"b23f7252",
X"83e7f051",
X"f8ee3f83",
X"e0800881",
X"ff0651ff",
X"add03f84",
X"3d0d04ff",
X"b13d0d80",
X"d13df805",
X"51f9973f",
X"83e9f408",
X"810583e9",
X"f40c80cf",
X"3d33cf11",
X"7081ff06",
X"51565674",
X"832688ed",
X"38758f06",
X"ff055675",
X"83e7ec08",
X"2e9b3875",
X"83269638",
X"7583e7ec",
X"0c758429",
X"83ea9005",
X"70085355",
X"7551fa96",
X"3f807624",
X"88c93875",
X"842983ea",
X"90055574",
X"08802e88",
X"ba3883e7",
X"ec088429",
X"83ea9005",
X"70080288",
X"0582b905",
X"33525b55",
X"7480d22e",
X"84b13874",
X"80d22490",
X"3874bf2e",
X"9c387480",
X"d02e81d7",
X"3887f839",
X"7480d32e",
X"80d23874",
X"80d72e81",
X"c63887e7",
X"390282bb",
X"05330284",
X"0582ba05",
X"33718280",
X"29055656",
X"ffaccc3f",
X"80c151ff",
X"ac843ff6",
X"e73f860b",
X"83e7f034",
X"815283e7",
X"f051ffad",
X"a73f8151",
X"fde43f74",
X"8938860b",
X"83ea8c0c",
X"8739a80b",
X"83ea8c0c",
X"ffac983f",
X"80c151ff",
X"abd03ff6",
X"b33f900b",
X"83ea8733",
X"81065656",
X"74802e83",
X"38985683",
X"e9fc3383",
X"e9fd3371",
X"882b0756",
X"59748180",
X"2e098106",
X"9c3883e9",
X"fa3383e9",
X"fb337188",
X"2b075657",
X"ad807527",
X"8c387581",
X"80075685",
X"3975a007",
X"567583e7",
X"f034ff0b",
X"83e7f134",
X"e00b83e7",
X"f234800b",
X"83e7f334",
X"845283e7",
X"f051ffac",
X"9b3f8451",
X"869e3902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"5659ffab",
X"8a3f7951",
X"ffb5f73f",
X"83e08008",
X"802e8b38",
X"80ce51ff",
X"aab43f85",
X"f23980c1",
X"51ffaaaa",
X"3fffab9f",
X"3fffa9d2",
X"3f83eaa0",
X"08588375",
X"259b3883",
X"e9fc3383",
X"e9fd3371",
X"882b07fc",
X"1771297a",
X"05838005",
X"5a51578d",
X"39748180",
X"2918ff80",
X"05588180",
X"57805676",
X"762e9338",
X"ffaa833f",
X"83e08008",
X"83e7f017",
X"34811656",
X"ea39ffa9",
X"f13f83e0",
X"800881ff",
X"06775383",
X"e7f05256",
X"f4d63f83",
X"e0800881",
X"ff065575",
X"752e0981",
X"06818a38",
X"ffa9f03f",
X"80c151ff",
X"a9a83fff",
X"aa9d3f77",
X"527951ff",
X"b4863f80",
X"5e80d13d",
X"fdf40554",
X"765383e7",
X"f0527951",
X"ffb2933f",
X"0282b905",
X"33558158",
X"7480d72e",
X"098106bd",
X"3880d13d",
X"fdf00554",
X"76538f3d",
X"70537a52",
X"59ffb398",
X"3f805676",
X"762ea238",
X"751983e7",
X"f0173371",
X"33707232",
X"70307080",
X"2570307e",
X"06811d5d",
X"5e515151",
X"525b55db",
X"3982ac51",
X"e4a23f77",
X"802e8638",
X"80c35184",
X"3980ce51",
X"ffa8a33f",
X"ffa9983f",
X"ffa7cb3f",
X"83dd3902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"59558070",
X"5d59ffa8",
X"be3f80c1",
X"51ffa7f6",
X"3f83ea88",
X"08792e82",
X"de3883ea",
X"a80880fc",
X"055580fd",
X"52745186",
X"d73f83e0",
X"80085b77",
X"8224b238",
X"ff187087",
X"2b83ffff",
X"800680f7",
X"e00583e7",
X"f0595755",
X"81805575",
X"70810557",
X"33777081",
X"055934ff",
X"157081ff",
X"06515574",
X"ea38828d",
X"397782e8",
X"2e81ab38",
X"7782e92e",
X"09810681",
X"b23880f6",
X"9851ffad",
X"f93f7858",
X"77873270",
X"30707207",
X"80257a8a",
X"32703070",
X"72078025",
X"73075354",
X"5a515755",
X"75802e97",
X"38787826",
X"9238a00b",
X"83e7f01a",
X"34811970",
X"81ff065a",
X"55eb3981",
X"187081ff",
X"0659558a",
X"7827ffbc",
X"388f5883",
X"e7eb1833",
X"83e7f019",
X"34ff1870",
X"81ff0659",
X"55778426",
X"ea389058",
X"800b83e7",
X"f0193481",
X"187081ff",
X"0670982b",
X"52595574",
X"8025e938",
X"80c6557a",
X"858f2484",
X"3880c255",
X"7483e7f0",
X"3480f10b",
X"83e7f334",
X"810b83e7",
X"f4347a83",
X"e7f1347a",
X"882c5574",
X"83e7f234",
X"80cb3982",
X"f0782580",
X"c4387780",
X"fd29fd97",
X"d3055279",
X"51ffb0b4",
X"3f80d13d",
X"fdec0554",
X"80fd5383",
X"e7f05279",
X"51ffafec",
X"3f7b8119",
X"59567580",
X"fc248338",
X"78587788",
X"2c557483",
X"e8ed3477",
X"83e8ee34",
X"7583e8ef",
X"34818059",
X"80cc3983",
X"eaa00857",
X"8378259b",
X"3883e9fc",
X"3383e9fd",
X"3371882b",
X"07fc1a71",
X"29790583",
X"80055951",
X"598d3977",
X"81802917",
X"ff800557",
X"81805976",
X"527951ff",
X"afc23f80",
X"d13dfdec",
X"05547853",
X"83e7f052",
X"7951ffae",
X"fb3f7851",
X"f6b83fff",
X"a5b53fff",
X"a3e83f8b",
X"3983e9f0",
X"08810583",
X"e9f00c80",
X"d13d0d04",
X"f6d93fea",
X"af3ff939",
X"fc3d0d76",
X"78718429",
X"83ea9005",
X"70085153",
X"5353709e",
X"3880ce72",
X"3480cf0b",
X"81133480",
X"ce0b8213",
X"3480c50b",
X"83133470",
X"84133480",
X"e73983ea",
X"a4133354",
X"80d27234",
X"73822a70",
X"81065151",
X"80cf5370",
X"843880d7",
X"53728113",
X"34a00b82",
X"13347383",
X"06517081",
X"2e9e3870",
X"81248838",
X"70802e8f",
X"389f3970",
X"822e9238",
X"70832e92",
X"38933980",
X"d8558e39",
X"80d35589",
X"3980cd55",
X"843980c4",
X"55748313",
X"3480c40b",
X"84133480",
X"0b851334",
X"863d0d04",
X"fd3d0d75",
X"5380730c",
X"800b8414",
X"0c800b88",
X"140c87a6",
X"80337081",
X"ff067081",
X"2a813271",
X"81327181",
X"06718106",
X"3184180c",
X"55567083",
X"2a813271",
X"822a8132",
X"71810671",
X"81063177",
X"0c525451",
X"5187a090",
X"33700981",
X"0688150c",
X"51853d0d",
X"04fe3d0d",
X"74765452",
X"7151ffa0",
X"3f72812e",
X"a2388173",
X"268d3872",
X"822eab38",
X"72832e9f",
X"38e63971",
X"08e23884",
X"1208dd38",
X"881208d8",
X"38a03988",
X"1208812e",
X"098106cc",
X"38943988",
X"1208812e",
X"8d387108",
X"89388412",
X"08802eff",
X"b738843d",
X"0d04fc3d",
X"0d767853",
X"54815380",
X"55873971",
X"10731054",
X"52737226",
X"5172802e",
X"a7387080",
X"2e863871",
X"8025e838",
X"72802e98",
X"38717426",
X"89387372",
X"31757407",
X"56547281",
X"2a72812a",
X"5353e539",
X"73517883",
X"38745170",
X"83e0800c",
X"863d0d04",
X"fe3d0d80",
X"53755274",
X"51ffa33f",
X"843d0d04",
X"fe3d0d81",
X"53755274",
X"51ff933f",
X"843d0d04",
X"fb3d0d77",
X"79555580",
X"56747625",
X"86387430",
X"55815673",
X"80258838",
X"73307681",
X"32575480",
X"53735274",
X"51fee73f",
X"83e08008",
X"5475802e",
X"873883e0",
X"80083054",
X"7383e080",
X"0c873d0d",
X"04fa3d0d",
X"787a5755",
X"80577477",
X"25863874",
X"30558157",
X"759f2c54",
X"81537574",
X"32743152",
X"7451feaa",
X"3f83e080",
X"08547680",
X"2e873883",
X"e0800830",
X"547383e0",
X"800c883d",
X"0d040000",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002aef",
X"00002b30",
X"00002b52",
X"00002b79",
X"00002b79",
X"00002b79",
X"00002b79",
X"00002bea",
X"00002c3c",
X"25732025",
X"73000000",
X"2e2e0000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"54757262",
X"6f3a2564",
X"78000000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"66726565",
X"7a65722e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"6e616d65",
X"20000000",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00003a4c",
X"00003a50",
X"00003a58",
X"00003a64",
X"00003a70",
X"00003a7c",
X"00003a88",
X"00003a8c",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"2f737973",
X"74656d2f",
X"726f6d2f",
X"61746172",
X"69383030",
X"00000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
